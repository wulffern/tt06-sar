* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
*+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
*+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7]
*+ ui_in[0] uo_out[6] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=240.8616 ps=1.269k w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=244.62 ps=1.28028k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X51 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X52 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X56 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X58 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X63 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X65 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X66 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X72 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X74 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X76 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X77 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X78 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X79 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 VPWR SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X88 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X90 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X95 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X96 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X97 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X98 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R8 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X99 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X100 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X101 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X106 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X107 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X108 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X114 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X115 SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X116 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 VGND SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X118 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R10 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X119 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X120 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X121 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X122 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X124 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X125 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X130 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X131 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X132 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X134 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X135 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X136 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X137 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X146 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X147 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X148 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X149 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X150 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X155 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R13 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X158 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X160 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X163 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X166 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R14 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X167 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X169 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X174 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X175 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R15 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X176 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X177 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X178 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X181 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X185 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X186 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X188 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X193 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X194 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X195 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X198 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R16 uio_oe[0] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R17 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X199 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X201 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R18 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X205 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X206 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X207 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 VGND SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R19 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X212 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X213 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X214 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X216 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X221 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X223 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X225 SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X228 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X229 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X230 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X232 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X233 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X235 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X236 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X237 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X239 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X244 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X246 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X250 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X253 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X255 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X260 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X263 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X266 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X267 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X268 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X270 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X275 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X276 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X278 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X280 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R23 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R24 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X282 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X284 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X286 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X288 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X292 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X294 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X295 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X300 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X307 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X308 VPWR SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X309 VGND SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X310 SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X311 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X312 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X313 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X314 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R25 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R26 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X316 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X318 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X321 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X322 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XB2.XA3.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X324 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R27 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X328 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X333 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X337 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X338 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X341 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X342 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X344 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R29 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X346 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X347 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X348 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X349 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X351 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X352 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R30 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X359 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X360 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X364 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R31 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X365 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X366 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R32 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X368 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X370 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X371 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X372 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X373 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X374 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X375 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X376 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X377 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X378 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X379 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R34 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X381 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X382 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X384 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X385 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X386 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X387 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R35 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X388 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X389 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X390 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X391 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X393 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X394 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X395 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X400 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X402 SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X404 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R36 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R37 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X407 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X410 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X413 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X414 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X416 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X417 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X418 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X419 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X420 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X421 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X422 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R38 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X423 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X424 SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X425 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X426 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X427 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X428 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X429 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X433 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X434 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X435 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X436 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X437 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X440 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X441 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X442 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R41 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X443 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X447 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X449 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X450 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X452 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X453 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X454 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X455 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R42 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X457 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R43 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X458 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X459 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X462 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X463 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X465 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X468 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R44 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X470 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X471 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X472 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X473 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X474 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X477 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X478 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X479 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X480 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X481 VGND SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X482 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X484 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X486 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X489 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X491 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X492 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X493 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X494 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X496 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R46 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X498 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X499 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X500 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X501 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X502 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X503 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X505 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X506 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X508 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R48 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X509 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X510 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X511 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X512 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X513 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X514 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X515 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X516 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X517 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X519 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X520 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X521 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X522 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R49 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X525 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X526 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X527 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X528 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X530 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X532 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X533 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X536 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X537 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XA20.XA10.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X540 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X541 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X544 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R51 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X545 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X548 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X553 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X554 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X557 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X558 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X560 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X561 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X562 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X564 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X565 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X567 SUNSAR_CAPT8B_CV_0.XA2.MN0.G SUNSAR_CAPT8B_CV_0.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X568 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X569 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X570 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X571 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X572 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X573 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X574 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X575 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X578 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X579 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X580 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X581 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X582 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X583 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X584 SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R53 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X586 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X587 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X588 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X589 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X590 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X591 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X592 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R54 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X593 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X594 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X595 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X596 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X598 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VGND SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X601 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X602 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X603 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X604 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X605 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X606 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X609 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X610 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X612 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X613 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X614 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X616 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X618 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X619 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X621 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X624 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X625 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X626 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X631 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X632 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R55 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X635 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X637 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X640 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X642 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X644 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X645 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X647 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X648 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X649 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X650 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X652 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X653 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X654 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X655 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X656 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R57 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R58 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X657 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X658 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X660 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X661 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X663 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X664 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X665 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X666 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X667 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X669 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X670 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X671 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X674 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X675 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X676 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X677 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X679 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X680 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X681 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X682 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X683 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X684 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X685 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R60 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X686 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X687 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X688 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X690 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X691 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X693 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X694 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X695 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X696 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X697 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X699 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X700 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X701 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X704 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X705 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R61 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X706 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X707 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X709 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X710 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X713 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X714 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R62 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X715 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X716 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X717 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X718 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X719 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X720 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X721 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X722 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X723 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X726 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X727 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X728 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X729 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X730 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X731 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X732 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X733 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X734 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X735 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X738 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X739 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R65 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X740 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X741 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X742 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X743 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X745 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X746 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X747 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X749 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X751 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X752 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X753 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X754 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X755 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R67 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X758 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X759 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X760 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X762 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X763 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X765 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X766 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X767 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X768 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X769 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X770 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R68 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X771 VGND SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X773 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X774 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X776 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X777 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X778 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X779 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X780 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X781 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X782 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X783 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X786 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X787 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X788 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X790 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X791 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X792 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X793 SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X794 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X796 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X798 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X800 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X802 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X804 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X809 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X810 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X811 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X813 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X814 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X816 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X817 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X818 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X819 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X821 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X822 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X823 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X824 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X825 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X826 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X828 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X829 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R70 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X830 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X831 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X832 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X833 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X834 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R71 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X835 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X836 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X837 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X838 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X839 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X842 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X843 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X844 SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X845 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X847 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X848 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X849 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X850 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X852 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X853 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X854 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X855 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X858 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X859 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X862 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X864 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X865 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X866 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X867 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X868 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X870 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X872 VGND SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X873 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X874 VPWR SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X875 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X876 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X877 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X878 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R72 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X879 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X880 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X881 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X883 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X884 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X886 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X887 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R73 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X888 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X889 VGND SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X890 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R74 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X892 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X893 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X894 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X895 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X896 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R75 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X897 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X899 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X901 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X902 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R76 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X903 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X904 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X905 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X906 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X909 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X910 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X911 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X912 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X913 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X914 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R77 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X915 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X917 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X918 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X919 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X920 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X922 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X923 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X924 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X925 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X926 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R78 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X928 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X929 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X930 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X931 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R79 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X932 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X933 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X934 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X935 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X936 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X937 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X939 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X940 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X941 SUNSAR_SAR8B_CV_0.XB1.XA3.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X942 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X944 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X945 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R80 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X946 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X947 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X948 VGND SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X949 SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X950 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X951 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X952 TIE_L SUNSAR_CAPT8B_CV_0.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X953 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X954 SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X955 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X957 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R81 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X958 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X959 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X961 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X962 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X963 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X964 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X965 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X967 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X970 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X971 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X972 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X974 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X975 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X976 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R82 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X977 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X978 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X980 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X982 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X983 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X984 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X985 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X986 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X987 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X988 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R83 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X991 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X993 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X994 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X995 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X997 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R84 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X999 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1000 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1001 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1002 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1004 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1005 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1008 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1013 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1014 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R85 uio_out[0] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X1016 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1018 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1019 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1020 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1021 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1022 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1023 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1024 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1025 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1029 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1030 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1033 VGND SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1034 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1035 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1036 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1037 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 VPWR uo_out[7] 1.27659f
C1 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.204048f
C3 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.316693f
C4 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.142061f
C5 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR 0.106927f
C6 a_15210_34716# VPWR 0.399819f
C7 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_4390# 0.15559f
C8 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C9 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D VPWR 0.108436f
C10 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C11 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.26479f
C12 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38576f
C13 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C14 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.301485f
C15 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y uo_out[6] 0.306905f
C16 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR 0.106927f
C17 a_15210_31196# VPWR 0.44007f
C18 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.649845f
C19 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.179089f
C20 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C21 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C22 a_3782_40296# VPWR 0.457343f
C23 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[6] 0.258218f
C24 SUNSAR_CAPT8B_CV_0.XE10.QN VPWR 0.901622f
C25 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.375196f
C26 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR 0.722887f
C27 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.55251f
C28 SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR 2.64054f
C29 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y a_16382_42408# 0.113479f
C30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.702226f
C31 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.126806f
C32 SUNSAR_SAR8B_CV_0.D<3> VPWR 5.17056f
C33 a_13842_34716# VPWR 0.399819f
C34 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233744f
C35 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C36 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VPWR 0.279205f
C37 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.669708f
C38 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.379175p
C39 a_16542_5974# VPWR 0.449888f
C40 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR 2.95305f
C41 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR 0.930839f
C42 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.635098f
C43 a_13842_31196# VPWR 0.44007f
C44 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C45 SUNSAR_CAPT8B_CV_0.XD09.QN VPWR 0.901622f
C46 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.220689f
C47 SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D VPWR 0.101979f
C48 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR 2.7271f
C49 a_5150_41880# VPWR 0.395781f
C50 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C51 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.15651f
C52 a_3782_44168# VPWR 0.3405f
C53 SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR 1.63909f
C54 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.CKN 0.102131f
C55 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C56 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3686# 0.16579f
C57 a_23942_44344# VPWR 0.342053f
C58 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VPWR 1.77562f
C59 a_5130_27852# VPWR 0.358413f
C60 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C61 a_23942_40648# VPWR 0.489094f
C62 SUNSAR_CAPT8B_CV_0.XB07.QN uo_out[7] 0.263255f
C63 SUNSAR_CAPT8B_CV_0.XC08.QN VPWR 0.901622f
C64 SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D VPWR 0.119314f
C65 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR 2.72582f
C66 a_3782_41880# VPWR 0.395781f
C67 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.63636f
C68 a_20250_28908# VPWR 0.395394f
C69 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C70 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.2165f
C71 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.702226f
C72 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.255261f
C73 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.363295f
C74 SUNSAR_SAR8B_CV_0.XA6.ENO a_17730_28556# 0.132757f
C75 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.318734f
C76 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D VPWR 0.104609f
C77 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.143148f
C78 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C79 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.57155f
C80 SUNSAR_CAPT8B_CV_0.XE10.XA4.A a_10190_42760# 0.111734f
C81 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y a_5150_41880# 0.100592f
C82 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR 0.808658f
C83 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_2768# 0.172147f
C84 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR 0.106927f
C85 SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR 1.2202f
C86 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.55251f
C87 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.241356f
C88 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.178114f
C89 a_3762_27852# VPWR 0.358599f
C90 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C91 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_2928# 0.105547f
C92 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.59087f
C93 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C94 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.29297f
C95 SUNSAR_CAPT8B_CV_0.XB07.QN VPWR 0.901622f
C96 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.383512f
C97 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR 0.725614f
C98 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR 2.72889f
C99 a_18882_28908# VPWR 0.395394f
C100 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C101 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.327909f
C102 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.380687f
C103 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.267238f
C104 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.204048f
C105 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43816# 0.129239f
C106 SUNSAR_SAR8B_CV_0.D<4> VPWR 5.15123f
C107 a_10170_34716# VPWR 0.399819f
C108 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.M3.G 0.151329f
C109 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.07223f
C110 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.164325f
C111 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.440586f
C112 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y uo_out[7] 0.308722f
C113 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR 0.93081f
C114 a_10170_31196# VPWR 0.44007f
C115 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.393076f
C116 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C117 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C118 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.2622f
C119 SUNSAR_CAPT8B_CV_0.XA2.MN0.G VPWR 0.667429f
C120 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR 0.722887f
C121 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 3.55251f
C122 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D VPWR 0.118162f
C123 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35420# 0.160931f
C124 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.09966f
C125 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C126 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y a_12710_42408# 0.111909f
C127 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.702226f
C128 SUNSAR_SAR8B_CV_0.XA5.ENO a_16362_28556# 0.135353f
C129 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D 0.109021f
C130 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR 0.106927f
C131 a_8802_34716# VPWR 0.399819f
C132 SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR 1.63909f
C133 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.ENO 0.409858f
C134 a_9990_5622# VPWR 0.470814f
C135 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y uo_out[7] 0.248979f
C136 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VPWR 1.77562f
C137 SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR 1.22023f
C138 a_8802_31196# VPWR 0.44007f
C139 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 0.595738f
C140 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C141 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.88588f
C142 a_20250_33836# VPWR 0.407174f
C143 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VPWR 1.20019f
C144 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.126085f
C145 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_5130_35420# 0.133834f
C146 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C147 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.17528f
C148 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C149 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR 0.106927f
C150 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C151 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C152 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.41635f
C153 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR 2.9531f
C154 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.649845f
C155 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.179089f
C156 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.746324f
C157 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.431984f
C158 a_20270_44168# VPWR 0.340085f
C159 a_20270_40648# VPWR 0.492579f
C160 a_18882_33836# VPWR 0.409601f
C161 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA8.A 0.527529f
C162 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.233892f
C163 a_15210_28908# VPWR 0.395394f
C164 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C165 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.297363f
C166 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y a_11342_42408# 0.113479f
C167 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.11382f
C168 a_16542_2630# VPWR 0.448659f
C169 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.702226f
C170 SUNSAR_SAR8B_CV_0.D<5> VPWR 5.14531f
C171 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.M3.G 0.1501f
C172 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VPWR 0.271482f
C173 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C174 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_4038# 0.135393f
C175 SUNSAR_CAPT8B_CV_0.XD09.XA4.A a_8822_42760# 0.113305f
C176 a_9990_5974# VPWR 0.451043f
C177 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR 0.765792f
C178 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR 0.930839f
C179 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.744161f
C180 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.07164f
C181 a_18902_44168# VPWR 0.3405f
C182 a_18902_40648# VPWR 0.491225f
C183 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR 0.106927f
C184 a_13842_28908# VPWR 0.395394f
C185 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.19724f
C186 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C187 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.419738f
C188 a_5130_34716# VPWR 0.399819f
C189 SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR 1.63909f
C190 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C191 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y a_17750_42408# 0.100131f
C192 a_23922_26796# VPWR 0.442318f
C193 a_5130_31196# VPWR 0.44007f
C194 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_ON 2.96993f
C195 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 54.2173f
C196 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR 0.106927f
C197 SUNSAR_SAR8B_CV_0.SARN ua[0] 1.02347f
C198 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_3762_35420# 0.133834f
C199 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80606f
C200 TIE_L1 uo_out[5] 0.366299f
C201 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C202 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.702226f
C203 a_8822_44168# VPWR 0.3405f
C204 SUNSAR_SAR8B_CV_0.XA4.ENO a_12690_28556# 0.132757f
C205 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP 0.596437f
C206 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.318734f
C207 a_3762_34716# VPWR 0.399819f
C208 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D VPWR 0.104609f
C209 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.ENO 0.438277f
C210 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.174845f
C211 a_20270_43816# VPWR 0.391817f
C212 SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR 1.2202f
C213 a_3762_31196# VPWR 0.44007f
C214 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.178114f
C215 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.625035f
C216 SUNSAR_SAR8B_CV_0.SARN ua[1] 0.806872f
C217 a_15210_33836# VPWR 0.409601f
C218 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35420# 0.160931f
C219 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.665724f
C220 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C221 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.419738f
C222 SUNSAR_SAR8B_CV_0.D<6> VPWR 5.17441f
C223 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VPWR 0.271482f
C224 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.587991f
C225 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.EN 0.343905f
C226 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.250503f
C227 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.ENO 0.116058f
C228 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR 0.93081f
C229 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.39306f
C230 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C231 a_15230_44168# VPWR 0.340085f
C232 a_15230_40648# VPWR 0.492579f
C233 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.375196f
C234 a_13842_33836# VPWR 0.409601f
C235 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.55251f
C236 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.63636f
C237 a_10170_28908# VPWR 0.395394f
C238 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y a_7670_42408# 0.111909f
C239 TIE_L1 uo_out[7] 0.461734f
C240 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.74594f
C241 SUNSAR_SAR8B_CV_0.XA3.ENO a_11322_28556# 0.135353f
C242 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR 0.106927f
C243 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR 3.91346f
C244 SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR 1.63909f
C245 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_4742# 0.156331f
C246 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.55251f
C247 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.CKN 0.41624f
C248 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.ENO 0.111173f
C249 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.849501f
C250 a_20250_26796# VPWR 0.441753f
C251 a_21402_36828# SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.104051f
C252 SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR 1.22023f
C253 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR 6.94539f
C254 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA2.Y 0.241356f
C255 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.419738f
C256 a_13862_44168# VPWR 0.3405f
C257 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.294852f
C258 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR 0.106927f
C259 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA8.A 0.527529f
C260 a_8802_28908# VPWR 0.395394f
C261 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.34383f
C262 a_9990_2630# VPWR 0.447504f
C263 TIE_L1 VPWR 0.115195f
C264 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.86675f
C265 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.204048f
C266 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR 0.106927f
C267 a_23922_34892# VPWR 0.395601f
C268 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_4742# 0.156331f
C269 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C270 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_2768# 0.172147f
C271 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D 0.101001f
C272 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.134182f
C273 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.ENO 0.111217f
C274 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.ENO 0.893904f
C275 a_18882_26796# VPWR 0.442908f
C276 a_23922_31724# VPWR 0.412398f
C277 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.179089f
C278 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.419738f
C279 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.26537f
C280 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 6.86675f
C281 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR 0.106927f
C282 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.39041f
C283 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C284 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y a_6302_42408# 0.113479f
C285 a_16542_2982# VPWR 0.490338f
C286 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C287 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.748719f
C288 SUNSAR_SAR8B_CV_0.D<7> VPWR 3.61291f
C289 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D VPWR 0.104609f
C290 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C291 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.ENO 0.503825f
C292 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.ENO 0.952619f
C293 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.ENO 0.111173f
C294 SUNSAR_CAPT8B_CV_0.XC08.XA4.A a_5150_42760# 0.111734f
C295 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.310451f
C296 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR 0.930839f
C297 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.744161f
C298 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO 0.144331f
C299 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.419738f
C300 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 0.625175f
C301 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.268769f
C302 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.383512f
C303 a_10170_33836# VPWR 0.409601f
C304 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.352238f
C305 SUNSAR_SAR8B_CV_0.XA7.ENO VPWR 4.77251f
C306 SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR 1.63909f
C307 SUNSAR_CAPT8B_CV_0.XA4.MN0.S SUNSAR_CAPT8B_CV_0.XA4.Y 0.206292f
C308 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.ENO 1.02916f
C309 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.ENO 0.111217f
C310 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.426291f
C311 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.449584f
C312 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.15234f
C313 SUNSAR_SAR8B_CV_0.XA4.CEO VPWR 2.30385f
C314 SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR 2.62711f
C315 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.649845f
C316 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.419738f
C317 SUNSAR_SAR8B_CV_0.XA2.XA10.Y a_7650_36300# 0.13253f
C318 a_8802_33836# VPWR 0.409601f
C319 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.2165f
C320 a_5130_28908# VPWR 0.395394f
C321 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.165965f
C322 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.136678f
C323 SUNSAR_SAR8B_CV_0.XB2.XA3.B ua[0] 0.241597f
C324 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C325 SUNSAR_SAR8B_CV_0.XA2.ENO a_7650_28556# 0.132757f
C326 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C327 a_23942_41880# VPWR 0.398828f
C328 SUNSAR_SAR8B_CV_0.XA6.ENO VPWR 5.54203f
C329 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN 0.143148f
C330 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.ENO 0.952619f
C331 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.ENO 0.111173f
C332 a_15210_26796# VPWR 0.441753f
C333 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.340491f
C334 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR 0.720133f
C335 SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR 1.2202f
C336 SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR 2.62329f
C337 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.178114f
C338 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP 0.435464f
C339 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D 0.252966f
C340 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR 0.106927f
C341 a_3762_28908# VPWR 0.395394f
C342 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189112f
C343 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.52234f
C344 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S ua[0] 0.100365f
C345 SUNSAR_CAPT8B_CV_0.XA4.Y clk 0.206733f
C346 SUNSAR_SAR8B_CV_0.XA5.ENO VPWR 4.84607f
C347 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_3728# 0.172147f
C348 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.62595f
C349 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.ENO 1.02916f
C350 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.ENO 0.111217f
C351 a_13842_26796# VPWR 0.442908f
C352 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.449584f
C353 SUNSAR_SAR8B_CV_0.XA3.CEO VPWR 1.06031f
C354 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR 0.93081f
C355 SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR 2.62342f
C356 SUNSAR_SAR8B_CV_0.XA1.XA10.Y a_6282_36300# 0.13402f
C357 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.137975f
C358 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 27.1625f
C359 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR 0.106927f
C360 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y a_2630_42408# 0.111909f
C361 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.SARN 0.108405f
C362 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C363 SUNSAR_SAR8B_CV_0.XA1.ENO a_6282_28556# 0.135353f
C364 SUNSAR_SAR8B_CV_0.XA4.ENO VPWR 5.52623f
C365 SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR 1.63909f
C366 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VPWR 0.271482f
C367 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.55251f
C368 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.ENO 0.438277f
C369 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.CKN 0.200119f
C370 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.ENO 0.952619f
C371 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.ENO 0.111173f
C372 SUNSAR_CAPT8B_CV_0.XB07.XA4.A a_3782_42760# 0.113305f
C373 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARP 0.506551f
C374 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR 0.723762f
C375 SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR 1.22398f
C376 SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR 2.62342f
C377 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.241356f
C378 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.625035f
C379 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.276413f
C380 a_5130_33836# VPWR 0.409601f
C381 a_9990_2982# VPWR 0.491909f
C382 SUNSAR_SAR8B_CV_0.XB1.XA3.B ua[1] 0.241597f
C383 a_20270_41880# VPWR 0.395781f
C384 SUNSAR_SAR8B_CV_0.XA3.ENO VPWR 4.84607f
C385 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_6768# 0.105547f
C386 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D 0.101001f
C387 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.ENO 1.04628f
C388 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.12241f
C389 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6519f
C390 a_17730_36828# SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.10248f
C391 SUNSAR_SAR8B_CV_0.XA2.CEO VPWR 2.30393f
C392 SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR 2.62342f
C393 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.393125f
C394 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35068# 0.129098f
C395 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO 0.144331f
C396 a_3762_33836# VPWR 0.409601f
C397 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.127551f
C398 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.86675f
C399 SUNSAR_SAR8B_CV_0.XB1.TIE_L ua[0] 1.05246f
C400 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA8.A 0.527529f
C401 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D VPWR 0.104609f
C402 a_16542_3334# VPWR 0.380282f
C403 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S ua[1] 0.100365f
C404 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.107567f
C405 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA10.Y 0.303978f
C406 SUNSAR_SAR8B_CV_0.XA2.ENO VPWR 5.52623f
C407 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D VPWR 0.104609f
C408 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.CKN 0.41624f
C409 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.432466f
C410 a_10170_26796# VPWR 0.441753f
C411 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR 0.720114f
C412 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 6.86675f
C413 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR 0.94014f
C414 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR 2.62393f
C415 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_4688# 0.172147f
C416 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.449584f
C417 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.105016f
C418 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D 0.152518f
C419 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR 0.106927f
C420 SUNSAR_SAR8B_CV_0.XB1.TIE_L ua[1] 0.704356f
C421 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.109613f
C422 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.13078f
C423 SUNSAR_SAR8B_CV_0.XA1.ENO VPWR 4.84607f
C424 SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR 1.63909f
C425 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_5094# 0.160184f
C426 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_4688# 0.172147f
C427 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VPWR 0.271482f
C428 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 0.250503f
C429 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y a_12710_42408# 0.100131f
C430 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.55251f
C431 a_8802_26796# VPWR 0.442908f
C432 SUNSAR_SAR8B_CV_0.XA1.CEO VPWR 1.0603f
C433 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.11641f
C434 a_23922_35948# VPWR 0.390687f
C435 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR 2.62403f
C436 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.649845f
C437 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.449584f
C438 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.671839f
C439 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.284482f
C440 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.375025f
C441 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 13.6523f
C442 SUNSAR_SAR8B_CV_0.SARN VPWR 0.132799f
C443 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR 0.106927f
C444 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D VPWR 0.104609f
C445 SUNSAR_SAR8B_CV_0.XA0.ENO a_2610_28556# 0.132757f
C446 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.131536f
C447 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.109137f
C448 SUNSAR_SAR8B_CV_0.XA0.ENO VPWR 5.52718f
C449 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_5094# 0.160184f
C450 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.ENO 0.503825f
C451 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.104933f
C452 a_16362_36828# SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.104051f
C453 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR 0.728492f
C454 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.152052f
C455 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.143675f
C456 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.744161f
C457 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO 0.144331f
C458 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.449584f
C459 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 0.625175f
C460 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D 0.150467f
C461 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.10225f
C462 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.227625f
C463 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.16676f
C464 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C465 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.352238f
C466 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 1.62434f
C467 SUNSAR_SAR8B_CV_0.XA0.CEO VPWR 2.30575f
C468 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.339883f
C469 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.180903f
C470 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.144778f
C471 a_20250_32076# VPWR 0.433941f
C472 a_20250_28204# VPWR 0.361706f
C473 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.11099f
C474 SUNSAR_SAR8B_CV_0.XA0.XA10.Y a_2610_36300# 0.13253f
C475 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.372599f
C476 a_23942_42408# VPWR 0.3915f
C477 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1615f
C478 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C479 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.45828f
C480 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.143023f
C481 a_20250_35068# VPWR 0.391458f
C482 SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR 1.63909f
C483 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D VPWR 0.104609f
C484 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.432466f
C485 a_5130_26796# VPWR 0.441753f
C486 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.139471f
C487 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 27.1615f
C488 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_6608# 0.172147f
C489 a_20250_35948# VPWR 0.414756f
C490 a_18882_32076# VPWR 0.436368f
C491 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 4.28648f
C492 a_18882_28204# VPWR 0.36179f
C493 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35068# 0.127528f
C494 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_5648# 0.172147f
C495 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.180455f
C496 TIE_L clk 0.150303f
C497 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VPWR 0.405511f
C498 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA8.A 0.527529f
C499 SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D VPWR 0.101979f
C500 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.109613f
C501 a_9990_3334# VPWR 0.380282f
C502 a_18882_35068# VPWR 0.394528f
C503 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_5648# 0.172147f
C504 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.M3.G 0.224309f
C505 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.12241f
C506 a_3762_26796# VPWR 0.442908f
C507 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 54.2165f
C508 a_20250_37180# VPWR 0.469114f
C509 a_18882_35948# VPWR 0.417826f
C510 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.252047f
C511 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.791379f
C512 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D 0.104122f
C513 TIE_L uo_out[0] 0.280844f
C514 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.449584f
C515 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 3.57448f
C516 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR 1.70987f
C517 SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D VPWR 0.119314f
C518 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.155424f
C519 a_21422_41000# SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.115667f
C520 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.110962f
C521 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.142977f
C522 SUNSAR_CAPT8B_CV_0.XA4.Y VPWR 1.18734f
C523 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.ENO 0.434116f
C524 a_18882_37180# VPWR 0.473682f
C525 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.154232f
C526 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.63636f
C527 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.08082f
C528 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.11884f
C529 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D 0.155821f
C530 TIE_L uo_out[1] 0.50141f
C531 a_20270_42408# VPWR 0.391292f
C532 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR 0.725614f
C533 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D VPWR 0.104609f
C534 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.CEO 0.301665f
C535 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C536 a_20270_41000# SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.156079f
C537 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.175642f
C538 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.133602f
C539 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.M3.G 0.263588f
C540 a_23922_27148# VPWR 0.483246f
C541 a_12690_36828# SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.10248f
C542 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.3401f
C543 a_15210_32076# VPWR 0.436368f
C544 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO 0.144331f
C545 a_15210_28204# VPWR 0.361706f
C546 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C547 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON a_20250_30316# 0.127528f
C548 TIE_L uo_out[2] 0.162449f
C549 a_18902_42408# VPWR 0.391292f
C550 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6519f
C551 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR 0.722887f
C552 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.227625f
C553 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR 1.56028f
C554 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C555 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.142956f
C556 a_15210_35068# VPWR 0.394528f
C557 a_20270_43288# VPWR 0.394205f
C558 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_5446# 0.102604f
C559 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VPWR 0.271482f
C560 a_15210_35948# VPWR 0.417826f
C561 a_13842_32076# VPWR 0.436368f
C562 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.744161f
C563 a_13842_28204# VPWR 0.36179f
C564 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_6608# 0.172147f
C565 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C566 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03123f
C567 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.276413f
C568 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D 0.150467f
C569 TIE_L uo_out[3] 0.188109f
C570 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR 4.36162f
C571 SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D VPWR 0.101979f
C572 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR 0.183853f
C573 a_12710_41000# SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.114097f
C574 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.133602f
C575 a_13842_35068# VPWR 0.394528f
C576 a_18902_43288# VPWR 0.394205f
C577 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_5446# 0.101033f
C578 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_2928# 0.105547f
C579 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.12241f
C580 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.ENO 0.793076f
C581 a_15210_37180# VPWR 0.474036f
C582 a_13842_35948# VPWR 0.417826f
C583 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.649845f
C584 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35068# 0.129098f
C585 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_3888# 0.105547f
C586 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.199516f
C587 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C588 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON a_18882_30316# 0.129098f
C589 TIE_L uo_out[4] 0.333172f
C590 a_23922_34540# VPWR 0.502044f
C591 SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D VPWR 0.119314f
C592 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D VPWR 0.104609f
C593 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR 1.5612f
C594 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.142977f
C595 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D VPWR 0.104609f
C596 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.CKN 0.200119f
C597 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.ENO 0.491653f
C598 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.432466f
C599 a_20250_27148# VPWR 0.470364f
C600 a_13842_37180# VPWR 0.473697f
C601 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6519f
C602 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO 0.144331f
C603 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.233892f
C604 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.20727f
C605 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C606 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C607 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03123f
C608 TIE_L uo_out[5] 1.32477f
C609 a_15230_42408# VPWR 0.391292f
C610 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR 0.728421f
C611 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.227625f
C612 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.545186f
C613 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR 0.183853f
C614 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.189429f
C615 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.133602f
C616 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VPWR 0.271482f
C617 a_18882_27148# VPWR 0.471462f
C618 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.290432f
C619 a_10170_32076# VPWR 0.436368f
C620 a_10170_28204# VPWR 0.361706f
C621 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.CKN 0.153964f
C622 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.215251f
C623 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C624 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.377598f
C625 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.284482f
C626 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D 0.104122f
C627 TIE_L uo_out[6] 0.203535f
C628 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C629 a_13862_42408# VPWR 0.391292f
C630 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.55251f
C631 SUNSAR_SAR8B_CV_0.XB1.TIE_L VPWR 7.37316f
C632 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA8.A 0.527529f
C633 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARN 0.64474f
C634 a_16542_4038# VPWR 0.379979f
C635 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.11826f
C636 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.191868f
C637 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.142956f
C638 a_10170_35068# VPWR 0.394528f
C639 a_15230_43288# VPWR 0.394205f
C640 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.146492f
C641 a_10170_35948# VPWR 0.417826f
C642 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.182595f
C643 a_8802_32076# VPWR 0.436368f
C644 a_8802_28204# VPWR 0.36179f
C645 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.178111f
C646 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03107f
C647 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D 0.155821f
C648 TIE_L uo_out[7] 0.462706f
C649 a_18902_41000# SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.15757f
C650 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.137745f
C651 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.175642f
C652 a_11342_41000# SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.115667f
C653 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.133602f
C654 SUNSAR_SAR8B_CV_0.XA20.XA2.CO a_23922_30844# 0.100515f
C655 a_13862_43288# VPWR 0.394205f
C656 a_8802_35068# VPWR 0.394528f
C657 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_3888# 0.105547f
C658 SUNSAR_CAPT8B_CV_0.XA4.MN0.S SUNSAR_CAPT8B_CV_0.XA3.Y 0.300065f
C659 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.ENO 1.2771f
C660 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y a_7670_42408# 0.100131f
C661 a_10170_37180# VPWR 0.474068f
C662 a_8802_35948# VPWR 0.417826f
C663 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_4848# 0.105547f
C664 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.50324f
C665 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.293159f
C666 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON a_15210_30316# 0.127528f
C667 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.474658f
C668 TIE_L VPWR 0.401306f
C669 a_20250_36828# VPWR 0.392512f
C670 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.412143f
C671 a_17750_41000# SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.114097f
C672 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.4271f
C673 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C674 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.162703f
C675 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C676 SUNSAR_SAR8B_CV_0.XB2.M3.G ua[0] 0.765539f
C677 a_10190_41000# SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.156079f
C678 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.142977f
C679 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D VPWR 0.104609f
C680 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.ENO 0.11341f
C681 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y 0.22339f
C682 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.432466f
C683 a_15210_27148# VPWR 0.470364f
C684 a_8802_37180# VPWR 0.473729f
C685 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.152052f
C686 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.324105f
C687 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.321724f
C688 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.63636f
C689 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35068# 0.127528f
C690 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C691 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.791351f
C692 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.CEO 0.432008f
C693 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D 0.150467f
C694 a_10190_42408# VPWR 0.391292f
C695 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR 0.112098f
C696 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D VPWR 0.104609f
C697 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.133602f
C698 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.M3.G 0.224309f
C699 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.12241f
C700 a_13842_27148# VPWR 0.471462f
C701 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.339883f
C702 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.37807f
C703 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.CEO 0.138f
C704 a_5130_32076# VPWR 0.436368f
C705 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO 0.144331f
C706 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.146458f
C707 a_5130_28204# VPWR 0.361706f
C708 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.228326f
C709 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.158152f
C710 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON a_13842_30316# 0.129098f
C711 a_8822_42408# VPWR 0.391292f
C712 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR 0.112858f
C713 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.55251f
C714 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.227625f
C715 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.142956f
C716 a_10190_43288# VPWR 0.394205f
C717 a_5130_35068# VPWR 0.394528f
C718 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C719 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.267144f
C720 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.724217f
C721 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_5808# 0.105547f
C722 a_5130_35948# VPWR 0.417826f
C723 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.158152f
C724 SUNSAR_SAR8B_CV_0.DONE ui_in[0] 0.175856f
C725 a_3762_32076# VPWR 0.436368f
C726 a_3762_28204# VPWR 0.36179f
C727 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C728 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.CKN 0.153964f
C729 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR 4.24834f
C730 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA8.A 0.527529f
C731 a_18882_36828# VPWR 0.395703f
C732 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C733 a_9990_4038# VPWR 0.379979f
C734 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.133602f
C735 a_8822_43288# VPWR 0.394205f
C736 a_3762_35068# VPWR 0.394528f
C737 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_4848# 0.105547f
C738 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.ENO 1.2771f
C739 a_5130_37180# VPWR 0.474051f
C740 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.386137f
C741 a_3762_35948# VPWR 0.417826f
C742 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_5808# 0.105547f
C743 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<0> 0.492001f
C744 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C745 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1615f
C746 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.220689f
C747 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D 0.104122f
C748 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.145483f
C749 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.205884f
C750 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D VPWR 0.104609f
C751 a_16382_41000# SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.115667f
C752 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.238636f
C753 SUNSAR_SAR8B_CV_0.XB1.M3.G ua[1] 0.762388f
C754 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR 2.50821f
C755 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.142977f
C756 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VPWR 0.271482f
C757 a_10170_27148# VPWR 0.470364f
C758 a_3762_37180# VPWR 0.473713f
C759 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.154232f
C760 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.722427f
C761 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.220689f
C762 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C763 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR 0.618979f
C764 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO 0.144331f
C765 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VPWR 0.429492f
C766 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C767 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.791379f
C768 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.10132f
C769 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.112859f
C770 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D 0.155821f
C771 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.276413f
C772 a_5150_42408# VPWR 0.391292f
C773 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.694484f
C774 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.227625f
C775 a_15230_41000# SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.156079f
C776 SUNSAR_SAR8B_CV_0.XB2.CKN VPWR 2.34497f
C777 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.133602f
C778 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.12241f
C779 a_8802_27148# VPWR 0.471462f
C780 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.3401f
C781 SUNSAR_SAR8B_CV_0.XA20.XA10.B VPWR 1.13456f
C782 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR 0.324111f
C783 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR 0.137646f
C784 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.143554f
C785 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35068# 0.129098f
C786 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.55251f
C787 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.228332f
C788 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.34399f
C789 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.11263f
C790 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.377598f
C791 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON a_10170_30316# 0.127528f
C792 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.145483f
C793 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR 4.25569f
C794 a_3782_42408# VPWR 0.391292f
C795 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.2165f
C796 SUNSAR_SAR8B_CV_0.SARP ua[1] 1.01251f
C797 a_15210_36828# VPWR 0.395582f
C798 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31666f
C799 a_8822_41000# SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.15757f
C800 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C801 a_5150_43288# VPWR 0.394205f
C802 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR 2.1352f
C803 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C804 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.393665f
C805 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.200058f
C806 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.432466f
C807 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.103734f
C808 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.722417f
C809 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_6768# 0.105547f
C810 SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR 0.774301f
C811 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.377598f
C812 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR 2.30036f
C813 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VPWR 1.06002f
C814 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<1> 0.297507f
C815 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.193518f
C816 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.209352f
C817 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.112859f
C818 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D 0.150467f
C819 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.204048f
C820 a_13842_36828# VPWR 0.395703f
C821 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.111867f
C822 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_34540# 0.103065f
C823 a_7670_41000# SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.114097f
C824 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.133602f
C825 a_3782_43288# VPWR 0.394205f
C826 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y uo_out[0] 0.245915f
C827 SUNSAR_SAR8B_CV_0.XA6.DONE VPWR 0.246222f
C828 a_20250_30316# VPWR 0.403745f
C829 a_22790_41880# SUNSAR_CAPT8B_CV_0.XA4.Y 0.111538f
C830 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.241356f
C831 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.EN 0.176398f
C832 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.ENO 1.2771f
C833 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO 1.43919f
C834 a_20250_37532# VPWR 0.454392f
C835 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.107427f
C836 SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR 0.780003f
C837 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR 2.31184f
C838 a_10190_41000# VPWR 0.388175f
C839 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR 0.138148f
C840 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.11263f
C841 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.238862f
C842 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.293159f
C843 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.284482f
C844 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON a_8802_30316# 0.129098f
C845 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.145483f
C846 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR 0.686731f
C847 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.205884f
C848 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y uo_out[0] 0.307374f
C849 SUNSAR_SAR8B_CV_0.XA5.DONE VPWR 0.245452f
C850 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C851 a_18882_30316# VPWR 0.403802f
C852 a_5130_27148# VPWR 0.470364f
C853 a_18882_37532# VPWR 0.458267f
C854 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.722427f
C855 SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR 0.779986f
C856 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR 2.31184f
C857 a_8822_41000# VPWR 0.388256f
C858 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.63636f
C859 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VPWR 1.06875f
C860 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.112859f
C861 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.372578f
C862 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.437693f
C863 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.CEO 0.432008f
C864 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VPWR 0.898003f
C865 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D VPWR 0.104609f
C866 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.182408f
C867 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.86675f
C868 SUNSAR_SAR8B_CV_0.XA4.DONE VPWR 0.246222f
C869 a_3762_27148# VPWR 0.471462f
C870 SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR 0.780003f
C871 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR 2.31184f
C872 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR 0.137646f
C873 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<2> 0.297715f
C874 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.228326f
C875 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.11263f
C876 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.158152f
C877 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.SARP 0.122781f
C878 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.145483f
C879 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.126354f
C880 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VPWR 0.898003f
C881 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.86675f
C882 a_10170_36828# VPWR 0.396003f
C883 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.301485f
C884 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.291229f
C885 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.227625f
C886 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C887 SUNSAR_SAR8B_CV_0.XB1.CKN VPWR 2.34497f
C888 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.SARP 0.147435f
C889 SUNSAR_CAPT8B_CV_0.XA3.Y VPWR 0.86364f
C890 SUNSAR_SAR8B_CV_0.XA3.DONE VPWR 0.245452f
C891 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G 0.22339f
C892 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.432466f
C893 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.722417f
C894 SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR 0.779986f
C895 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR 2.31184f
C896 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.145738f
C897 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35068# 0.127528f
C898 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.441867f
C899 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VPWR 1.05322f
C900 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.437693f
C901 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.242472f
C902 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.2165f
C903 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN 0.253395f
C904 TIE_L TIE_L1 0.284231f
C905 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.318734f
C906 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VPWR 0.898003f
C907 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR 0.112858f
C908 a_8802_36828# VPWR 0.396052f
C909 a_13862_41000# SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.15757f
C910 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.11536f
C911 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR 2.50821f
C912 a_6302_41000# SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.115667f
C913 TIE_L2 uo_out[7] 0.106093f
C914 a_23942_43640# VPWR 0.412992f
C915 SUNSAR_SAR8B_CV_0.XA2.DONE VPWR 0.246222f
C916 a_15210_30316# VPWR 0.404384f
C917 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y a_2630_42408# 0.100131f
C918 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.12241f
C919 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C920 a_15210_37532# VPWR 0.459479f
C921 a_17750_43816# SUNSAR_CAPT8B_CV_0.XH13.QN 0.127669f
C922 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.386137f
C923 SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR 0.780003f
C924 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR 2.31184f
C925 a_5150_41000# VPWR 0.388161f
C926 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR 0.138148f
C927 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.437693f
C928 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C929 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.145483f
C930 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON a_5130_30316# 0.127528f
C931 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR 0.112858f
C932 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VPWR 0.898003f
C933 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.205884f
C934 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D VPWR 0.104609f
C935 SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR 0.665006f
C936 a_5150_41000# SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.156079f
C937 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP 0.123668f
C938 TIE_L2 VPWR 0.106973f
C939 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y uo_out[1] 0.305961f
C940 SUNSAR_SAR8B_CV_0.XA1.DONE VPWR 0.245452f
C941 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C942 SUNSAR_SAR8B_CV_0.XA7.XA10.Y a_21402_36300# 0.13402f
C943 a_13842_30316# VPWR 0.404384f
C944 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA1.CEO 0.303978f
C945 a_20250_27500# VPWR 0.382397f
C946 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.738812f
C947 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.152052f
C948 a_13842_37532# VPWR 0.458324f
C949 SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR 0.779986f
C950 SUNSAR_SAR8B_CV_0.DONE VPWR 7.82595f
C951 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR 2.31184f
C952 a_3782_41000# VPWR 0.388256f
C953 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35420# 0.160931f
C954 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.233892f
C955 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.441867f
C956 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VPWR 1.06875f
C957 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<3> 0.297504f
C958 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.437693f
C959 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.791351f
C960 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.297144f
C961 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR 4.2492f
C962 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VPWR 0.898003f
C963 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.227625f
C964 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23942_42760# 0.101843f
C965 a_16542_4566# VPWR 0.413433f
C966 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y uo_out[1] 0.248461f
C967 SUNSAR_SAR8B_CV_0.XA0.DONE VPWR 0.247527f
C968 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.CEO 0.13078f
C969 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.241356f
C970 a_18882_27500# VPWR 0.382189f
C971 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.280191f
C972 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.339883f
C973 a_16382_43816# SUNSAR_CAPT8B_CV_0.XG12.QN 0.129239f
C974 SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR 0.784656f
C975 a_23942_41000# VPWR 0.390551f
C976 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR 2.31184f
C977 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.143554f
C978 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_20250_35420# 0.133834f
C979 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR 0.137646f
C980 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.228332f
C981 a_18902_43816# VPWR 0.391817f
C982 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON a_3762_30316# 0.129098f
C983 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.204048f
C984 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.145483f
C985 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VPWR 0.898003f
C986 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 27.1615f
C987 a_5130_36828# VPWR 0.395767f
C988 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22790_42760# 0.13379f
C989 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.301485f
C990 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR 0.106927f
C991 a_23922_35420# VPWR 0.416528f
C992 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C993 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.393049f
C994 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.738798f
C995 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.152045f
C996 a_23922_36300# VPWR 0.472384f
C997 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR 4.6743f
C998 a_23942_41352# VPWR 0.376408f
C999 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VPWR 1.05322f
C1000 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.331207f
C1001 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.276252f
C1002 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VPWR 0.898003f
C1003 a_3762_36828# VPWR 0.395857f
C1004 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.254583f
C1005 SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR 0.665006f
C1006 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.464697f
C1007 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.159359f
C1008 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR 2.95296f
C1009 a_10170_30316# VPWR 0.404384f
C1010 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA0.CEO 0.352238f
C1011 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.12241f
C1012 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C1013 a_10170_37532# VPWR 0.459599f
C1014 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6519f
C1015 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.107427f
C1016 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35068# 0.129098f
C1017 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR 0.138148f
C1018 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<4> 0.297602f
C1019 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C1020 ua[1] ua[0] 3.85017f
C1021 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.145483f
C1022 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR 4.27988f
C1023 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VPWR 0.898003f
C1024 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.205884f
C1025 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.42393f
C1026 SUNSAR_SAR8B_CV_0.EN a_20250_29612# 0.142592f
C1027 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VPWR 1.77563f
C1028 a_8802_30316# VPWR 0.404384f
C1029 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.CK 1.59176f
C1030 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.432466f
C1031 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.649845f
C1032 a_15210_27500# VPWR 0.382397f
C1033 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.740872f
C1034 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.154232f
C1035 a_8802_37532# VPWR 0.458443f
C1036 a_20270_41000# VPWR 0.388156f
C1037 a_20250_32956# VPWR 0.433941f
C1038 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_18882_35420# 0.133834f
C1039 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y 0.342913f
C1040 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.63636f
C1041 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VPWR 1.06875f
C1042 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.108751f
C1043 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 3.86364f
C1044 a_15230_43816# VPWR 0.391817f
C1045 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.318734f
C1046 a_23942_42760# VPWR 0.388156f
C1047 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA10.Y 0.381914f
C1048 SUNSAR_SAR8B_CV_0.SARP VPWR 0.139564f
C1049 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y a_15230_41880# 0.100592f
C1050 a_9990_4566# VPWR 0.413433f
C1051 SUNSAR_SAR8B_CV_0.EN a_18882_29612# 0.143959f
C1052 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.324243f
C1053 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR 0.106927f
C1054 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y uo_out[2] 0.246879f
C1055 a_20250_35420# VPWR 0.39661f
C1056 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.744161f
C1057 a_13842_27500# VPWR 0.382189f
C1058 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C1059 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.3401f
C1060 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.55251f
C1061 a_12710_43816# SUNSAR_CAPT8B_CV_0.XF11.QN 0.127669f
C1062 a_20250_36300# VPWR 0.395776f
C1063 a_18902_41000# VPWR 0.388256f
C1064 a_18882_32956# VPWR 0.436368f
C1065 a_20270_41352# VPWR 0.394053f
C1066 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35420# 0.160931f
C1067 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR 0.137646f
C1068 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.227341f
C1069 a_13862_43816# VPWR 0.391817f
C1070 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.204048f
C1071 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.176792f
C1072 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN 0.538639f
C1073 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6519f
C1074 SUNSAR_SAR8B_CV_0.DONE SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.227625f
C1075 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.301485f
C1076 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.174995f
C1077 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VPWR 0.452478f
C1078 a_3782_41000# SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.15757f
C1079 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1080 a_5150_44168# VPWR 0.340085f
C1081 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR 0.714341f
C1082 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y uo_out[2] 0.305131f
C1083 a_18882_35420# VPWR 0.39968f
C1084 SUNSAR_SAR8B_CV_0.XA6.XA10.Y a_17730_36300# 0.13253f
C1085 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.215804f
C1086 a_18882_36300# VPWR 0.399161f
C1087 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.55251f
C1088 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.145738f
C1089 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_22790_43640# 0.127669f
C1090 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VPWR 1.05322f
C1091 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<5> 0.297941f
C1092 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C1093 SUNSAR_CAPT8B_CV_0.XA4.MN0.S clk 0.438597f
C1094 a_20250_29612# VPWR 0.398044f
C1095 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.475004f
C1096 a_2630_41000# SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.114097f
C1097 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C1098 SUNSAR_SAR8B_CV_0.XA7.CEO VPWR 1.1111f
C1099 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VPWR 1.77562f
C1100 a_5130_30316# VPWR 0.404384f
C1101 a_22790_41000# SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.11811f
C1102 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 1.15994f
C1103 a_5130_37532# VPWR 0.459538f
C1104 a_11342_43816# SUNSAR_CAPT8B_CV_0.XE10.QN 0.129239f
C1105 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[0] 0.247314f
C1106 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR 0.138148f
C1107 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.118161f
C1108 clk ui_in[0] 0.169609f
C1109 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.SARP 0.257526f
C1110 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.30776f
C1111 a_20270_42760# VPWR 0.391454f
C1112 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.205884f
C1113 a_18882_29612# VPWR 0.397362f
C1114 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.232115f
C1115 SUNSAR_SAR8B_CV_0.EN a_15210_29612# 0.143959f
C1116 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1117 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CN1 0.466806f
C1118 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR 0.723713f
C1119 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR 2.95303f
C1120 SUNSAR_SAR8B_CV_0.XA5.XA10.Y a_16362_36300# 0.13402f
C1121 a_3762_30316# VPWR 0.404384f
C1122 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.393063f
C1123 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA6.ENO 0.291697f
C1124 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.432466f
C1125 a_10170_27500# VPWR 0.382397f
C1126 a_3762_37532# VPWR 0.458382f
C1127 a_15230_41000# VPWR 0.388156f
C1128 a_15210_32956# VPWR 0.436368f
C1129 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35068# 0.127528f
C1130 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VPWR 1.06875f
C1131 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C1132 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.13041f
C1133 a_10190_43816# VPWR 0.391817f
C1134 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.128204f
C1135 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.318734f
C1136 a_10190_41352# VPWR 0.394053f
C1137 a_18902_42760# VPWR 0.391454f
C1138 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR 0.112858f
C1139 SUNSAR_CAPT8B_CV_0.XI14.XA4.A a_20270_42760# 0.111734f
C1140 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR 0.519052f
C1141 SUNSAR_SAR8B_CV_0.EN a_13842_29612# 0.143959f
C1142 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C1143 SUNSAR_SAR8B_CV_0.XA6.CEO VPWR 2.28789f
C1144 a_15210_35420# VPWR 0.39968f
C1145 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.241356f
C1146 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.12241f
C1147 a_8802_27500# VPWR 0.382189f
C1148 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 54.2165f
C1149 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C1150 a_15210_36300# VPWR 0.398846f
C1151 a_13862_41000# VPWR 0.388256f
C1152 a_13842_32956# VPWR 0.436368f
C1153 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.143554f
C1154 a_23922_28556# VPWR 0.499441f
C1155 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<6> 0.298165f
C1156 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.227352f
C1157 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.118161f
C1158 a_8822_43816# VPWR 0.391817f
C1159 a_8822_41352# VPWR 0.394053f
C1160 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR 0.112858f
C1161 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA10.Y 0.303978f
C1162 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.55549f
C1163 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.726497f
C1164 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.301485f
C1165 a_16542_4918# VPWR 0.470354f
C1166 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CN1 0.466806f
C1167 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1168 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR 0.720096f
C1169 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR 0.106927f
C1170 a_13842_35420# VPWR 0.39968f
C1171 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y uo_out[3] 0.309657f
C1172 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR 6.88568f
C1173 a_23942_40296# VPWR 0.452344f
C1174 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.118152f
C1175 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.26609f
C1176 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.386305f
C1177 a_13842_36300# VPWR 0.399161f
C1178 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 54.2165f
C1179 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35420# 0.160931f
C1180 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.129613f
C1181 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.363295f
C1182 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR 4.24508f
C1183 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.13078f
C1184 a_15210_29612# VPWR 0.397362f
C1185 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_3334# 0.120042f
C1186 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.SARP 0.102632f
C1187 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C1188 SUNSAR_SAR8B_CV_0.XA5.CEO VPWR 1.0603f
C1189 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR 2.95304f
C1190 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y uo_out[3] 0.249907f
C1191 a_23922_30844# VPWR 0.425847f
C1192 a_11322_36828# SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.104051f
C1193 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.744161f
C1194 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.170578f
C1195 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C1196 a_7670_43816# SUNSAR_CAPT8B_CV_0.XD09.QN 0.127669f
C1197 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_15210_35420# 0.133834f
C1198 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.118226f
C1199 uo_out[1] uo_out[0] 0.366897f
C1200 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 1.62434f
C1201 a_15230_42760# VPWR 0.391454f
C1202 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.205884f
C1203 a_13842_29612# VPWR 0.397362f
C1204 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_3334# 0.113134f
C1205 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR 0.519052f
C1206 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1207 SUNSAR_SAR8B_CV_0.EN a_10170_29612# 0.143959f
C1208 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CN1 0.466806f
C1209 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR 0.723728f
C1210 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VPWR 1.77562f
C1211 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.649845f
C1212 a_5130_27500# VPWR 0.382397f
C1213 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.166192f
C1214 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.152052f
C1215 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.473354f
C1216 a_10170_32956# VPWR 0.436368f
C1217 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.63636f
C1218 a_20250_28556# VPWR 0.406628f
C1219 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.D<7> 0.294651f
C1220 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.530644f
C1221 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 4.0111f
C1222 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.13041f
C1223 a_5150_41352# VPWR 0.394053f
C1224 a_13862_42760# VPWR 0.391454f
C1225 SUNSAR_CAPT8B_CV_0.XH13.XA4.A a_18902_42760# 0.113305f
C1226 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VPWR 0.452478f
C1227 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.504801f
C1228 SUNSAR_SAR8B_CV_0.EN a_8802_29612# 0.143959f
C1229 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR 0.106927f
C1230 a_10170_35420# VPWR 0.39968f
C1231 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR 2.45124f
C1232 a_3762_27500# VPWR 0.382189f
C1233 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.166272f
C1234 a_20270_40296# VPWR 0.455248f
C1235 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145339f
C1236 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.149144f
C1237 a_6302_43816# SUNSAR_CAPT8B_CV_0.XC08.QN 0.129239f
C1238 a_10170_36300# VPWR 0.398846f
C1239 a_8802_32956# VPWR 0.436368f
C1240 a_18882_28556# VPWR 0.406628f
C1241 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CP0 0.331282f
C1242 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.638386f
C1243 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C1244 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.118161f
C1245 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.204048f
C1246 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.316693f
C1247 a_3782_41352# VPWR 0.394053f
C1248 SUNSAR_SAR8B_CV_0.EN ui_in[0] 0.969482f
C1249 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR 4.25322f
C1250 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18344f
C1251 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_2982# 0.158066f
C1252 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.301485f
C1253 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARN 0.591428f
C1254 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CN1 0.466806f
C1255 a_8802_35420# VPWR 0.39968f
C1256 SUNSAR_SAR8B_CV_0.XA4.XA10.Y a_12690_36300# 0.13253f
C1257 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR 2.44986f
C1258 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.166192f
C1259 a_18902_40296# VPWR 0.457343f
C1260 SUNSAR_CAPT8B_CV_0.XI14.QN uo_out[0] 0.25785f
C1261 a_8802_36300# VPWR 0.399161f
C1262 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 6.86675f
C1263 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.40569f
C1264 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_13842_35420# 0.133834f
C1265 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C1266 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C1267 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.2199f
C1268 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.129613f
C1269 VPWR ua[0] 0.493296f
C1270 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.126806f
C1271 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.293873f
C1272 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.318734f
C1273 a_10170_29612# VPWR 0.397362f
C1274 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.EN 0.315968f
C1275 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 6.86675f
C1276 a_9990_4918# VPWR 0.468783f
C1277 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARP 0.524159f
C1278 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y uo_out[4] 0.246349f
C1279 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VPWR 1.77562f
C1280 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR 2.45309f
C1281 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.241356f
C1282 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.166272f
C1283 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C1284 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35420# 0.160931f
C1285 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.118226f
C1286 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.398331f
C1287 VPWR ua[1] 0.225132f
C1288 uo_out[3] uo_out[2] 0.110956f
C1289 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_23922_29964# 0.151031f
C1290 SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR 0.635621f
C1291 a_10190_42760# VPWR 0.391454f
C1292 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.205884f
C1293 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C1294 a_8802_29612# VPWR 0.397362f
C1295 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.106828f
C1296 SUNSAR_SAR8B_CV_0.EN a_5130_29612# 0.143959f
C1297 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CN1 0.466806f
C1298 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y uo_out[4] 0.305131f
C1299 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR 2.95308f
C1300 SUNSAR_SAR8B_CV_0.XA3.XA10.Y a_11322_36300# 0.13402f
C1301 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR 2.45309f
C1302 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.393049f
C1303 a_7650_36828# SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.10248f
C1304 a_20250_27852# VPWR 0.358413f
C1305 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.166192f
C1306 a_5150_43816# VPWR 0.391817f
C1307 SUNSAR_CAPT8B_CV_0.XH13.QN uo_out[1] 0.254135f
C1308 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.375196f
C1309 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.EN 0.208884f
C1310 a_18902_41880# VPWR 0.395781f
C1311 a_5130_32956# VPWR 0.436368f
C1312 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.233892f
C1313 a_15210_28556# VPWR 0.406628f
C1314 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C1315 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.13041f
C1316 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.25689f
C1317 a_13862_40648# VPWR 0.491225f
C1318 VPWR ui_in[0] 1.19322f
C1319 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_22770_29964# 0.134249f
C1320 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.363295f
C1321 a_8822_42760# VPWR 0.391454f
C1322 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR 0.112858f
C1323 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1324 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D 0.107674f
C1325 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y a_10190_41880# 0.100592f
C1326 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARP 0.187721f
C1327 SUNSAR_SAR8B_CV_0.EN a_3762_29612# 0.143959f
C1328 a_5130_35420# VPWR 0.39968f
C1329 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR 2.45309f
C1330 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.105035f
C1331 a_18882_27852# VPWR 0.358599f
C1332 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.206912f
C1333 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C1334 a_15230_40296# VPWR 0.455577f
C1335 a_3782_43816# VPWR 0.391817f
C1336 a_5130_36300# VPWR 0.398846f
C1337 a_3762_32956# VPWR 0.436368f
C1338 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C1339 a_13842_28556# VPWR 0.406628f
C1340 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.327152f
C1341 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.118161f
C1342 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.79343f
C1343 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C1344 VPWR clk 0.645958f
C1345 uo_out[4] uo_out[3] 0.862834f
C1346 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.204048f
C1347 SUNSAR_SAR8B_CV_0.D<0> VPWR 5.48841f
C1348 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR 0.112858f
C1349 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87301f
C1350 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.379175p
C1351 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_2982# 0.158066f
C1352 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.174995f
C1353 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.301485f
C1354 a_16542_5270# VPWR 0.489055f
C1355 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.535136f
C1356 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR 0.106927f
C1357 a_3762_35420# VPWR 0.39968f
C1358 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR 2.45309f
C1359 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.649845f
C1360 a_13862_40296# VPWR 0.457343f
C1361 SUNSAR_CAPT8B_CV_0.XG12.QN uo_out[2] 0.254418f
C1362 a_3762_36300# VPWR 0.399161f
C1363 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1615f
C1364 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.129613f
C1365 SUNSAR_CAPT8B_CV_0.XA5.XA2.A a_22790_42408# 0.10248f
C1366 VPWR uo_out[0] 1.19196f
C1367 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.318734f
C1368 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR 0.106927f
C1369 a_5130_29612# VPWR 0.397362f
C1370 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.26479f
C1371 SUNSAR_CAPT8B_CV_0.XG12.XA4.A a_15230_42760# 0.111734f
C1372 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 27.1615f
C1373 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR 2.95307f
C1374 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR 2.45309f
C1375 a_6282_36828# SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.104051f
C1376 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.744161f
C1377 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.303428f
C1378 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR 11.7183f
C1379 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.383512f
C1380 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR 4.93712f
C1381 a_15230_41880# VPWR 0.395781f
C1382 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.118226f
C1383 VPWR uo_out[1] 1.02322f
C1384 a_10190_40648# VPWR 0.492624f
C1385 uo_out[5] uo_out[4] 1.16362f
C1386 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.316693f
C1387 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.M3.G 0.36754f
C1388 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR 0.106927f
C1389 a_5150_42760# VPWR 0.391454f
C1390 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR 3.09787f
C1391 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C1392 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.205884f
C1393 a_3762_29612# VPWR 0.397362f
C1394 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1395 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.669708f
C1396 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3334# 0.163985f
C1397 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_3334# 0.114704f
C1398 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.787331f
C1399 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.589705f
C1400 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.107823f
C1401 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.559553f
C1402 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y uo_out[5] 0.30523f
C1403 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VPWR 1.77562f
C1404 SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D VPWR 0.106794f
C1405 a_18902_41352# VPWR 0.394053f
C1406 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR 2.45309f
C1407 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.183415f
C1408 a_15210_27852# VPWR 0.358413f
C1409 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.244517f
C1410 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_3728# 0.172147f
C1411 a_23942_43992# VPWR 0.388156f
C1412 SUNSAR_CAPT8B_CV_0.XF11.QN uo_out[3] 0.267395f
C1413 a_23922_36652# VPWR 0.449853f
C1414 a_23922_33132# VPWR 0.415713f
C1415 a_13862_41880# VPWR 0.395781f
C1416 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.63636f
C1417 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.527529f
C1418 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35420# 0.160931f
C1419 a_10170_28556# VPWR 0.406628f
C1420 SUNSAR_CAPT8B_CV_0.XA4.MN0.S SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.138433f
C1421 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.13041f
C1422 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.394834f
C1423 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y a_21422_42408# 0.113479f
C1424 a_8822_40648# VPWR 0.491225f
C1425 uo_out[6] uo_out[4] 0.84361f
C1426 VPWR uo_out[2] 1.02322f
C1427 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.126806f
C1428 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_28556# 0.140127f
C1429 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.55251f
C1430 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.CMP_OP 7.93512f
C1431 SUNSAR_SAR8B_CV_0.D<1> VPWR 5.18522f
C1432 a_3782_42760# VPWR 0.391454f
C1433 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.433299f
C1434 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_3334# 0.118471f
C1435 a_9990_5270# VPWR 0.490626f
C1436 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C1437 SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR 0.658328f
C1438 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y uo_out[5] 0.245678f
C1439 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR 0.106927f
C1440 a_20270_41880# SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.100592f
C1441 a_13842_27852# VPWR 0.358599f
C1442 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C1443 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C1444 a_10190_40296# VPWR 0.455675f
C1445 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] 0.172623f
C1446 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_10170_35420# 0.133834f
C1447 a_8802_28556# VPWR 0.406628f
C1448 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.327909f
C1449 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.118161f
C1450 uo_out[6] uo_out[5] 0.327382f
C1451 uo_out[7] uo_out[4] 0.121957f
C1452 VPWR uo_out[3] 1.25759f
C1453 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1615f
C1454 a_20250_34716# VPWR 0.396749f
C1455 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C1456 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR 0.337652f
C1457 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.301485f
C1458 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR 0.808658f
C1459 a_10190_44168# VPWR 0.340085f
C1460 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.40569f
C1461 a_20250_31196# VPWR 0.437f
C1462 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.393055f
C1463 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA4.Y 0.504864f
C1464 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.240612f
C1465 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.18614f
C1466 a_8822_40296# VPWR 0.457343f
C1467 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.205975f
C1468 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[4] 0.249063f
C1469 SUNSAR_CAPT8B_CV_0.XI14.QN VPWR 0.901631f
C1470 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR 0.718455f
C1471 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6519f
C1472 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR 2.66621f
C1473 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y clk 0.210661f
C1474 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.449584f
C1475 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 5.19722f
C1476 uo_out[7] uo_out[5] 1.57818f
C1477 VPWR uo_out[4] 1.03096f
C1478 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.363295f
C1479 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB1.M3.G 0.175967f
C1480 SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR 9.342111f
C1481 a_18882_34716# VPWR 0.399819f
C1482 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.CKN 0.102131f
C1483 a_23922_29964# VPWR 0.429137f
C1484 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1485 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_4038# 0.135393f
C1486 SUNSAR_CAPT8B_CV_0.XF11.XA4.A a_13862_42760# 0.113305f
C1487 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6519f
C1488 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VPWR 1.77562f
C1489 SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR 1.20972f
C1490 a_15230_41352# VPWR 0.394053f
C1491 a_18882_31196# VPWR 0.44007f
C1492 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 0.241356f
C1493 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.178114f
C1494 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C1495 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.145048f
C1496 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.328435f
C1497 SUNSAR_CAPT8B_CV_0.XH13.QN VPWR 0.901622f
C1498 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.293159f
C1499 SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D VPWR 0.101562f
C1500 a_10190_41880# VPWR 0.395781f
C1501 SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR 2.64055f
C1502 a_5150_40648# VPWR 0.492592f
C1503 uo_out[7] uo_out[6] 2.38922f
C1504 VPWR uo_out[5] 1.0281f
C1505 SUNSAR_SAR8B_CV_0.D<2> VPWR 5.20829f
C1506 SUNSAR_SAR8B_CV_0.EN VPWR 41.784603f
C1507 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.98135f
C1508 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3334# 0.163985f
C1509 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3686# 0.16579f
C1510 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR 2.95303f
C1511 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR 0.924613f
C1512 a_13862_41352# VPWR 0.394053f
C1513 a_2610_36828# SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.10248f
C1514 a_10170_27852# VPWR 0.358413f
C1515 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C1516 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.693521f
C1517 SUNSAR_CAPT8B_CV_0.XG12.QN VPWR 0.901622f
C1518 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[5] 0.248535f
C1519 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.CEO 0.432008f
C1520 SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D VPWR 0.119314f
C1521 a_8822_41880# VPWR 0.395781f
C1522 SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR 2.64054f
C1523 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_8802_35420# 0.133834f
C1524 a_5130_28556# VPWR 0.406628f
C1525 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.449584f
C1526 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y a_17750_42408# 0.111909f
C1527 a_3782_40648# VPWR 0.491225f
C1528 VPWR uo_out[6] 1.34623f
C1529 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.55251f
C1530 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.SARP 5.22744f
C1531 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C1532 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.318734f
C1533 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR 0.106927f
C1534 a_23942_43112# VPWR 0.393308f
C1535 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_4390# 0.15559f
C1536 a_16542_5622# VPWR 0.472384f
C1537 SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR 1.22023f
C1538 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y uo_out[6] 0.251051f
C1539 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.744161f
C1540 a_8802_27852# VPWR 0.358599f
C1541 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C1542 a_5150_40296# VPWR 0.455605f
C1543 SUNSAR_CAPT8B_CV_0.XF11.QN VPWR 0.901622f
C1544 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.158152f
C1545 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR 0.725614f
C1546 SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR 2.64055f
C1547 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35420# 0.160931f
C1548 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA8.A 0.527529f
C1549 a_3762_28556# VPWR 0.406628f
C1550 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.327152f
C1551 ua[2] VGND 0.117454f
C1552 ua[3] VGND 0.117454f
C1553 ua[4] VGND 0.118698f
C1554 ua[5] VGND 0.120088f
C1555 ua[6] VGND 0.120088f
C1556 ua[7] VGND 0.111009f
C1557 ua[0] VGND 7.66672f
C1558 ua[1] VGND 6.98607f
C1559 ui_in[0] VGND 5.69254f
C1560 clk VGND 6.42293f
C1561 uo_out[0] VGND 2.81872f
C1562 uo_out[1] VGND 1.77173f
C1563 uo_out[2] VGND 1.57211f
C1564 uo_out[3] VGND 1.79184f
C1565 uo_out[4] VGND 1.64454f
C1566 uo_out[5] VGND 2.45226f
C1567 uo_out[6] VGND 2.74323f
C1568 uo_out[7] VGND 3.47431f
C1569 VPWR VGND 0.65886p
C1570 TIE_L1 VGND 1.5148f
C1571 TIE_L2 VGND 1.73849f
C1572 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93609f
C1573 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93609f
C1574 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.5533f
C1575 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.5533f
C1576 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.334839f
C1577 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.334839f
C1578 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.469f
C1579 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.469f
C1580 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43533f
C1581 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43533f
C1582 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67745f
C1583 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67745f
C1584 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.6684f
C1585 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.6684f
C1586 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.574499f
C1587 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.574499f
C1588 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33412f
C1589 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33412f
C1590 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.469f
C1591 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.469f
C1592 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43533f
C1593 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43533f
C1594 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67745f
C1595 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67745f
C1596 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.6684f
C1597 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.6684f
C1598 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.575099f
C1599 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.575099f
C1600 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33412f
C1601 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33412f
C1602 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.469f
C1603 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.469f
C1604 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43533f
C1605 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43533f
C1606 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67745f
C1607 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67745f
C1608 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.6684f
C1609 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.6684f
C1610 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.571799f
C1611 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.571799f
C1612 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33412f
C1613 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33412f
C1614 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.471901f
C1615 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.471901f
C1616 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.439809f
C1617 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44253f
C1618 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.3859f
C1619 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.38266f
C1620 a_15390_2630# VGND 0.542161f $ **FLOATING
C1621 a_13950_2630# VGND 0.427094f $ **FLOATING
C1622 a_12582_2630# VGND 0.426679f $ **FLOATING
C1623 a_11142_2630# VGND 0.543317f $ **FLOATING
C1624 a_15390_2982# VGND 0.491607f $ **FLOATING
C1625 a_13950_2982# VGND 0.352472f $ **FLOATING
C1626 a_12582_2982# VGND 0.352472f $ **FLOATING
C1627 a_11142_2982# VGND 0.490037f $ **FLOATING
C1628 a_15390_3334# VGND 0.374919f $ **FLOATING
C1629 a_13950_3334# VGND 0.352438f $ **FLOATING
C1630 a_12582_3334# VGND 0.352438f $ **FLOATING
C1631 a_11142_3334# VGND 0.374919f $ **FLOATING
C1632 a_13950_3686# VGND 0.352418f $ **FLOATING
C1633 a_12582_3686# VGND 0.352418f $ **FLOATING
C1634 SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND 41.5268f
C1635 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.70146f
C1636 SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND 41.5268f
C1637 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.70146f
C1638 a_15390_4038# VGND 0.397033f $ **FLOATING
C1639 a_13950_4038# VGND 0.354407f $ **FLOATING
C1640 a_12582_4038# VGND 0.354407f $ **FLOATING
C1641 a_11142_4038# VGND 0.397033f $ **FLOATING
C1642 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VGND 37.7832f
C1643 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.38998f
C1644 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D VGND 0.103625f
C1645 a_13950_4390# VGND 0.352432f $ **FLOATING
C1646 a_12582_4390# VGND 0.352432f $ **FLOATING
C1647 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D VGND 0.103625f
C1648 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.38998f
C1649 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VGND 37.7832f
C1650 SUNSAR_SAR8B_CV_0.XB2.M3.G VGND 3.1165f
C1651 a_15390_4566# VGND 0.389036f $ **FLOATING
C1652 SUNSAR_SAR8B_CV_0.XB1.M3.G VGND 3.07938f
C1653 a_11142_4566# VGND 0.389036f $ **FLOATING
C1654 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VGND 0.970036f
C1655 a_13950_4742# VGND 0.352456f $ **FLOATING
C1656 a_12582_4742# VGND 0.352456f $ **FLOATING
C1657 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND 0.7964f
C1658 a_15390_4918# VGND 0.470144f $ **FLOATING
C1659 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND 0.7964f
C1660 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VGND 0.970036f
C1661 a_11142_4918# VGND 0.471715f $ **FLOATING
C1662 a_13950_5094# VGND 0.353103f $ **FLOATING
C1663 a_12582_5094# VGND 0.353103f $ **FLOATING
C1664 a_15390_5270# VGND 0.492927f $ **FLOATING
C1665 a_11142_5270# VGND 0.491356f $ **FLOATING
C1666 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND 0.596866f
C1667 a_13950_5446# VGND 0.433341f $ **FLOATING
C1668 a_12582_5446# VGND 0.433756f $ **FLOATING
C1669 a_15390_5622# VGND 0.47219f $ **FLOATING
C1670 a_15390_5974# VGND 0.541341f $ **FLOATING
C1671 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND 0.596866f
C1672 a_11142_5622# VGND 0.47376f $ **FLOATING
C1673 a_11142_5974# VGND 0.540186f $ **FLOATING
C1674 a_22770_26796# VGND 0.529341f $ **FLOATING
C1675 a_21402_26796# VGND 0.531659f $ **FLOATING
C1676 a_17730_26796# VGND 0.530834f $ **FLOATING
C1677 a_16362_26796# VGND 0.531989f $ **FLOATING
C1678 a_12690_26796# VGND 0.530834f $ **FLOATING
C1679 a_11322_26796# VGND 0.531989f $ **FLOATING
C1680 a_7650_26796# VGND 0.530213f $ **FLOATING
C1681 a_6282_26796# VGND 0.530979f $ **FLOATING
C1682 a_2610_26796# VGND 0.531178f $ **FLOATING
C1683 a_22770_27148# VGND 0.499848f $ **FLOATING
C1684 a_21402_27148# VGND 0.467094f $ **FLOATING
C1685 a_17730_27148# VGND 0.471508f $ **FLOATING
C1686 a_16362_27148# VGND 0.467722f $ **FLOATING
C1687 a_12690_27148# VGND 0.471508f $ **FLOATING
C1688 a_11322_27148# VGND 0.467722f $ **FLOATING
C1689 a_7650_27148# VGND 0.470266f $ **FLOATING
C1690 a_6282_27148# VGND 0.465734f $ **FLOATING
C1691 a_2610_27148# VGND 0.47123f $ **FLOATING
C1692 a_21402_27500# VGND 0.385968f $ **FLOATING
C1693 a_17730_27500# VGND 0.387712f $ **FLOATING
C1694 a_16362_27500# VGND 0.386249f $ **FLOATING
C1695 a_12690_27500# VGND 0.387712f $ **FLOATING
C1696 a_11322_27500# VGND 0.386249f $ **FLOATING
C1697 a_7650_27500# VGND 0.38671f $ **FLOATING
C1698 a_6282_27500# VGND 0.384229f $ **FLOATING
C1699 a_2610_27500# VGND 0.387675f $ **FLOATING
C1700 a_21402_27852# VGND 0.370125f $ **FLOATING
C1701 a_17730_27852# VGND 0.370785f $ **FLOATING
C1702 a_16362_27852# VGND 0.368771f $ **FLOATING
C1703 a_12690_27852# VGND 0.370785f $ **FLOATING
C1704 a_11322_27852# VGND 0.368771f $ **FLOATING
C1705 a_7650_27852# VGND 0.369543f $ **FLOATING
C1706 a_6282_27852# VGND 0.366751f $ **FLOATING
C1707 a_2610_27852# VGND 0.370508f $ **FLOATING
C1708 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D VGND 0.506947f
C1709 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D VGND 0.502211f
C1710 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D VGND 0.477244f
C1711 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D VGND 0.502211f
C1712 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D VGND 0.477244f
C1713 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D VGND 0.502211f
C1714 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D VGND 0.477244f
C1715 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D VGND 0.502211f
C1716 a_21402_28204# VGND 0.405715f $ **FLOATING
C1717 a_17730_28204# VGND 0.406284f $ **FLOATING
C1718 a_16362_28204# VGND 0.406284f $ **FLOATING
C1719 a_12690_28204# VGND 0.406284f $ **FLOATING
C1720 a_11322_28204# VGND 0.406284f $ **FLOATING
C1721 a_7650_28204# VGND 0.405133f $ **FLOATING
C1722 a_6282_28204# VGND 0.404355f $ **FLOATING
C1723 a_2610_28204# VGND 0.406098f $ **FLOATING
C1724 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND 0.608956f
C1725 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND 0.741242f
C1726 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND 0.749251f
C1727 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND 0.735502f
C1728 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND 0.749251f
C1729 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND 0.735502f
C1730 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND 0.746591f
C1731 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND 0.73057f
C1732 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND 0.74895f
C1733 a_22770_28556# VGND 0.401649f $ **FLOATING
C1734 a_21402_28556# VGND 0.387558f $ **FLOATING
C1735 a_17730_28556# VGND 0.388127f $ **FLOATING
C1736 a_16362_28556# VGND 0.388127f $ **FLOATING
C1737 a_12690_28556# VGND 0.388127f $ **FLOATING
C1738 a_11322_28556# VGND 0.388127f $ **FLOATING
C1739 a_7650_28556# VGND 0.386976f $ **FLOATING
C1740 a_6282_28556# VGND 0.386198f $ **FLOATING
C1741 a_2610_28556# VGND 0.38794f $ **FLOATING
C1742 a_21402_28908# VGND 0.394283f $ **FLOATING
C1743 a_17730_28908# VGND 0.394852f $ **FLOATING
C1744 a_16362_28908# VGND 0.394852f $ **FLOATING
C1745 a_12690_28908# VGND 0.394852f $ **FLOATING
C1746 a_11322_28908# VGND 0.394852f $ **FLOATING
C1747 a_7650_28908# VGND 0.393701f $ **FLOATING
C1748 a_6282_28908# VGND 0.392923f $ **FLOATING
C1749 a_2610_28908# VGND 0.394666f $ **FLOATING
C1750 SUNSAR_SAR8B_CV_0.SARP VGND 70.097496f
C1751 a_21402_29612# VGND 0.395457f $ **FLOATING
C1752 a_17730_29612# VGND 0.396116f $ **FLOATING
C1753 a_16362_29612# VGND 0.395588f $ **FLOATING
C1754 a_12690_29612# VGND 0.396116f $ **FLOATING
C1755 a_11322_29612# VGND 0.395588f $ **FLOATING
C1756 a_7650_29612# VGND 0.394965f $ **FLOATING
C1757 a_6282_29612# VGND 0.393746f $ **FLOATING
C1758 a_2610_29612# VGND 0.395923f $ **FLOATING
C1759 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318647f
C1760 a_22770_29964# VGND 0.400512f $ **FLOATING
C1761 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D VGND 0.103281f
C1762 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VGND 1.27143f
C1763 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D VGND 0.100021f
C1764 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VGND 1.26503f
C1765 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D VGND 0.100021f
C1766 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VGND 1.26391f
C1767 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D VGND 0.100021f
C1768 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VGND 1.26503f
C1769 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D VGND 0.100021f
C1770 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VGND 1.26391f
C1771 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D VGND 0.100021f
C1772 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VGND 1.25938f
C1773 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D VGND 0.100021f
C1774 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VGND 1.25329f
C1775 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D VGND 0.100021f
C1776 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VGND 1.26407f
C1777 a_21402_30316# VGND 0.401758f $ **FLOATING
C1778 a_17730_30316# VGND 0.401074f $ **FLOATING
C1779 a_16362_30316# VGND 0.401074f $ **FLOATING
C1780 a_12690_30316# VGND 0.401074f $ **FLOATING
C1781 a_11322_30316# VGND 0.401074f $ **FLOATING
C1782 a_7650_30316# VGND 0.399923f $ **FLOATING
C1783 a_6282_30316# VGND 0.399145f $ **FLOATING
C1784 a_2610_30316# VGND 0.400881f $ **FLOATING
C1785 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND 15.315499f
C1786 a_22770_30844# VGND 0.421853f $ **FLOATING
C1787 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND 2.24318f
C1788 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND 2.22194f
C1789 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND 2.22198f
C1790 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND 2.22194f
C1791 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND 2.22198f
C1792 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND 2.20909f
C1793 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND 2.19751f
C1794 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND 2.21827f
C1795 a_21402_31196# VGND 0.4255f $ **FLOATING
C1796 a_17730_31196# VGND 0.426069f $ **FLOATING
C1797 a_16362_31196# VGND 0.426069f $ **FLOATING
C1798 a_12690_31196# VGND 0.426069f $ **FLOATING
C1799 a_11322_31196# VGND 0.426069f $ **FLOATING
C1800 a_7650_31196# VGND 0.424917f $ **FLOATING
C1801 a_6282_31196# VGND 0.42414f $ **FLOATING
C1802 a_2610_31196# VGND 0.425876f $ **FLOATING
C1803 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND 19.4783f
C1804 a_22770_31724# VGND 0.423601f $ **FLOATING
C1805 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.99939f
C1806 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.97987f
C1807 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.97901f
C1808 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.97987f
C1809 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.97901f
C1810 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.85828f
C1811 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.37577f
C1812 a_21402_32076# VGND 0.426091f $ **FLOATING
C1813 a_17730_32076# VGND 0.42666f $ **FLOATING
C1814 a_16362_32076# VGND 0.42666f $ **FLOATING
C1815 a_12690_32076# VGND 0.42666f $ **FLOATING
C1816 a_11322_32076# VGND 0.42666f $ **FLOATING
C1817 a_7650_32076# VGND 0.42666f $ **FLOATING
C1818 a_6282_32076# VGND 0.42666f $ **FLOATING
C1819 a_2610_32076# VGND 0.426468f $ **FLOATING
C1820 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND 1.55564f
C1821 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C1822 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND 3.19736f
C1823 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND 3.22974f
C1824 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND 3.22835f
C1825 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND 3.22974f
C1826 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND 3.22835f
C1827 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND 3.22678f
C1828 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND 3.22545f
C1829 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND 3.31413f
C1830 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND 2.68549f
C1831 a_21402_32956# VGND 0.426069f $ **FLOATING
C1832 a_17730_32956# VGND 0.426069f $ **FLOATING
C1833 a_16362_32956# VGND 0.426069f $ **FLOATING
C1834 a_12690_32956# VGND 0.426069f $ **FLOATING
C1835 a_11322_32956# VGND 0.426069f $ **FLOATING
C1836 a_7650_32956# VGND 0.426069f $ **FLOATING
C1837 a_6282_32956# VGND 0.426069f $ **FLOATING
C1838 a_2610_32956# VGND 0.425876f $ **FLOATING
C1839 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND 2.85099f
C1840 a_22770_33132# VGND 0.403395f $ **FLOATING
C1841 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 3.01164f
C1842 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.01628f
C1843 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.01641f
C1844 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.01628f
C1845 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.01641f
C1846 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.54669f
C1847 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.78758f
C1848 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 12.1041f
C1849 a_21402_33836# VGND 0.426756f $ **FLOATING
C1850 a_17730_33836# VGND 0.426756f $ **FLOATING
C1851 a_16362_33836# VGND 0.426756f $ **FLOATING
C1852 a_12690_33836# VGND 0.426756f $ **FLOATING
C1853 a_11322_33836# VGND 0.426756f $ **FLOATING
C1854 a_7650_33836# VGND 0.426756f $ **FLOATING
C1855 a_6282_33836# VGND 0.426756f $ **FLOATING
C1856 a_2610_33836# VGND 0.426472f $ **FLOATING
C1857 SUNSAR_SAR8B_CV_0.SARN VGND 71.1589f
C1858 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND 0.149691f
C1859 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND 0.515385f
C1860 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C1861 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND 0.149691f
C1862 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.72791f
C1863 a_22770_34540# VGND 0.39377f $ **FLOATING
C1864 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND 0.102f
C1865 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND 0.149691f
C1866 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 4.1719f
C1867 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND 0.149691f
C1868 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.27991f
C1869 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND 0.102f
C1870 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND 0.102f
C1871 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND 0.149691f
C1872 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.31299f
C1873 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND 0.149691f
C1874 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.68294f
C1875 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND 0.102f
C1876 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND 0.102f
C1877 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND 0.149691f
C1878 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 4.25175f
C1879 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND 0.149691f
C1880 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 10.150401f
C1881 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND 0.102f
C1882 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND 0.102f
C1883 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND 0.102f
C1884 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 8.127279f
C1885 a_21402_34716# VGND 0.39476f $ **FLOATING
C1886 a_17730_34716# VGND 0.39476f $ **FLOATING
C1887 a_16362_34716# VGND 0.39476f $ **FLOATING
C1888 a_12690_34716# VGND 0.39476f $ **FLOATING
C1889 a_11322_34716# VGND 0.39476f $ **FLOATING
C1890 a_7650_34716# VGND 0.39476f $ **FLOATING
C1891 a_6282_34716# VGND 0.39476f $ **FLOATING
C1892 a_2610_34716# VGND 0.394567f $ **FLOATING
C1893 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND 4.75219f
C1894 a_22770_34892# VGND 0.394644f $ **FLOATING
C1895 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.67603f
C1896 SUNSAR_SAR8B_CV_0.XA6.ENO VGND 4.51439f
C1897 SUNSAR_SAR8B_CV_0.XA5.ENO VGND 4.46191f
C1898 SUNSAR_SAR8B_CV_0.XA4.ENO VGND 4.27708f
C1899 SUNSAR_SAR8B_CV_0.XA3.ENO VGND 4.50282f
C1900 SUNSAR_SAR8B_CV_0.XA2.ENO VGND 4.42572f
C1901 SUNSAR_SAR8B_CV_0.XA1.ENO VGND 4.44437f
C1902 SUNSAR_SAR8B_CV_0.XA0.ENO VGND 4.39222f
C1903 a_21402_35068# VGND 0.389563f $ **FLOATING
C1904 a_17730_35068# VGND 0.389563f $ **FLOATING
C1905 a_16362_35068# VGND 0.389563f $ **FLOATING
C1906 a_12690_35068# VGND 0.389563f $ **FLOATING
C1907 a_11322_35068# VGND 0.389563f $ **FLOATING
C1908 a_7650_35068# VGND 0.389563f $ **FLOATING
C1909 a_6282_35068# VGND 0.389563f $ **FLOATING
C1910 a_2610_35068# VGND 0.38937f $ **FLOATING
C1911 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND 4.54316f
C1912 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C1913 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C1914 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C1915 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C1916 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C1917 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C1918 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557214f
C1919 a_22770_35420# VGND 0.395535f $ **FLOATING
C1920 a_21402_35420# VGND 0.389041f $ **FLOATING
C1921 a_17730_35420# VGND 0.388925f $ **FLOATING
C1922 a_16362_35420# VGND 0.389297f $ **FLOATING
C1923 a_12690_35420# VGND 0.388925f $ **FLOATING
C1924 a_11322_35420# VGND 0.389297f $ **FLOATING
C1925 a_7650_35420# VGND 0.388925f $ **FLOATING
C1926 a_6282_35420# VGND 0.389297f $ **FLOATING
C1927 a_2610_35420# VGND 0.389015f $ **FLOATING
C1928 SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND 1.07685f
C1929 SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D VGND 0.112889f
C1930 SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND 1.50901f
C1931 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VGND 1.53168f
C1932 SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND 1.50964f
C1933 SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D VGND 0.112889f
C1934 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VGND 1.54335f
C1935 SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D VGND 0.112889f
C1936 SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND 1.51005f
C1937 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VGND 1.53305f
C1938 SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND 1.50964f
C1939 SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D VGND 0.112889f
C1940 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VGND 1.54335f
C1941 SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D VGND 0.112889f
C1942 SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND 1.51005f
C1943 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VGND 1.53305f
C1944 SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND 1.50964f
C1945 SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D VGND 0.112889f
C1946 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VGND 1.54335f
C1947 SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D VGND 0.112889f
C1948 SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND 1.51005f
C1949 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VGND 1.53305f
C1950 SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND 1.51935f
C1951 SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D VGND 0.112889f
C1952 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VGND 1.61753f
C1953 a_22770_35948# VGND 0.414038f $ **FLOATING
C1954 a_21402_35948# VGND 0.390722f $ **FLOATING
C1955 a_17730_35948# VGND 0.391291f $ **FLOATING
C1956 a_16362_35948# VGND 0.391291f $ **FLOATING
C1957 a_12690_35948# VGND 0.391291f $ **FLOATING
C1958 a_11322_35948# VGND 0.391291f $ **FLOATING
C1959 a_7650_35948# VGND 0.391291f $ **FLOATING
C1960 a_6282_35948# VGND 0.391291f $ **FLOATING
C1961 a_2610_35948# VGND 0.391099f $ **FLOATING
C1962 SUNSAR_SAR8B_CV_0.XA20.XA10.B VGND 0.789814f
C1963 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C1964 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C1965 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C1966 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C1967 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C1968 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C1969 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C1970 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.895311f
C1971 a_22770_36300# VGND 0.472701f $ **FLOATING
C1972 a_21402_36300# VGND 0.393831f $ **FLOATING
C1973 a_17730_36300# VGND 0.394738f $ **FLOATING
C1974 a_16362_36300# VGND 0.3944f $ **FLOATING
C1975 a_12690_36300# VGND 0.394718f $ **FLOATING
C1976 a_11322_36300# VGND 0.3944f $ **FLOATING
C1977 a_7650_36300# VGND 0.394715f $ **FLOATING
C1978 a_6282_36300# VGND 0.3944f $ **FLOATING
C1979 a_2610_36300# VGND 0.394523f $ **FLOATING
C1980 a_22770_36652# VGND 0.542245f $ **FLOATING
C1981 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND 0.881626f
C1982 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND 0.884627f
C1983 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND 0.877071f
C1984 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND 0.884604f
C1985 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND 0.877059f
C1986 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND 0.884603f
C1987 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND 0.877071f
C1988 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND 0.892649f
C1989 SUNSAR_SAR8B_CV_0.XB1.TIE_L VGND 32.9183f
C1990 a_21402_36828# VGND 0.414041f $ **FLOATING
C1991 a_17730_36828# VGND 0.413952f $ **FLOATING
C1992 a_16362_36828# VGND 0.413659f $ **FLOATING
C1993 a_12690_36828# VGND 0.413942f $ **FLOATING
C1994 a_11322_36828# VGND 0.413658f $ **FLOATING
C1995 a_7650_36828# VGND 0.413944f $ **FLOATING
C1996 a_6282_36828# VGND 0.413659f $ **FLOATING
C1997 a_2610_36828# VGND 0.413594f $ **FLOATING
C1998 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND 1.08552f
C1999 SUNSAR_SAR8B_CV_0.XA7.CEO VGND 2.06017f
C2000 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND 1.10839f
C2001 SUNSAR_SAR8B_CV_0.XA6.CEO VGND 1.45333f
C2002 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND 1.06778f
C2003 SUNSAR_SAR8B_CV_0.XA5.CEO VGND 1.71757f
C2004 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND 1.10834f
C2005 SUNSAR_SAR8B_CV_0.XA4.CEO VGND 1.52588f
C2006 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND 1.06777f
C2007 SUNSAR_SAR8B_CV_0.XA3.CEO VGND 1.71756f
C2008 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND 1.10835f
C2009 SUNSAR_SAR8B_CV_0.XA2.CEO VGND 1.52589f
C2010 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND 1.06778f
C2011 SUNSAR_SAR8B_CV_0.XA1.CEO VGND 1.71756f
C2012 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND 1.11927f
C2013 SUNSAR_SAR8B_CV_0.XA0.CEO VGND 1.53308f
C2014 a_21402_37180# VGND 0.47501f $ **FLOATING
C2015 a_17730_37180# VGND 0.474809f $ **FLOATING
C2016 a_16362_37180# VGND 0.476355f $ **FLOATING
C2017 a_12690_37180# VGND 0.47479f $ **FLOATING
C2018 a_11322_37180# VGND 0.476354f $ **FLOATING
C2019 a_7650_37180# VGND 0.474794f $ **FLOATING
C2020 a_6282_37180# VGND 0.476355f $ **FLOATING
C2021 a_2610_37180# VGND 0.474277f $ **FLOATING
C2022 a_21402_37532# VGND 0.546649f $ **FLOATING
C2023 a_17730_37532# VGND 0.548986f $ **FLOATING
C2024 a_16362_37532# VGND 0.547631f $ **FLOATING
C2025 a_12690_37532# VGND 0.548815f $ **FLOATING
C2026 a_11322_37532# VGND 0.547631f $ **FLOATING
C2027 a_7650_37532# VGND 0.548857f $ **FLOATING
C2028 a_6282_37532# VGND 0.547634f $ **FLOATING
C2029 a_2610_37532# VGND 0.546853f $ **FLOATING
C2030 a_22790_40296# VGND 0.546732f $ **FLOATING
C2031 a_21422_40296# VGND 0.54563f $ **FLOATING
C2032 a_17750_40296# VGND 0.546813f $ **FLOATING
C2033 a_16382_40296# VGND 0.547966f $ **FLOATING
C2034 a_12710_40296# VGND 0.546813f $ **FLOATING
C2035 a_11342_40296# VGND 0.547969f $ **FLOATING
C2036 a_7670_40296# VGND 0.54681f $ **FLOATING
C2037 a_6302_40296# VGND 0.547966f $ **FLOATING
C2038 a_2630_40296# VGND 0.54539f $ **FLOATING
C2039 a_22790_40648# VGND 0.492438f $ **FLOATING
C2040 a_21422_40648# VGND 0.49034f $ **FLOATING
C2041 a_17750_40648# VGND 0.492453f $ **FLOATING
C2042 a_16382_40648# VGND 0.490883f $ **FLOATING
C2043 a_12710_40648# VGND 0.492453f $ **FLOATING
C2044 a_11342_40648# VGND 0.490883f $ **FLOATING
C2045 a_7670_40648# VGND 0.492453f $ **FLOATING
C2046 a_6302_40648# VGND 0.490883f $ **FLOATING
C2047 a_2630_40648# VGND 0.492826f $ **FLOATING
C2048 SUNSAR_SAR8B_CV_0.DONE VGND 20.737402f
C2049 a_22790_41000# VGND 0.388777f $ **FLOATING
C2050 a_21422_41000# VGND 0.388174f $ **FLOATING
C2051 a_17750_41000# VGND 0.388174f $ **FLOATING
C2052 a_16382_41000# VGND 0.388174f $ **FLOATING
C2053 a_12710_41000# VGND 0.388174f $ **FLOATING
C2054 a_11342_41000# VGND 0.388174f $ **FLOATING
C2055 a_7670_41000# VGND 0.388174f $ **FLOATING
C2056 a_6302_41000# VGND 0.388174f $ **FLOATING
C2057 a_2630_41000# VGND 0.388638f $ **FLOATING
C2058 a_22790_41352# VGND 0.374594f $ **FLOATING
C2059 a_21422_41352# VGND 0.393558f $ **FLOATING
C2060 a_17750_41352# VGND 0.393558f $ **FLOATING
C2061 a_16382_41352# VGND 0.393558f $ **FLOATING
C2062 a_12710_41352# VGND 0.393558f $ **FLOATING
C2063 a_11342_41352# VGND 0.393558f $ **FLOATING
C2064 a_7670_41352# VGND 0.393558f $ **FLOATING
C2065 a_6302_41352# VGND 0.393558f $ **FLOATING
C2066 a_2630_41352# VGND 0.394022f $ **FLOATING
C2067 SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND 0.803097f
C2068 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND 0.107737f
C2069 SUNSAR_SAR8B_CV_0.D<0> VGND 5.87227f
C2070 SUNSAR_SAR8B_CV_0.D<1> VGND 13.789701f
C2071 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND 0.107643f
C2072 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND 0.107643f
C2073 SUNSAR_SAR8B_CV_0.D<2> VGND 12.5832f
C2074 SUNSAR_SAR8B_CV_0.D<3> VGND 11.4395f
C2075 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND 0.107643f
C2076 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND 0.107643f
C2077 SUNSAR_SAR8B_CV_0.D<4> VGND 11.8306f
C2078 SUNSAR_SAR8B_CV_0.D<5> VGND 12.7012f
C2079 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND 0.107643f
C2080 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND 0.107643f
C2081 SUNSAR_SAR8B_CV_0.D<6> VGND 12.0145f
C2082 SUNSAR_SAR8B_CV_0.D<7> VGND 17.833302f
C2083 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND 0.107643f
C2084 a_22790_41880# VGND 0.394408f $ **FLOATING
C2085 a_21422_41880# VGND 0.395138f $ **FLOATING
C2086 a_17750_41880# VGND 0.395707f $ **FLOATING
C2087 a_16382_41880# VGND 0.395707f $ **FLOATING
C2088 a_12710_41880# VGND 0.395707f $ **FLOATING
C2089 a_11342_41880# VGND 0.395707f $ **FLOATING
C2090 a_7670_41880# VGND 0.395707f $ **FLOATING
C2091 a_6302_41880# VGND 0.395707f $ **FLOATING
C2092 a_2630_41880# VGND 0.396052f $ **FLOATING
C2093 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND 1.96193f
C2094 a_22790_42408# VGND 0.410698f $ **FLOATING
C2095 a_21422_42408# VGND 0.389697f $ **FLOATING
C2096 a_17750_42408# VGND 0.390266f $ **FLOATING
C2097 a_16382_42408# VGND 0.390266f $ **FLOATING
C2098 a_12710_42408# VGND 0.390266f $ **FLOATING
C2099 a_11342_42408# VGND 0.390266f $ **FLOATING
C2100 a_7670_42408# VGND 0.390266f $ **FLOATING
C2101 a_6302_42408# VGND 0.390266f $ **FLOATING
C2102 a_2630_42408# VGND 0.390612f $ **FLOATING
C2103 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C2104 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND 1.28758f
C2105 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND 1.27933f
C2106 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND 1.27933f
C2107 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND 1.27933f
C2108 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND 1.27933f
C2109 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND 1.27933f
C2110 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND 1.27933f
C2111 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND 1.29578f
C2112 a_22790_42760# VGND 0.378208f $ **FLOATING
C2113 a_21422_42760# VGND 0.393027f $ **FLOATING
C2114 a_17750_42760# VGND 0.393596f $ **FLOATING
C2115 a_16382_42760# VGND 0.393596f $ **FLOATING
C2116 a_12710_42760# VGND 0.393596f $ **FLOATING
C2117 a_11342_42760# VGND 0.393596f $ **FLOATING
C2118 a_7670_42760# VGND 0.393596f $ **FLOATING
C2119 a_6302_42760# VGND 0.393596f $ **FLOATING
C2120 a_2630_42760# VGND 0.393942f $ **FLOATING
C2121 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 24.7108f
C2122 SUNSAR_SAR8B_CV_0.EN VGND 11.027699f
C2123 a_22790_43112# VGND 0.388427f $ **FLOATING
C2124 SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND 1.29446f
C2125 SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND 1.29655f
C2126 SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND 1.29655f
C2127 SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND 1.29655f
C2128 SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND 1.29655f
C2129 SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND 1.29655f
C2130 SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND 1.29655f
C2131 SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND 1.29893f
C2132 SUNSAR_CAPT8B_CV_0.XA4.Y VGND 2.38165f
C2133 a_21422_43288# VGND 0.394124f $ **FLOATING
C2134 a_17750_43288# VGND 0.394693f $ **FLOATING
C2135 a_16382_43288# VGND 0.394693f $ **FLOATING
C2136 a_12710_43288# VGND 0.394693f $ **FLOATING
C2137 a_11342_43288# VGND 0.394693f $ **FLOATING
C2138 a_7670_43288# VGND 0.394693f $ **FLOATING
C2139 a_6302_43288# VGND 0.394693f $ **FLOATING
C2140 a_2630_43288# VGND 0.395039f $ **FLOATING
C2141 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D VGND 0.103608f
C2142 SUNSAR_CAPT8B_CV_0.XA3.Y VGND 1.65429f
C2143 a_22790_43640# VGND 0.387806f $ **FLOATING
C2144 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND 0.112889f
C2145 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND 2.60322f
C2146 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VGND 1.6954f
C2147 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND 0.112889f
C2148 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VGND 1.69797f
C2149 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND 2.58593f
C2150 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND 0.112889f
C2151 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND 2.6374f
C2152 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VGND 1.69797f
C2153 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND 0.112889f
C2154 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VGND 1.69797f
C2155 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND 2.63726f
C2156 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND 0.112889f
C2157 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND 2.59274f
C2158 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VGND 1.69797f
C2159 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND 0.112889f
C2160 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VGND 1.69797f
C2161 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND 2.5926f
C2162 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND 0.112889f
C2163 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND 2.6374f
C2164 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VGND 1.69797f
C2165 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND 0.112889f
C2166 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VGND 1.69726f
C2167 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND 2.70316f
C2168 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.891538f
C2169 a_21422_43816# VGND 0.390629f $ **FLOATING
C2170 a_17750_43816# VGND 0.391198f $ **FLOATING
C2171 a_16382_43816# VGND 0.391198f $ **FLOATING
C2172 a_12710_43816# VGND 0.391198f $ **FLOATING
C2173 a_11342_43816# VGND 0.391198f $ **FLOATING
C2174 a_7670_43816# VGND 0.391198f $ **FLOATING
C2175 a_6302_43816# VGND 0.391198f $ **FLOATING
C2176 a_2630_43816# VGND 0.391544f $ **FLOATING
C2177 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 24.566801f
C2178 a_22790_43992# VGND 0.384235f $ **FLOATING
C2179 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.26356f
C2180 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.26291f
C2181 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.26291f
C2182 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.26291f
C2183 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26291f
C2184 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C2185 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C2186 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C2187 SUNSAR_CAPT8B_CV_0.XA2.MN0.G VGND 0.651712f
C2188 a_21422_44168# VGND 0.425534f $ **FLOATING
C2189 a_17750_44168# VGND 0.425449f $ **FLOATING
C2190 a_16382_44168# VGND 0.425864f $ **FLOATING
C2191 a_12710_44168# VGND 0.425449f $ **FLOATING
C2192 a_11342_44168# VGND 0.425864f $ **FLOATING
C2193 a_7670_44168# VGND 0.425449f $ **FLOATING
C2194 a_6302_44168# VGND 0.425864f $ **FLOATING
C2195 a_2630_44168# VGND 0.426034f $ **FLOATING
C2196 TIE_L VGND 6.84182f
C2197 a_22790_44344# VGND 0.423601f $ **FLOATING
.ends

