VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_TT06_SAR_wulffern
  CLASS BLOCK ;
  FOREIGN tt_um_TT06_SAR_wulffern ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.156000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 6.156000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.615600 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.388800 ;
    ANTENNADIFFAREA 1.231200 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.000 5.000 157.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 111.430 221.590 118.630 222.470 ;
        RECT 10.630 200.910 17.830 221.590 ;
      LAYER nwell ;
        RECT 17.830 200.910 30.430 221.590 ;
      LAYER pwell ;
        RECT 30.430 200.910 43.030 221.590 ;
      LAYER nwell ;
        RECT 43.030 200.910 55.630 221.590 ;
      LAYER pwell ;
        RECT 55.630 200.910 68.230 221.590 ;
      LAYER nwell ;
        RECT 68.230 200.910 80.830 221.590 ;
      LAYER pwell ;
        RECT 80.830 200.910 93.430 221.590 ;
      LAYER nwell ;
        RECT 93.430 200.910 106.030 221.590 ;
      LAYER pwell ;
        RECT 106.030 200.910 118.630 221.590 ;
      LAYER nwell ;
        RECT 118.630 200.910 125.830 222.470 ;
      LAYER pwell ;
        RECT 135.355 199.205 142.555 207.565 ;
      LAYER nwell ;
        RECT 142.555 199.205 149.755 207.565 ;
      LAYER pwell ;
        RECT 10.530 133.410 17.730 188.410 ;
      LAYER nwell ;
        RECT 17.730 133.410 30.330 188.410 ;
      LAYER pwell ;
        RECT 30.330 133.410 42.930 188.410 ;
      LAYER nwell ;
        RECT 42.930 133.410 55.530 188.410 ;
      LAYER pwell ;
        RECT 55.530 133.410 68.130 188.410 ;
      LAYER nwell ;
        RECT 68.130 133.410 80.730 188.410 ;
      LAYER pwell ;
        RECT 80.730 133.410 93.330 188.410 ;
      LAYER nwell ;
        RECT 93.330 133.410 105.930 188.410 ;
      LAYER pwell ;
        RECT 105.930 184.010 113.130 188.410 ;
        RECT 105.930 133.410 118.530 184.010 ;
      LAYER nwell ;
        RECT 118.530 133.410 125.730 184.010 ;
        RECT 47.430 12.580 54.630 30.620 ;
      LAYER pwell ;
        RECT 54.630 27.980 61.830 30.620 ;
        RECT 74.430 27.980 81.630 30.620 ;
        RECT 54.630 12.580 81.630 27.980 ;
      LAYER nwell ;
        RECT 81.630 12.580 88.830 30.620 ;
      LAYER li1 ;
        RECT 60.120 224.020 136.740 224.320 ;
        RECT 112.640 223.020 135.510 223.320 ;
        RECT 10.990 202.620 12.070 221.150 ;
        RECT 15.310 220.320 20.350 220.660 ;
        RECT 13.150 219.880 14.870 220.220 ;
        RECT 21.430 219.880 22.510 220.220 ;
        RECT 14.530 218.900 14.870 219.880 ;
        RECT 15.310 219.440 16.390 219.780 ;
        RECT 19.270 219.440 20.350 219.780 ;
        RECT 14.530 218.560 20.350 218.900 ;
        RECT 13.150 218.120 14.230 218.460 ;
        RECT 15.310 217.680 16.390 218.020 ;
        RECT 13.150 217.240 14.230 217.580 ;
        RECT 15.310 216.800 16.390 217.140 ;
        RECT 16.690 216.260 17.030 218.560 ;
        RECT 20.650 218.120 22.510 218.460 ;
        RECT 19.270 217.680 20.350 218.020 ;
        RECT 19.270 216.800 20.350 217.140 ;
        RECT 15.310 215.920 20.350 216.260 ;
        RECT 13.150 215.480 14.230 215.820 ;
        RECT 13.930 215.140 14.870 215.480 ;
        RECT 13.150 214.600 14.230 214.940 ;
        RECT 13.150 212.840 14.230 213.180 ;
        RECT 14.530 211.420 14.870 215.140 ;
        RECT 15.310 215.040 16.390 215.380 ;
        RECT 19.270 215.040 20.350 215.380 ;
        RECT 15.310 214.160 16.390 214.500 ;
        RECT 19.270 214.160 20.350 214.500 ;
        RECT 15.310 213.280 20.350 213.620 ;
        RECT 15.310 212.400 16.390 212.740 ;
        RECT 19.270 212.400 20.350 212.740 ;
        RECT 15.310 211.520 20.350 211.860 ;
        RECT 13.150 211.080 14.870 211.420 ;
        RECT 13.150 210.200 14.230 210.540 ;
        RECT 13.150 208.440 14.230 208.780 ;
        RECT 13.150 207.560 14.230 207.900 ;
        RECT 14.530 206.580 14.870 211.080 ;
        RECT 15.310 210.640 16.390 210.980 ;
        RECT 15.310 209.760 16.390 210.100 ;
        RECT 16.690 209.220 17.030 211.520 ;
        RECT 19.270 210.640 20.350 210.980 ;
        RECT 19.270 209.760 20.350 210.100 ;
        RECT 15.310 208.880 20.350 209.220 ;
        RECT 20.650 208.780 20.990 218.120 ;
        RECT 21.430 217.240 22.510 217.580 ;
        RECT 21.430 215.480 22.510 215.820 ;
        RECT 21.430 214.600 22.510 214.940 ;
        RECT 21.430 212.840 22.510 213.180 ;
        RECT 21.430 211.080 22.510 211.420 ;
        RECT 21.430 210.200 22.510 210.540 ;
        RECT 20.650 208.440 22.510 208.780 ;
        RECT 15.310 208.000 16.390 208.340 ;
        RECT 19.270 208.000 20.350 208.340 ;
        RECT 15.310 207.120 16.390 207.460 ;
        RECT 19.270 207.120 20.350 207.460 ;
        RECT 20.650 206.580 20.990 208.440 ;
        RECT 21.430 207.560 22.510 207.900 ;
        RECT 14.530 206.240 20.990 206.580 ;
        RECT 13.150 205.800 14.230 206.140 ;
        RECT 21.430 205.800 22.510 206.140 ;
        RECT 15.310 205.360 16.390 205.700 ;
        RECT 19.270 205.360 20.350 205.700 ;
        RECT 20.650 205.460 21.730 205.800 ;
        RECT 20.650 204.820 20.990 205.460 ;
        RECT 15.310 204.480 20.990 204.820 ;
        RECT 13.150 204.040 14.230 204.380 ;
        RECT 21.430 204.040 22.510 204.380 ;
        RECT 15.310 203.600 16.390 203.940 ;
        RECT 19.270 203.600 20.350 203.940 ;
        RECT 14.530 202.720 16.390 203.060 ;
        RECT 19.270 202.720 20.990 203.060 ;
        RECT 14.530 202.620 14.870 202.720 ;
        RECT 10.990 202.280 14.870 202.620 ;
        RECT 10.990 201.350 12.070 202.280 ;
        RECT 14.530 202.180 14.870 202.280 ;
        RECT 20.650 202.620 20.990 202.720 ;
        RECT 23.590 202.620 24.670 221.150 ;
        RECT 27.910 220.320 32.950 220.660 ;
        RECT 25.750 219.880 26.830 220.220 ;
        RECT 33.390 219.880 35.110 220.220 ;
        RECT 27.910 219.440 28.990 219.780 ;
        RECT 31.870 219.440 32.950 219.780 ;
        RECT 33.390 218.900 33.730 219.880 ;
        RECT 27.910 218.560 33.730 218.900 ;
        RECT 25.750 218.120 27.610 218.460 ;
        RECT 25.750 217.240 26.830 217.580 ;
        RECT 25.750 215.480 26.830 215.820 ;
        RECT 25.750 214.600 26.830 214.940 ;
        RECT 25.750 212.840 26.830 213.180 ;
        RECT 25.750 211.080 26.830 211.420 ;
        RECT 25.750 210.200 26.830 210.540 ;
        RECT 27.270 208.780 27.610 218.120 ;
        RECT 27.910 217.680 28.990 218.020 ;
        RECT 27.910 216.800 28.990 217.140 ;
        RECT 31.230 216.260 31.570 218.560 ;
        RECT 34.030 218.120 35.110 218.460 ;
        RECT 31.870 217.680 32.950 218.020 ;
        RECT 34.030 217.240 35.110 217.580 ;
        RECT 31.870 216.800 32.950 217.140 ;
        RECT 27.910 215.920 32.950 216.260 ;
        RECT 34.030 215.480 35.110 215.820 ;
        RECT 27.910 215.040 28.990 215.380 ;
        RECT 31.870 215.040 32.950 215.380 ;
        RECT 33.390 215.140 34.330 215.480 ;
        RECT 27.910 214.160 28.990 214.500 ;
        RECT 31.870 214.160 32.950 214.500 ;
        RECT 27.910 213.280 32.950 213.620 ;
        RECT 27.910 212.400 28.990 212.740 ;
        RECT 31.870 212.400 32.950 212.740 ;
        RECT 27.910 211.520 32.950 211.860 ;
        RECT 27.910 210.640 28.990 210.980 ;
        RECT 27.910 209.760 28.990 210.100 ;
        RECT 31.230 209.220 31.570 211.520 ;
        RECT 33.390 211.420 33.730 215.140 ;
        RECT 34.030 214.600 35.110 214.940 ;
        RECT 34.030 212.840 35.110 213.180 ;
        RECT 33.390 211.080 35.110 211.420 ;
        RECT 31.870 210.640 32.950 210.980 ;
        RECT 31.870 209.760 32.950 210.100 ;
        RECT 27.910 208.880 32.950 209.220 ;
        RECT 25.750 208.440 27.610 208.780 ;
        RECT 25.750 207.560 26.830 207.900 ;
        RECT 27.270 206.580 27.610 208.440 ;
        RECT 27.910 208.000 28.990 208.340 ;
        RECT 31.870 208.000 32.950 208.340 ;
        RECT 27.910 207.120 28.990 207.460 ;
        RECT 31.870 207.120 32.950 207.460 ;
        RECT 33.390 206.580 33.730 211.080 ;
        RECT 34.030 210.200 35.110 210.540 ;
        RECT 34.030 208.440 35.110 208.780 ;
        RECT 34.030 207.560 35.110 207.900 ;
        RECT 27.270 206.240 33.730 206.580 ;
        RECT 25.750 205.800 26.830 206.140 ;
        RECT 34.030 205.800 35.110 206.140 ;
        RECT 26.530 205.460 27.610 205.800 ;
        RECT 27.270 204.820 27.610 205.460 ;
        RECT 27.910 205.360 28.990 205.700 ;
        RECT 31.870 205.360 32.950 205.700 ;
        RECT 27.270 204.480 32.950 204.820 ;
        RECT 25.750 204.040 26.830 204.380 ;
        RECT 34.030 204.040 35.110 204.380 ;
        RECT 27.910 203.600 28.990 203.940 ;
        RECT 31.870 203.600 32.950 203.940 ;
        RECT 27.270 202.720 28.990 203.060 ;
        RECT 31.870 202.720 33.730 203.060 ;
        RECT 27.270 202.620 27.610 202.720 ;
        RECT 20.650 202.280 27.610 202.620 ;
        RECT 20.650 202.180 20.990 202.280 ;
        RECT 14.530 201.840 16.390 202.180 ;
        RECT 19.270 201.840 20.990 202.180 ;
        RECT 23.590 201.350 24.670 202.280 ;
        RECT 27.270 202.180 27.610 202.280 ;
        RECT 33.390 202.620 33.730 202.720 ;
        RECT 36.190 202.620 37.270 221.150 ;
        RECT 40.510 220.320 45.550 220.660 ;
        RECT 38.350 219.880 40.070 220.220 ;
        RECT 46.630 219.880 47.710 220.220 ;
        RECT 39.730 218.900 40.070 219.880 ;
        RECT 40.510 219.440 41.590 219.780 ;
        RECT 44.470 219.440 45.550 219.780 ;
        RECT 39.730 218.560 45.550 218.900 ;
        RECT 38.350 218.120 39.430 218.460 ;
        RECT 40.510 217.680 41.590 218.020 ;
        RECT 38.350 217.240 39.430 217.580 ;
        RECT 40.510 216.800 41.590 217.140 ;
        RECT 41.890 216.260 42.230 218.560 ;
        RECT 45.850 218.120 47.710 218.460 ;
        RECT 44.470 217.680 45.550 218.020 ;
        RECT 44.470 216.800 45.550 217.140 ;
        RECT 40.510 215.920 45.550 216.260 ;
        RECT 38.350 215.480 39.430 215.820 ;
        RECT 39.130 215.140 40.070 215.480 ;
        RECT 38.350 214.600 39.430 214.940 ;
        RECT 38.350 212.840 39.430 213.180 ;
        RECT 39.730 211.420 40.070 215.140 ;
        RECT 40.510 215.040 41.590 215.380 ;
        RECT 44.470 215.040 45.550 215.380 ;
        RECT 40.510 214.160 41.590 214.500 ;
        RECT 44.470 214.160 45.550 214.500 ;
        RECT 40.510 213.280 45.550 213.620 ;
        RECT 40.510 212.400 41.590 212.740 ;
        RECT 44.470 212.400 45.550 212.740 ;
        RECT 40.510 211.520 45.550 211.860 ;
        RECT 38.350 211.080 40.070 211.420 ;
        RECT 38.350 210.200 39.430 210.540 ;
        RECT 38.350 208.440 39.430 208.780 ;
        RECT 38.350 207.560 39.430 207.900 ;
        RECT 39.730 206.580 40.070 211.080 ;
        RECT 40.510 210.640 41.590 210.980 ;
        RECT 40.510 209.760 41.590 210.100 ;
        RECT 41.890 209.220 42.230 211.520 ;
        RECT 44.470 210.640 45.550 210.980 ;
        RECT 44.470 209.760 45.550 210.100 ;
        RECT 40.510 208.880 45.550 209.220 ;
        RECT 45.850 208.780 46.190 218.120 ;
        RECT 46.630 217.240 47.710 217.580 ;
        RECT 46.630 215.480 47.710 215.820 ;
        RECT 46.630 214.600 47.710 214.940 ;
        RECT 46.630 212.840 47.710 213.180 ;
        RECT 46.630 211.080 47.710 211.420 ;
        RECT 46.630 210.200 47.710 210.540 ;
        RECT 45.850 208.440 47.710 208.780 ;
        RECT 40.510 208.000 41.590 208.340 ;
        RECT 44.470 208.000 45.550 208.340 ;
        RECT 40.510 207.120 41.590 207.460 ;
        RECT 44.470 207.120 45.550 207.460 ;
        RECT 45.850 206.580 46.190 208.440 ;
        RECT 46.630 207.560 47.710 207.900 ;
        RECT 39.730 206.240 46.190 206.580 ;
        RECT 38.350 205.800 39.430 206.140 ;
        RECT 46.630 205.800 47.710 206.140 ;
        RECT 40.510 205.360 41.590 205.700 ;
        RECT 44.470 205.360 45.550 205.700 ;
        RECT 45.850 205.460 46.930 205.800 ;
        RECT 45.850 204.820 46.190 205.460 ;
        RECT 40.510 204.480 46.190 204.820 ;
        RECT 38.350 204.040 39.430 204.380 ;
        RECT 46.630 204.040 47.710 204.380 ;
        RECT 40.510 203.600 41.590 203.940 ;
        RECT 44.470 203.600 45.550 203.940 ;
        RECT 39.730 202.720 41.590 203.060 ;
        RECT 44.470 202.720 46.190 203.060 ;
        RECT 39.730 202.620 40.070 202.720 ;
        RECT 33.390 202.280 40.070 202.620 ;
        RECT 33.390 202.180 33.730 202.280 ;
        RECT 27.270 201.840 28.990 202.180 ;
        RECT 31.870 201.840 33.730 202.180 ;
        RECT 36.190 201.350 37.270 202.280 ;
        RECT 39.730 202.180 40.070 202.280 ;
        RECT 45.850 202.620 46.190 202.720 ;
        RECT 48.790 202.620 49.870 221.150 ;
        RECT 53.110 220.320 58.150 220.660 ;
        RECT 50.950 219.880 52.030 220.220 ;
        RECT 58.590 219.880 60.310 220.220 ;
        RECT 53.110 219.440 54.190 219.780 ;
        RECT 57.070 219.440 58.150 219.780 ;
        RECT 58.590 218.900 58.930 219.880 ;
        RECT 53.110 218.560 58.930 218.900 ;
        RECT 50.950 218.120 52.810 218.460 ;
        RECT 50.950 217.240 52.030 217.580 ;
        RECT 50.950 215.480 52.030 215.820 ;
        RECT 50.950 214.600 52.030 214.940 ;
        RECT 50.950 212.840 52.030 213.180 ;
        RECT 50.950 211.080 52.030 211.420 ;
        RECT 50.950 210.200 52.030 210.540 ;
        RECT 52.470 208.780 52.810 218.120 ;
        RECT 53.110 217.680 54.190 218.020 ;
        RECT 53.110 216.800 54.190 217.140 ;
        RECT 56.430 216.260 56.770 218.560 ;
        RECT 59.230 218.120 60.310 218.460 ;
        RECT 57.070 217.680 58.150 218.020 ;
        RECT 59.230 217.240 60.310 217.580 ;
        RECT 57.070 216.800 58.150 217.140 ;
        RECT 53.110 215.920 58.150 216.260 ;
        RECT 59.230 215.480 60.310 215.820 ;
        RECT 53.110 215.040 54.190 215.380 ;
        RECT 57.070 215.040 58.150 215.380 ;
        RECT 58.590 215.140 59.530 215.480 ;
        RECT 53.110 214.160 54.190 214.500 ;
        RECT 57.070 214.160 58.150 214.500 ;
        RECT 53.110 213.280 58.150 213.620 ;
        RECT 53.110 212.400 54.190 212.740 ;
        RECT 57.070 212.400 58.150 212.740 ;
        RECT 53.110 211.520 58.150 211.860 ;
        RECT 53.110 210.640 54.190 210.980 ;
        RECT 53.110 209.760 54.190 210.100 ;
        RECT 56.430 209.220 56.770 211.520 ;
        RECT 58.590 211.420 58.930 215.140 ;
        RECT 59.230 214.600 60.310 214.940 ;
        RECT 59.230 212.840 60.310 213.180 ;
        RECT 58.590 211.080 60.310 211.420 ;
        RECT 57.070 210.640 58.150 210.980 ;
        RECT 57.070 209.760 58.150 210.100 ;
        RECT 53.110 208.880 58.150 209.220 ;
        RECT 50.950 208.440 52.810 208.780 ;
        RECT 50.950 207.560 52.030 207.900 ;
        RECT 52.470 206.580 52.810 208.440 ;
        RECT 53.110 208.000 54.190 208.340 ;
        RECT 57.070 208.000 58.150 208.340 ;
        RECT 53.110 207.120 54.190 207.460 ;
        RECT 57.070 207.120 58.150 207.460 ;
        RECT 58.590 206.580 58.930 211.080 ;
        RECT 59.230 210.200 60.310 210.540 ;
        RECT 59.230 208.440 60.310 208.780 ;
        RECT 59.230 207.560 60.310 207.900 ;
        RECT 52.470 206.240 58.930 206.580 ;
        RECT 50.950 205.800 52.030 206.140 ;
        RECT 59.230 205.800 60.310 206.140 ;
        RECT 51.730 205.460 52.810 205.800 ;
        RECT 52.470 204.820 52.810 205.460 ;
        RECT 53.110 205.360 54.190 205.700 ;
        RECT 57.070 205.360 58.150 205.700 ;
        RECT 52.470 204.480 58.150 204.820 ;
        RECT 50.950 204.040 52.030 204.380 ;
        RECT 59.230 204.040 60.310 204.380 ;
        RECT 53.110 203.600 54.190 203.940 ;
        RECT 57.070 203.600 58.150 203.940 ;
        RECT 52.470 202.720 54.190 203.060 ;
        RECT 57.070 202.720 58.930 203.060 ;
        RECT 52.470 202.620 52.810 202.720 ;
        RECT 45.850 202.280 52.810 202.620 ;
        RECT 45.850 202.180 46.190 202.280 ;
        RECT 39.730 201.840 41.590 202.180 ;
        RECT 44.470 201.840 46.190 202.180 ;
        RECT 48.790 201.350 49.870 202.280 ;
        RECT 52.470 202.180 52.810 202.280 ;
        RECT 58.590 202.620 58.930 202.720 ;
        RECT 61.390 202.620 62.470 221.150 ;
        RECT 65.710 220.320 70.750 220.660 ;
        RECT 63.550 219.880 65.270 220.220 ;
        RECT 71.830 219.880 72.910 220.220 ;
        RECT 64.930 218.900 65.270 219.880 ;
        RECT 65.710 219.440 66.790 219.780 ;
        RECT 69.670 219.440 70.750 219.780 ;
        RECT 64.930 218.560 70.750 218.900 ;
        RECT 63.550 218.120 64.630 218.460 ;
        RECT 65.710 217.680 66.790 218.020 ;
        RECT 63.550 217.240 64.630 217.580 ;
        RECT 65.710 216.800 66.790 217.140 ;
        RECT 67.090 216.260 67.430 218.560 ;
        RECT 71.050 218.120 72.910 218.460 ;
        RECT 69.670 217.680 70.750 218.020 ;
        RECT 69.670 216.800 70.750 217.140 ;
        RECT 65.710 215.920 70.750 216.260 ;
        RECT 63.550 215.480 64.630 215.820 ;
        RECT 64.330 215.140 65.270 215.480 ;
        RECT 63.550 214.600 64.630 214.940 ;
        RECT 63.550 212.840 64.630 213.180 ;
        RECT 64.930 211.420 65.270 215.140 ;
        RECT 65.710 215.040 66.790 215.380 ;
        RECT 69.670 215.040 70.750 215.380 ;
        RECT 65.710 214.160 66.790 214.500 ;
        RECT 69.670 214.160 70.750 214.500 ;
        RECT 65.710 213.280 70.750 213.620 ;
        RECT 65.710 212.400 66.790 212.740 ;
        RECT 69.670 212.400 70.750 212.740 ;
        RECT 65.710 211.520 70.750 211.860 ;
        RECT 63.550 211.080 65.270 211.420 ;
        RECT 63.550 210.200 64.630 210.540 ;
        RECT 63.550 208.440 64.630 208.780 ;
        RECT 63.550 207.560 64.630 207.900 ;
        RECT 64.930 206.580 65.270 211.080 ;
        RECT 65.710 210.640 66.790 210.980 ;
        RECT 65.710 209.760 66.790 210.100 ;
        RECT 67.090 209.220 67.430 211.520 ;
        RECT 69.670 210.640 70.750 210.980 ;
        RECT 69.670 209.760 70.750 210.100 ;
        RECT 65.710 208.880 70.750 209.220 ;
        RECT 71.050 208.780 71.390 218.120 ;
        RECT 71.830 217.240 72.910 217.580 ;
        RECT 71.830 215.480 72.910 215.820 ;
        RECT 71.830 214.600 72.910 214.940 ;
        RECT 71.830 212.840 72.910 213.180 ;
        RECT 71.830 211.080 72.910 211.420 ;
        RECT 71.830 210.200 72.910 210.540 ;
        RECT 71.050 208.440 72.910 208.780 ;
        RECT 65.710 208.000 66.790 208.340 ;
        RECT 69.670 208.000 70.750 208.340 ;
        RECT 65.710 207.120 66.790 207.460 ;
        RECT 69.670 207.120 70.750 207.460 ;
        RECT 71.050 206.580 71.390 208.440 ;
        RECT 71.830 207.560 72.910 207.900 ;
        RECT 64.930 206.240 71.390 206.580 ;
        RECT 63.550 205.800 64.630 206.140 ;
        RECT 71.830 205.800 72.910 206.140 ;
        RECT 65.710 205.360 66.790 205.700 ;
        RECT 69.670 205.360 70.750 205.700 ;
        RECT 71.050 205.460 72.130 205.800 ;
        RECT 71.050 204.820 71.390 205.460 ;
        RECT 65.710 204.480 71.390 204.820 ;
        RECT 63.550 204.040 64.630 204.380 ;
        RECT 71.830 204.040 72.910 204.380 ;
        RECT 65.710 203.600 66.790 203.940 ;
        RECT 69.670 203.600 70.750 203.940 ;
        RECT 64.930 202.720 66.790 203.060 ;
        RECT 69.670 202.720 71.390 203.060 ;
        RECT 64.930 202.620 65.270 202.720 ;
        RECT 58.590 202.280 65.270 202.620 ;
        RECT 58.590 202.180 58.930 202.280 ;
        RECT 52.470 201.840 54.190 202.180 ;
        RECT 57.070 201.840 58.930 202.180 ;
        RECT 61.390 201.350 62.470 202.280 ;
        RECT 64.930 202.180 65.270 202.280 ;
        RECT 71.050 202.620 71.390 202.720 ;
        RECT 73.990 202.620 75.070 221.150 ;
        RECT 78.310 220.320 83.350 220.660 ;
        RECT 76.150 219.880 77.230 220.220 ;
        RECT 83.790 219.880 85.510 220.220 ;
        RECT 78.310 219.440 79.390 219.780 ;
        RECT 82.270 219.440 83.350 219.780 ;
        RECT 83.790 218.900 84.130 219.880 ;
        RECT 78.310 218.560 84.130 218.900 ;
        RECT 76.150 218.120 78.010 218.460 ;
        RECT 76.150 217.240 77.230 217.580 ;
        RECT 76.150 215.480 77.230 215.820 ;
        RECT 76.150 214.600 77.230 214.940 ;
        RECT 76.150 212.840 77.230 213.180 ;
        RECT 76.150 211.080 77.230 211.420 ;
        RECT 76.150 210.200 77.230 210.540 ;
        RECT 77.670 208.780 78.010 218.120 ;
        RECT 78.310 217.680 79.390 218.020 ;
        RECT 78.310 216.800 79.390 217.140 ;
        RECT 81.630 216.260 81.970 218.560 ;
        RECT 84.430 218.120 85.510 218.460 ;
        RECT 82.270 217.680 83.350 218.020 ;
        RECT 84.430 217.240 85.510 217.580 ;
        RECT 82.270 216.800 83.350 217.140 ;
        RECT 78.310 215.920 83.350 216.260 ;
        RECT 84.430 215.480 85.510 215.820 ;
        RECT 78.310 215.040 79.390 215.380 ;
        RECT 82.270 215.040 83.350 215.380 ;
        RECT 83.790 215.140 84.730 215.480 ;
        RECT 78.310 214.160 79.390 214.500 ;
        RECT 82.270 214.160 83.350 214.500 ;
        RECT 78.310 213.280 83.350 213.620 ;
        RECT 78.310 212.400 79.390 212.740 ;
        RECT 82.270 212.400 83.350 212.740 ;
        RECT 78.310 211.520 83.350 211.860 ;
        RECT 78.310 210.640 79.390 210.980 ;
        RECT 78.310 209.760 79.390 210.100 ;
        RECT 81.630 209.220 81.970 211.520 ;
        RECT 83.790 211.420 84.130 215.140 ;
        RECT 84.430 214.600 85.510 214.940 ;
        RECT 84.430 212.840 85.510 213.180 ;
        RECT 83.790 211.080 85.510 211.420 ;
        RECT 82.270 210.640 83.350 210.980 ;
        RECT 82.270 209.760 83.350 210.100 ;
        RECT 78.310 208.880 83.350 209.220 ;
        RECT 76.150 208.440 78.010 208.780 ;
        RECT 76.150 207.560 77.230 207.900 ;
        RECT 77.670 206.580 78.010 208.440 ;
        RECT 78.310 208.000 79.390 208.340 ;
        RECT 82.270 208.000 83.350 208.340 ;
        RECT 78.310 207.120 79.390 207.460 ;
        RECT 82.270 207.120 83.350 207.460 ;
        RECT 83.790 206.580 84.130 211.080 ;
        RECT 84.430 210.200 85.510 210.540 ;
        RECT 84.430 208.440 85.510 208.780 ;
        RECT 84.430 207.560 85.510 207.900 ;
        RECT 77.670 206.240 84.130 206.580 ;
        RECT 76.150 205.800 77.230 206.140 ;
        RECT 84.430 205.800 85.510 206.140 ;
        RECT 76.930 205.460 78.010 205.800 ;
        RECT 77.670 204.820 78.010 205.460 ;
        RECT 78.310 205.360 79.390 205.700 ;
        RECT 82.270 205.360 83.350 205.700 ;
        RECT 77.670 204.480 83.350 204.820 ;
        RECT 76.150 204.040 77.230 204.380 ;
        RECT 84.430 204.040 85.510 204.380 ;
        RECT 78.310 203.600 79.390 203.940 ;
        RECT 82.270 203.600 83.350 203.940 ;
        RECT 77.670 202.720 79.390 203.060 ;
        RECT 82.270 202.720 84.130 203.060 ;
        RECT 77.670 202.620 78.010 202.720 ;
        RECT 71.050 202.280 78.010 202.620 ;
        RECT 71.050 202.180 71.390 202.280 ;
        RECT 64.930 201.840 66.790 202.180 ;
        RECT 69.670 201.840 71.390 202.180 ;
        RECT 73.990 201.350 75.070 202.280 ;
        RECT 77.670 202.180 78.010 202.280 ;
        RECT 83.790 202.620 84.130 202.720 ;
        RECT 86.590 202.620 87.670 221.150 ;
        RECT 90.910 220.320 95.950 220.660 ;
        RECT 88.750 219.880 90.470 220.220 ;
        RECT 97.030 219.880 98.110 220.220 ;
        RECT 90.130 218.900 90.470 219.880 ;
        RECT 90.910 219.440 91.990 219.780 ;
        RECT 94.870 219.440 95.950 219.780 ;
        RECT 90.130 218.560 95.950 218.900 ;
        RECT 88.750 218.120 89.830 218.460 ;
        RECT 90.910 217.680 91.990 218.020 ;
        RECT 88.750 217.240 89.830 217.580 ;
        RECT 90.910 216.800 91.990 217.140 ;
        RECT 92.290 216.260 92.630 218.560 ;
        RECT 96.250 218.120 98.110 218.460 ;
        RECT 94.870 217.680 95.950 218.020 ;
        RECT 94.870 216.800 95.950 217.140 ;
        RECT 90.910 215.920 95.950 216.260 ;
        RECT 88.750 215.480 89.830 215.820 ;
        RECT 89.530 215.140 90.470 215.480 ;
        RECT 88.750 214.600 89.830 214.940 ;
        RECT 88.750 212.840 89.830 213.180 ;
        RECT 90.130 211.420 90.470 215.140 ;
        RECT 90.910 215.040 91.990 215.380 ;
        RECT 94.870 215.040 95.950 215.380 ;
        RECT 90.910 214.160 91.990 214.500 ;
        RECT 94.870 214.160 95.950 214.500 ;
        RECT 90.910 213.280 95.950 213.620 ;
        RECT 90.910 212.400 91.990 212.740 ;
        RECT 94.870 212.400 95.950 212.740 ;
        RECT 90.910 211.520 95.950 211.860 ;
        RECT 88.750 211.080 90.470 211.420 ;
        RECT 88.750 210.200 89.830 210.540 ;
        RECT 88.750 208.440 89.830 208.780 ;
        RECT 88.750 207.560 89.830 207.900 ;
        RECT 90.130 206.580 90.470 211.080 ;
        RECT 90.910 210.640 91.990 210.980 ;
        RECT 90.910 209.760 91.990 210.100 ;
        RECT 92.290 209.220 92.630 211.520 ;
        RECT 94.870 210.640 95.950 210.980 ;
        RECT 94.870 209.760 95.950 210.100 ;
        RECT 90.910 208.880 95.950 209.220 ;
        RECT 96.250 208.780 96.590 218.120 ;
        RECT 97.030 217.240 98.110 217.580 ;
        RECT 97.030 215.480 98.110 215.820 ;
        RECT 97.030 214.600 98.110 214.940 ;
        RECT 97.030 212.840 98.110 213.180 ;
        RECT 97.030 211.080 98.110 211.420 ;
        RECT 97.030 210.200 98.110 210.540 ;
        RECT 96.250 208.440 98.110 208.780 ;
        RECT 90.910 208.000 91.990 208.340 ;
        RECT 94.870 208.000 95.950 208.340 ;
        RECT 90.910 207.120 91.990 207.460 ;
        RECT 94.870 207.120 95.950 207.460 ;
        RECT 96.250 206.580 96.590 208.440 ;
        RECT 97.030 207.560 98.110 207.900 ;
        RECT 90.130 206.240 96.590 206.580 ;
        RECT 88.750 205.800 89.830 206.140 ;
        RECT 97.030 205.800 98.110 206.140 ;
        RECT 90.910 205.360 91.990 205.700 ;
        RECT 94.870 205.360 95.950 205.700 ;
        RECT 96.250 205.460 97.330 205.800 ;
        RECT 96.250 204.820 96.590 205.460 ;
        RECT 90.910 204.480 96.590 204.820 ;
        RECT 88.750 204.040 89.830 204.380 ;
        RECT 97.030 204.040 98.110 204.380 ;
        RECT 90.910 203.600 91.990 203.940 ;
        RECT 94.870 203.600 95.950 203.940 ;
        RECT 90.130 202.720 91.990 203.060 ;
        RECT 94.870 202.720 96.590 203.060 ;
        RECT 90.130 202.620 90.470 202.720 ;
        RECT 83.790 202.280 90.470 202.620 ;
        RECT 83.790 202.180 84.130 202.280 ;
        RECT 77.670 201.840 79.390 202.180 ;
        RECT 82.270 201.840 84.130 202.180 ;
        RECT 86.590 201.350 87.670 202.280 ;
        RECT 90.130 202.180 90.470 202.280 ;
        RECT 96.250 202.620 96.590 202.720 ;
        RECT 99.190 202.620 100.270 221.150 ;
        RECT 103.510 220.320 108.550 220.660 ;
        RECT 101.350 219.880 102.430 220.220 ;
        RECT 108.990 219.880 110.710 220.220 ;
        RECT 103.510 219.440 104.590 219.780 ;
        RECT 107.470 219.440 108.550 219.780 ;
        RECT 108.990 218.900 109.330 219.880 ;
        RECT 103.510 218.560 109.330 218.900 ;
        RECT 101.350 218.120 103.210 218.460 ;
        RECT 101.350 217.240 102.430 217.580 ;
        RECT 101.350 215.480 102.430 215.820 ;
        RECT 101.350 214.600 102.430 214.940 ;
        RECT 101.350 212.840 102.430 213.180 ;
        RECT 101.350 211.080 102.430 211.420 ;
        RECT 101.350 210.200 102.430 210.540 ;
        RECT 102.870 208.780 103.210 218.120 ;
        RECT 103.510 217.680 104.590 218.020 ;
        RECT 103.510 216.800 104.590 217.140 ;
        RECT 106.830 216.260 107.170 218.560 ;
        RECT 109.630 218.120 110.710 218.460 ;
        RECT 107.470 217.680 108.550 218.020 ;
        RECT 109.630 217.240 110.710 217.580 ;
        RECT 107.470 216.800 108.550 217.140 ;
        RECT 103.510 215.920 108.550 216.260 ;
        RECT 109.630 215.480 110.710 215.820 ;
        RECT 103.510 215.040 104.590 215.380 ;
        RECT 107.470 215.040 108.550 215.380 ;
        RECT 108.990 215.140 109.930 215.480 ;
        RECT 103.510 214.160 104.590 214.500 ;
        RECT 107.470 214.160 108.550 214.500 ;
        RECT 103.510 213.280 108.550 213.620 ;
        RECT 103.510 212.400 104.590 212.740 ;
        RECT 107.470 212.400 108.550 212.740 ;
        RECT 103.510 211.520 108.550 211.860 ;
        RECT 103.510 210.640 104.590 210.980 ;
        RECT 103.510 209.760 104.590 210.100 ;
        RECT 106.830 209.220 107.170 211.520 ;
        RECT 108.990 211.420 109.330 215.140 ;
        RECT 109.630 214.600 110.710 214.940 ;
        RECT 109.630 212.840 110.710 213.180 ;
        RECT 108.990 211.080 110.710 211.420 ;
        RECT 107.470 210.640 108.550 210.980 ;
        RECT 107.470 209.760 108.550 210.100 ;
        RECT 103.510 208.880 108.550 209.220 ;
        RECT 101.350 208.440 103.210 208.780 ;
        RECT 101.350 207.560 102.430 207.900 ;
        RECT 102.870 206.580 103.210 208.440 ;
        RECT 103.510 208.000 104.590 208.340 ;
        RECT 107.470 208.000 108.550 208.340 ;
        RECT 103.510 207.120 104.590 207.460 ;
        RECT 107.470 207.120 108.550 207.460 ;
        RECT 108.990 206.580 109.330 211.080 ;
        RECT 109.630 210.200 110.710 210.540 ;
        RECT 109.630 208.440 110.710 208.780 ;
        RECT 109.630 207.560 110.710 207.900 ;
        RECT 102.870 206.240 109.330 206.580 ;
        RECT 101.350 205.800 102.430 206.140 ;
        RECT 109.630 205.800 110.710 206.140 ;
        RECT 102.130 205.460 103.210 205.800 ;
        RECT 102.870 204.820 103.210 205.460 ;
        RECT 103.510 205.360 104.590 205.700 ;
        RECT 107.470 205.360 108.550 205.700 ;
        RECT 102.870 204.480 108.550 204.820 ;
        RECT 101.350 204.040 102.430 204.380 ;
        RECT 109.630 204.040 110.710 204.380 ;
        RECT 103.510 203.600 104.590 203.940 ;
        RECT 107.470 203.600 108.550 203.940 ;
        RECT 102.870 202.720 104.590 203.060 ;
        RECT 107.470 202.720 109.330 203.060 ;
        RECT 102.870 202.620 103.210 202.720 ;
        RECT 96.250 202.280 103.210 202.620 ;
        RECT 96.250 202.180 96.590 202.280 ;
        RECT 90.130 201.840 91.990 202.180 ;
        RECT 94.870 201.840 96.590 202.180 ;
        RECT 99.190 201.350 100.270 202.280 ;
        RECT 102.870 202.180 103.210 202.280 ;
        RECT 108.990 202.620 109.330 202.720 ;
        RECT 111.790 202.620 112.870 222.030 ;
        RECT 116.110 221.200 117.190 221.540 ;
        RECT 120.070 221.200 121.790 221.540 ;
        RECT 121.450 221.100 121.790 221.200 ;
        RECT 113.950 220.760 115.030 221.100 ;
        RECT 121.450 220.760 123.310 221.100 ;
        RECT 116.110 220.320 117.190 220.660 ;
        RECT 120.070 220.320 121.150 220.660 ;
        RECT 116.110 219.440 121.150 219.780 ;
        RECT 113.950 219.000 115.670 219.340 ;
        RECT 122.230 219.000 123.310 219.340 ;
        RECT 115.330 218.020 115.670 219.000 ;
        RECT 116.110 218.560 117.190 218.900 ;
        RECT 120.070 218.560 121.150 218.900 ;
        RECT 115.330 217.680 117.830 218.020 ;
        RECT 120.070 217.680 121.150 218.020 ;
        RECT 113.950 217.240 115.030 217.580 ;
        RECT 117.490 217.140 117.830 217.680 ;
        RECT 122.230 217.240 123.310 217.580 ;
        RECT 116.110 216.800 117.190 217.140 ;
        RECT 117.490 216.800 121.150 217.140 ;
        RECT 113.950 216.360 115.030 216.700 ;
        RECT 122.230 216.360 123.310 216.700 ;
        RECT 116.110 215.920 117.190 216.260 ;
        RECT 120.070 215.920 121.150 216.260 ;
        RECT 116.110 215.040 121.150 215.380 ;
        RECT 113.950 214.600 115.810 214.940 ;
        RECT 122.230 214.600 123.310 214.940 ;
        RECT 115.470 213.960 115.810 214.600 ;
        RECT 116.110 214.160 117.190 214.500 ;
        RECT 120.070 214.160 121.150 214.500 ;
        RECT 115.470 213.620 116.410 213.960 ;
        RECT 116.110 213.280 121.150 213.620 ;
        RECT 113.950 212.840 115.670 213.180 ;
        RECT 122.230 212.840 123.310 213.180 ;
        RECT 113.950 211.080 115.030 211.420 ;
        RECT 115.330 210.980 115.670 212.840 ;
        RECT 116.110 212.400 117.190 212.740 ;
        RECT 120.070 212.400 121.150 212.740 ;
        RECT 116.110 211.520 117.190 211.860 ;
        RECT 117.490 211.520 121.150 211.860 ;
        RECT 117.490 210.980 117.830 211.520 ;
        RECT 122.230 211.080 123.310 211.420 ;
        RECT 115.330 210.640 117.830 210.980 ;
        RECT 120.070 210.640 121.150 210.980 ;
        RECT 113.950 210.200 115.030 210.540 ;
        RECT 122.230 210.200 123.310 210.540 ;
        RECT 116.110 209.760 117.190 210.100 ;
        RECT 120.070 209.760 121.150 210.100 ;
        RECT 116.110 208.880 121.150 209.220 ;
        RECT 113.950 208.440 115.670 208.780 ;
        RECT 122.230 208.440 123.310 208.780 ;
        RECT 113.950 207.560 115.030 207.900 ;
        RECT 115.330 207.460 115.670 208.440 ;
        RECT 116.110 208.000 117.190 208.340 ;
        RECT 120.070 208.000 121.150 208.340 ;
        RECT 122.230 207.560 123.310 207.900 ;
        RECT 115.330 207.120 121.150 207.460 ;
        RECT 116.110 206.240 121.150 206.580 ;
        RECT 113.950 205.800 115.030 206.140 ;
        RECT 122.230 205.800 123.310 206.140 ;
        RECT 116.110 205.360 117.190 205.700 ;
        RECT 120.070 205.360 121.150 205.700 ;
        RECT 116.110 204.480 121.150 204.820 ;
        RECT 113.950 204.040 115.030 204.380 ;
        RECT 122.230 204.040 123.310 204.380 ;
        RECT 116.110 203.600 117.190 203.940 ;
        RECT 120.070 203.600 121.150 203.940 ;
        RECT 115.330 202.720 117.190 203.060 ;
        RECT 120.070 202.720 121.790 203.060 ;
        RECT 115.330 202.620 115.670 202.720 ;
        RECT 108.990 202.280 115.670 202.620 ;
        RECT 108.990 202.180 109.330 202.280 ;
        RECT 102.870 201.840 104.590 202.180 ;
        RECT 107.470 201.840 109.330 202.180 ;
        RECT 111.790 201.350 112.870 202.280 ;
        RECT 115.330 202.180 115.670 202.280 ;
        RECT 121.450 202.620 121.790 202.720 ;
        RECT 124.390 202.620 125.470 222.030 ;
        RECT 121.450 202.280 125.470 202.620 ;
        RECT 121.450 202.180 121.790 202.280 ;
        RECT 115.330 201.840 117.190 202.180 ;
        RECT 120.070 201.840 121.790 202.180 ;
        RECT 124.390 201.350 125.470 202.280 ;
        RECT 11.530 200.510 132.450 200.850 ;
        RECT 11.530 199.070 124.930 199.990 ;
        RECT 2.630 4.260 2.970 198.550 ;
        RECT 3.690 197.630 132.570 198.550 ;
        RECT 3.690 194.030 132.570 194.950 ;
        RECT 3.690 6.960 4.610 194.030 ;
        RECT 7.290 190.430 128.970 191.350 ;
        RECT 7.290 10.560 8.210 190.430 ;
        RECT 10.890 187.040 11.970 187.970 ;
        RECT 14.430 187.140 16.290 187.480 ;
        RECT 19.170 187.140 20.890 187.480 ;
        RECT 14.430 187.040 14.770 187.140 ;
        RECT 10.890 186.700 14.770 187.040 ;
        RECT 10.890 135.120 11.970 186.700 ;
        RECT 14.430 186.600 14.770 186.700 ;
        RECT 20.550 187.040 20.890 187.140 ;
        RECT 23.490 187.040 24.570 187.970 ;
        RECT 27.170 187.140 28.890 187.480 ;
        RECT 31.770 187.140 33.630 187.480 ;
        RECT 27.170 187.040 27.510 187.140 ;
        RECT 20.550 186.700 27.510 187.040 ;
        RECT 20.550 186.600 20.890 186.700 ;
        RECT 14.430 186.260 16.290 186.600 ;
        RECT 19.170 186.260 20.890 186.600 ;
        RECT 19.170 185.720 20.090 185.890 ;
        RECT 15.210 185.380 20.250 185.720 ;
        RECT 13.050 184.940 14.770 185.280 ;
        RECT 21.330 184.940 22.410 185.280 ;
        RECT 13.050 183.180 14.130 183.520 ;
        RECT 14.430 183.080 14.770 184.940 ;
        RECT 15.210 184.500 16.290 184.840 ;
        RECT 19.170 184.500 20.250 184.840 ;
        RECT 15.210 183.620 16.290 183.960 ;
        RECT 16.590 183.620 20.250 183.960 ;
        RECT 16.590 183.080 16.930 183.620 ;
        RECT 21.330 183.180 22.410 183.520 ;
        RECT 14.430 182.740 16.930 183.080 ;
        RECT 19.170 182.740 20.250 183.080 ;
        RECT 13.050 182.300 14.130 182.640 ;
        RECT 21.330 182.300 22.410 182.640 ;
        RECT 13.830 181.960 14.770 182.300 ;
        RECT 14.430 181.320 14.770 181.960 ;
        RECT 15.210 181.860 16.290 182.200 ;
        RECT 19.170 181.860 20.250 182.200 ;
        RECT 14.430 180.980 20.250 181.320 ;
        RECT 13.050 180.540 14.130 180.880 ;
        RECT 21.330 180.540 22.410 180.880 ;
        RECT 13.830 180.200 14.770 180.540 ;
        RECT 14.430 179.560 14.770 180.200 ;
        RECT 15.210 180.100 16.290 180.440 ;
        RECT 19.170 180.100 20.250 180.440 ;
        RECT 14.430 179.220 16.930 179.560 ;
        RECT 19.170 179.220 20.250 179.560 ;
        RECT 13.050 178.780 14.130 179.120 ;
        RECT 16.590 178.680 16.930 179.220 ;
        RECT 21.330 178.780 22.410 179.120 ;
        RECT 15.210 178.340 16.290 178.680 ;
        RECT 16.590 178.340 20.250 178.680 ;
        RECT 13.050 177.900 14.130 178.240 ;
        RECT 21.330 177.900 22.410 178.240 ;
        RECT 13.420 176.480 13.760 177.900 ;
        RECT 15.210 177.460 16.290 177.800 ;
        RECT 19.170 177.460 20.250 177.800 ;
        RECT 15.210 176.580 20.250 176.920 ;
        RECT 13.050 176.140 14.770 176.480 ;
        RECT 21.330 176.140 22.410 176.480 ;
        RECT 14.430 175.160 14.770 176.140 ;
        RECT 15.210 175.700 16.290 176.040 ;
        RECT 19.170 175.700 20.250 176.040 ;
        RECT 14.430 174.820 20.250 175.160 ;
        RECT 13.050 174.380 14.130 174.720 ;
        RECT 21.330 174.380 22.410 174.720 ;
        RECT 15.210 173.940 16.290 174.280 ;
        RECT 19.170 173.940 20.250 174.280 ;
        RECT 15.210 173.060 20.250 173.400 ;
        RECT 13.050 172.620 14.130 172.960 ;
        RECT 13.420 172.080 13.760 172.620 ;
        RECT 15.210 172.180 16.290 172.520 ;
        RECT 13.050 171.740 14.130 172.080 ;
        RECT 13.420 171.200 13.760 171.740 ;
        RECT 15.210 171.300 16.290 171.640 ;
        RECT 13.050 170.860 14.130 171.200 ;
        RECT 13.420 170.320 13.760 170.860 ;
        RECT 15.210 170.420 16.290 170.760 ;
        RECT 13.050 169.980 14.130 170.320 ;
        RECT 16.590 169.880 16.930 173.060 ;
        RECT 21.330 172.620 22.410 172.960 ;
        RECT 19.170 172.180 20.250 172.520 ;
        RECT 21.700 172.080 22.040 172.620 ;
        RECT 21.330 171.740 22.410 172.080 ;
        RECT 19.170 171.300 20.250 171.640 ;
        RECT 21.330 170.860 22.410 171.200 ;
        RECT 19.170 170.420 20.250 170.760 ;
        RECT 21.700 170.320 22.040 170.860 ;
        RECT 20.550 169.980 22.410 170.320 ;
        RECT 15.210 169.540 16.290 169.880 ;
        RECT 16.590 169.540 20.250 169.880 ;
        RECT 15.210 168.660 16.290 169.000 ;
        RECT 19.170 168.660 20.250 169.000 ;
        RECT 13.050 168.220 14.130 168.560 ;
        RECT 13.420 167.680 13.760 168.220 ;
        RECT 15.210 167.780 20.250 168.120 ;
        RECT 13.050 167.340 14.130 167.680 ;
        RECT 13.420 166.800 13.760 167.340 ;
        RECT 15.210 166.900 16.290 167.240 ;
        RECT 13.050 166.460 14.130 166.800 ;
        RECT 13.420 165.920 13.760 166.460 ;
        RECT 16.590 166.360 16.930 167.780 ;
        RECT 19.170 166.900 20.250 167.240 ;
        RECT 18.160 166.360 18.500 166.650 ;
        RECT 20.550 166.360 20.890 169.980 ;
        RECT 21.330 168.220 22.410 168.560 ;
        RECT 21.700 167.680 22.040 168.220 ;
        RECT 21.330 167.340 22.410 167.680 ;
        RECT 21.700 166.800 22.040 167.340 ;
        RECT 21.330 166.460 22.410 166.800 ;
        RECT 15.210 166.020 20.890 166.360 ;
        RECT 13.050 165.580 14.770 165.920 ;
        RECT 18.160 165.730 18.500 166.020 ;
        RECT 21.700 165.920 22.040 166.460 ;
        RECT 21.330 165.580 22.410 165.920 ;
        RECT 13.050 163.820 14.130 164.160 ;
        RECT 13.420 163.280 13.760 163.820 ;
        RECT 13.050 162.940 14.130 163.280 ;
        RECT 13.420 162.400 13.760 162.940 ;
        RECT 13.050 162.060 14.130 162.400 ;
        RECT 13.420 161.520 13.760 162.060 ;
        RECT 14.430 161.960 14.770 165.580 ;
        RECT 15.210 165.140 16.290 165.480 ;
        RECT 19.170 165.140 20.250 165.480 ;
        RECT 15.210 164.260 16.290 164.600 ;
        RECT 19.170 164.260 20.250 164.600 ;
        RECT 21.330 163.820 22.410 164.160 ;
        RECT 15.210 163.380 20.250 163.720 ;
        RECT 15.210 162.500 16.290 162.840 ;
        RECT 16.590 161.960 16.930 163.380 ;
        RECT 21.700 163.280 22.040 163.820 ;
        RECT 21.330 162.940 22.410 163.280 ;
        RECT 19.170 162.500 20.250 162.840 ;
        RECT 21.700 162.400 22.040 162.940 ;
        RECT 17.375 161.960 17.715 162.250 ;
        RECT 21.330 162.060 22.410 162.400 ;
        RECT 14.430 161.620 20.250 161.960 ;
        RECT 13.050 161.180 14.130 161.520 ;
        RECT 17.375 161.330 17.715 161.620 ;
        RECT 21.700 161.520 22.040 162.060 ;
        RECT 21.330 161.180 22.410 161.520 ;
        RECT 15.210 160.740 16.290 161.080 ;
        RECT 19.170 160.740 20.250 161.080 ;
        RECT 15.210 159.860 16.290 160.200 ;
        RECT 19.170 159.860 20.250 160.200 ;
        RECT 13.050 159.420 14.130 159.760 ;
        RECT 21.330 159.420 22.410 159.760 ;
        RECT 13.420 158.880 13.760 159.420 ;
        RECT 15.210 158.980 20.250 159.320 ;
        RECT 13.050 158.540 14.130 158.880 ;
        RECT 13.420 158.000 13.760 158.540 ;
        RECT 15.210 158.100 16.290 158.440 ;
        RECT 13.050 157.660 14.130 158.000 ;
        RECT 16.590 157.850 16.930 158.980 ;
        RECT 21.700 158.880 22.040 159.420 ;
        RECT 21.330 158.540 22.410 158.880 ;
        RECT 19.170 158.100 20.250 158.440 ;
        RECT 21.700 158.000 22.040 158.540 ;
        RECT 13.420 157.120 13.760 157.660 ;
        RECT 16.590 157.560 17.000 157.850 ;
        RECT 21.330 157.660 22.410 158.000 ;
        RECT 15.210 157.220 20.250 157.560 ;
        RECT 13.050 156.780 14.770 157.120 ;
        RECT 16.660 156.930 17.000 157.220 ;
        RECT 21.700 157.120 22.040 157.660 ;
        RECT 21.330 156.780 22.410 157.120 ;
        RECT 13.050 155.020 14.130 155.360 ;
        RECT 13.420 154.480 13.760 155.020 ;
        RECT 13.050 154.140 14.130 154.480 ;
        RECT 13.420 153.600 13.760 154.140 ;
        RECT 13.050 153.260 14.130 153.600 ;
        RECT 13.420 152.720 13.760 153.260 ;
        RECT 14.430 153.160 14.770 156.780 ;
        RECT 15.210 156.340 16.290 156.680 ;
        RECT 19.170 156.340 20.250 156.680 ;
        RECT 15.210 155.460 16.290 155.800 ;
        RECT 19.170 155.460 20.250 155.800 ;
        RECT 21.330 155.020 22.410 155.360 ;
        RECT 15.210 154.580 20.250 154.920 ;
        RECT 15.210 153.700 16.290 154.040 ;
        RECT 16.590 153.160 16.930 154.580 ;
        RECT 21.700 154.480 22.040 155.020 ;
        RECT 21.330 154.140 22.410 154.480 ;
        RECT 19.170 153.700 20.250 154.040 ;
        RECT 21.700 153.600 22.040 154.140 ;
        RECT 21.330 153.260 22.410 153.600 ;
        RECT 14.430 152.820 20.250 153.160 ;
        RECT 21.700 152.720 22.040 153.260 ;
        RECT 13.050 152.380 14.130 152.720 ;
        RECT 20.690 152.380 22.410 152.720 ;
        RECT 15.210 151.940 16.290 152.280 ;
        RECT 19.170 151.940 20.250 152.280 ;
        RECT 20.690 151.400 21.030 152.380 ;
        RECT 15.210 151.060 21.030 151.400 ;
        RECT 13.050 150.620 14.130 150.960 ;
        RECT 21.330 150.620 23.050 150.960 ;
        RECT 15.210 150.180 16.290 150.520 ;
        RECT 19.170 150.180 20.250 150.520 ;
        RECT 21.700 150.080 22.040 150.620 ;
        RECT 13.050 149.740 14.770 150.080 ;
        RECT 21.330 149.740 22.410 150.080 ;
        RECT 12.410 148.860 14.130 149.200 ;
        RECT 12.410 138.640 12.750 148.860 ;
        RECT 13.050 147.100 14.130 147.440 ;
        RECT 14.430 146.560 14.770 149.740 ;
        RECT 15.210 149.300 16.290 149.640 ;
        RECT 19.170 149.300 20.250 149.640 ;
        RECT 21.700 149.200 22.040 149.740 ;
        RECT 21.330 148.860 22.410 149.200 ;
        RECT 15.210 148.420 16.290 148.760 ;
        RECT 19.170 148.420 20.250 148.760 ;
        RECT 15.210 147.540 20.250 147.880 ;
        RECT 22.710 147.440 23.050 150.620 ;
        RECT 21.330 147.100 23.050 147.440 ;
        RECT 15.210 146.660 16.290 147.000 ;
        RECT 19.170 146.660 20.250 147.000 ;
        RECT 21.700 146.560 22.040 147.100 ;
        RECT 13.050 146.220 14.770 146.560 ;
        RECT 21.330 146.220 22.410 146.560 ;
        RECT 13.050 145.340 14.130 145.680 ;
        RECT 14.430 144.360 14.770 146.220 ;
        RECT 15.210 145.780 16.290 146.120 ;
        RECT 19.170 145.780 20.250 146.120 ;
        RECT 21.700 145.680 22.040 146.220 ;
        RECT 21.330 145.340 22.410 145.680 ;
        RECT 15.210 144.900 16.290 145.240 ;
        RECT 19.170 144.900 20.250 145.240 ;
        RECT 14.430 144.020 20.250 144.360 ;
        RECT 13.050 143.580 14.130 143.920 ;
        RECT 21.330 143.580 22.410 143.920 ;
        RECT 13.830 143.240 14.770 143.580 ;
        RECT 14.430 142.600 14.770 143.240 ;
        RECT 15.210 143.140 16.290 143.480 ;
        RECT 19.170 143.140 20.250 143.480 ;
        RECT 14.430 142.260 18.870 142.600 ;
        RECT 19.170 142.260 20.250 142.600 ;
        RECT 13.050 141.820 14.130 142.160 ;
        RECT 15.210 141.380 16.290 141.720 ;
        RECT 15.210 140.500 16.290 140.840 ;
        RECT 13.050 140.060 14.130 140.400 ;
        RECT 15.210 139.620 16.930 139.960 ;
        RECT 16.590 139.080 16.930 139.620 ;
        RECT 15.210 138.740 16.930 139.080 ;
        RECT 12.410 138.300 14.130 138.640 ;
        RECT 15.210 137.860 16.290 138.200 ;
        RECT 16.590 137.320 16.930 138.740 ;
        RECT 18.530 138.200 18.870 142.260 ;
        RECT 20.550 141.820 22.410 142.160 ;
        RECT 19.170 141.380 20.250 141.720 ;
        RECT 19.540 140.840 19.880 141.380 ;
        RECT 19.170 140.500 20.250 140.840 ;
        RECT 19.170 139.620 20.250 139.960 ;
        RECT 19.540 139.080 19.880 139.620 ;
        RECT 19.170 138.740 20.250 139.080 ;
        RECT 18.530 137.860 20.250 138.200 ;
        RECT 15.210 136.980 16.930 137.320 ;
        RECT 19.170 136.980 20.250 137.320 ;
        RECT 13.050 136.540 14.130 136.880 ;
        RECT 20.550 136.440 20.890 141.820 ;
        RECT 21.330 140.060 22.410 140.400 ;
        RECT 21.330 138.300 22.410 138.640 ;
        RECT 22.710 136.880 23.050 147.100 ;
        RECT 21.330 136.540 23.050 136.880 ;
        RECT 15.210 136.100 20.890 136.440 ;
        RECT 14.430 135.220 16.290 135.560 ;
        RECT 19.170 135.220 20.890 135.560 ;
        RECT 14.430 135.120 14.770 135.220 ;
        RECT 10.890 134.780 14.770 135.120 ;
        RECT 10.890 133.850 11.970 134.780 ;
        RECT 14.430 134.680 14.770 134.780 ;
        RECT 20.550 135.120 20.890 135.220 ;
        RECT 23.490 135.120 24.570 186.700 ;
        RECT 27.170 186.600 27.510 186.700 ;
        RECT 33.290 187.040 33.630 187.140 ;
        RECT 36.090 187.040 37.170 187.970 ;
        RECT 39.630 187.140 41.490 187.480 ;
        RECT 44.370 187.140 46.090 187.480 ;
        RECT 39.630 187.040 39.970 187.140 ;
        RECT 33.290 186.700 39.970 187.040 ;
        RECT 33.290 186.600 33.630 186.700 ;
        RECT 27.170 186.260 28.890 186.600 ;
        RECT 31.770 186.260 33.630 186.600 ;
        RECT 27.810 185.380 32.850 185.720 ;
        RECT 25.650 184.940 26.730 185.280 ;
        RECT 33.290 184.940 35.010 185.280 ;
        RECT 27.810 184.500 28.890 184.840 ;
        RECT 31.770 184.500 32.850 184.840 ;
        RECT 27.810 183.620 31.470 183.960 ;
        RECT 31.770 183.620 32.850 183.960 ;
        RECT 25.650 183.180 26.730 183.520 ;
        RECT 31.130 183.080 31.470 183.620 ;
        RECT 33.290 183.080 33.630 184.940 ;
        RECT 33.930 183.180 35.010 183.520 ;
        RECT 27.810 182.740 28.890 183.080 ;
        RECT 31.130 182.740 33.630 183.080 ;
        RECT 25.650 182.300 26.730 182.640 ;
        RECT 33.930 182.300 35.010 182.640 ;
        RECT 27.810 181.860 28.890 182.200 ;
        RECT 31.770 181.860 32.850 182.200 ;
        RECT 33.290 181.960 34.230 182.300 ;
        RECT 33.290 181.320 33.630 181.960 ;
        RECT 27.810 180.980 33.630 181.320 ;
        RECT 25.650 180.540 26.730 180.880 ;
        RECT 33.930 180.540 35.010 180.880 ;
        RECT 27.810 180.100 28.890 180.440 ;
        RECT 31.770 180.100 32.850 180.440 ;
        RECT 33.290 180.200 34.230 180.540 ;
        RECT 33.290 179.560 33.630 180.200 ;
        RECT 27.810 179.220 28.890 179.560 ;
        RECT 31.130 179.220 33.630 179.560 ;
        RECT 25.650 178.780 26.730 179.120 ;
        RECT 31.130 178.680 31.470 179.220 ;
        RECT 33.930 178.780 35.010 179.120 ;
        RECT 27.810 178.340 31.470 178.680 ;
        RECT 31.770 178.340 32.850 178.680 ;
        RECT 25.650 177.900 26.730 178.240 ;
        RECT 33.930 177.900 35.010 178.240 ;
        RECT 27.810 177.460 28.890 177.800 ;
        RECT 31.770 177.460 32.850 177.800 ;
        RECT 27.810 176.580 32.850 176.920 ;
        RECT 34.300 176.480 34.640 177.900 ;
        RECT 25.650 176.140 26.730 176.480 ;
        RECT 33.290 176.140 35.010 176.480 ;
        RECT 27.810 175.700 28.890 176.040 ;
        RECT 31.770 175.700 32.850 176.040 ;
        RECT 33.290 175.160 33.630 176.140 ;
        RECT 27.810 174.820 33.630 175.160 ;
        RECT 25.650 174.380 26.730 174.720 ;
        RECT 33.930 174.380 35.010 174.720 ;
        RECT 27.810 173.940 28.890 174.280 ;
        RECT 31.770 173.940 32.850 174.280 ;
        RECT 27.810 173.060 32.850 173.400 ;
        RECT 25.650 172.620 26.730 172.960 ;
        RECT 26.020 172.080 26.360 172.620 ;
        RECT 27.810 172.180 28.890 172.520 ;
        RECT 25.650 171.740 26.730 172.080 ;
        RECT 27.810 171.300 28.890 171.640 ;
        RECT 25.650 170.860 26.730 171.200 ;
        RECT 26.020 170.320 26.360 170.860 ;
        RECT 27.810 170.420 28.890 170.760 ;
        RECT 25.650 169.980 27.510 170.320 ;
        RECT 25.650 168.220 26.730 168.560 ;
        RECT 26.020 167.680 26.360 168.220 ;
        RECT 25.650 167.340 26.730 167.680 ;
        RECT 26.020 166.800 26.360 167.340 ;
        RECT 25.650 166.460 26.730 166.800 ;
        RECT 26.020 165.920 26.360 166.460 ;
        RECT 27.170 166.360 27.510 169.980 ;
        RECT 31.130 169.880 31.470 173.060 ;
        RECT 33.930 172.620 35.010 172.960 ;
        RECT 31.770 172.180 32.850 172.520 ;
        RECT 34.300 172.080 34.640 172.620 ;
        RECT 33.930 171.740 35.010 172.080 ;
        RECT 31.770 171.300 32.850 171.640 ;
        RECT 34.300 171.200 34.640 171.740 ;
        RECT 33.930 170.860 35.010 171.200 ;
        RECT 31.770 170.420 32.850 170.760 ;
        RECT 34.300 170.320 34.640 170.860 ;
        RECT 33.930 169.980 35.010 170.320 ;
        RECT 27.810 169.540 31.470 169.880 ;
        RECT 31.770 169.540 32.850 169.880 ;
        RECT 27.810 168.660 28.890 169.000 ;
        RECT 31.770 168.660 32.850 169.000 ;
        RECT 33.930 168.220 35.010 168.560 ;
        RECT 27.810 167.780 32.850 168.120 ;
        RECT 27.810 166.900 28.890 167.240 ;
        RECT 29.560 166.360 29.900 166.650 ;
        RECT 31.130 166.360 31.470 167.780 ;
        RECT 34.300 167.680 34.640 168.220 ;
        RECT 33.930 167.340 35.010 167.680 ;
        RECT 31.770 166.900 32.850 167.240 ;
        RECT 34.300 166.800 34.640 167.340 ;
        RECT 33.930 166.460 35.010 166.800 ;
        RECT 27.170 166.020 32.850 166.360 ;
        RECT 25.650 165.580 26.730 165.920 ;
        RECT 29.560 165.730 29.900 166.020 ;
        RECT 34.300 165.920 34.640 166.460 ;
        RECT 33.290 165.580 35.010 165.920 ;
        RECT 27.810 165.140 28.890 165.480 ;
        RECT 31.770 165.140 32.850 165.480 ;
        RECT 27.810 164.260 28.890 164.600 ;
        RECT 31.770 164.260 32.850 164.600 ;
        RECT 25.650 163.820 26.730 164.160 ;
        RECT 26.020 163.280 26.360 163.820 ;
        RECT 27.810 163.380 32.850 163.720 ;
        RECT 25.650 162.940 26.730 163.280 ;
        RECT 26.020 162.400 26.360 162.940 ;
        RECT 27.810 162.500 28.890 162.840 ;
        RECT 25.650 162.060 26.730 162.400 ;
        RECT 26.020 161.520 26.360 162.060 ;
        RECT 30.345 161.960 30.685 162.250 ;
        RECT 31.130 161.960 31.470 163.380 ;
        RECT 31.770 162.500 32.850 162.840 ;
        RECT 33.290 161.960 33.630 165.580 ;
        RECT 33.930 163.820 35.010 164.160 ;
        RECT 34.300 163.280 34.640 163.820 ;
        RECT 33.930 162.940 35.010 163.280 ;
        RECT 34.300 162.400 34.640 162.940 ;
        RECT 33.930 162.060 35.010 162.400 ;
        RECT 27.810 161.620 33.630 161.960 ;
        RECT 25.650 161.180 26.730 161.520 ;
        RECT 30.345 161.330 30.685 161.620 ;
        RECT 34.300 161.520 34.640 162.060 ;
        RECT 33.930 161.180 35.010 161.520 ;
        RECT 27.810 160.740 28.890 161.080 ;
        RECT 31.770 160.740 32.850 161.080 ;
        RECT 27.810 159.860 28.890 160.200 ;
        RECT 31.770 159.860 32.850 160.200 ;
        RECT 25.650 159.420 26.730 159.760 ;
        RECT 33.930 159.420 35.010 159.760 ;
        RECT 26.020 158.880 26.360 159.420 ;
        RECT 27.810 158.980 32.850 159.320 ;
        RECT 25.650 158.540 26.730 158.880 ;
        RECT 26.020 158.000 26.360 158.540 ;
        RECT 27.810 158.100 28.890 158.440 ;
        RECT 25.650 157.660 26.730 158.000 ;
        RECT 31.130 157.850 31.470 158.980 ;
        RECT 34.300 158.880 34.640 159.420 ;
        RECT 33.930 158.540 35.010 158.880 ;
        RECT 31.770 158.100 32.850 158.440 ;
        RECT 34.300 158.000 34.640 158.540 ;
        RECT 26.020 157.120 26.360 157.660 ;
        RECT 31.060 157.560 31.470 157.850 ;
        RECT 33.930 157.660 35.010 158.000 ;
        RECT 27.810 157.220 32.850 157.560 ;
        RECT 25.650 156.780 26.730 157.120 ;
        RECT 31.060 156.930 31.400 157.220 ;
        RECT 34.300 157.120 34.640 157.660 ;
        RECT 33.290 156.780 35.010 157.120 ;
        RECT 27.810 156.340 28.890 156.680 ;
        RECT 31.770 156.340 32.850 156.680 ;
        RECT 27.810 155.460 28.890 155.800 ;
        RECT 31.770 155.460 32.850 155.800 ;
        RECT 25.650 155.020 26.730 155.360 ;
        RECT 26.020 154.480 26.360 155.020 ;
        RECT 27.810 154.580 32.850 154.920 ;
        RECT 25.650 154.140 26.730 154.480 ;
        RECT 26.020 153.600 26.360 154.140 ;
        RECT 27.810 153.700 28.890 154.040 ;
        RECT 25.650 153.260 26.730 153.600 ;
        RECT 26.020 152.720 26.360 153.260 ;
        RECT 31.130 153.160 31.470 154.580 ;
        RECT 31.770 153.700 32.850 154.040 ;
        RECT 33.290 153.160 33.630 156.780 ;
        RECT 33.930 155.020 35.010 155.360 ;
        RECT 34.300 154.480 34.640 155.020 ;
        RECT 33.930 154.140 35.010 154.480 ;
        RECT 34.300 153.600 34.640 154.140 ;
        RECT 33.930 153.260 35.010 153.600 ;
        RECT 27.810 152.820 33.630 153.160 ;
        RECT 34.300 152.720 34.640 153.260 ;
        RECT 25.650 152.380 27.370 152.720 ;
        RECT 33.930 152.380 35.010 152.720 ;
        RECT 27.030 151.400 27.370 152.380 ;
        RECT 27.810 151.940 28.890 152.280 ;
        RECT 31.770 151.940 32.850 152.280 ;
        RECT 27.030 151.060 32.850 151.400 ;
        RECT 25.010 150.620 26.730 150.960 ;
        RECT 33.930 150.620 35.010 150.960 ;
        RECT 25.010 147.440 25.350 150.620 ;
        RECT 26.020 150.080 26.360 150.620 ;
        RECT 27.810 150.180 28.890 150.520 ;
        RECT 31.770 150.180 32.850 150.520 ;
        RECT 25.650 149.740 26.730 150.080 ;
        RECT 33.290 149.740 35.010 150.080 ;
        RECT 26.020 149.200 26.360 149.740 ;
        RECT 27.810 149.300 28.890 149.640 ;
        RECT 31.770 149.300 32.850 149.640 ;
        RECT 25.650 148.860 26.730 149.200 ;
        RECT 27.810 148.420 28.890 148.760 ;
        RECT 31.770 148.420 32.850 148.760 ;
        RECT 27.810 147.540 32.850 147.880 ;
        RECT 25.010 147.100 26.730 147.440 ;
        RECT 25.010 136.880 25.350 147.100 ;
        RECT 26.020 146.560 26.360 147.100 ;
        RECT 27.810 146.660 28.890 147.000 ;
        RECT 31.770 146.660 32.850 147.000 ;
        RECT 33.290 146.560 33.630 149.740 ;
        RECT 33.930 148.860 35.650 149.200 ;
        RECT 33.930 147.100 35.010 147.440 ;
        RECT 25.650 146.220 26.730 146.560 ;
        RECT 33.290 146.220 35.010 146.560 ;
        RECT 26.020 145.680 26.360 146.220 ;
        RECT 27.810 145.780 28.890 146.120 ;
        RECT 31.770 145.780 32.850 146.120 ;
        RECT 25.650 145.340 26.730 145.680 ;
        RECT 27.810 144.900 28.890 145.240 ;
        RECT 31.770 144.900 32.850 145.240 ;
        RECT 33.290 144.360 33.630 146.220 ;
        RECT 33.930 145.340 35.010 145.680 ;
        RECT 27.810 144.020 33.630 144.360 ;
        RECT 25.650 143.580 26.730 143.920 ;
        RECT 33.930 143.580 35.010 143.920 ;
        RECT 27.810 143.140 28.890 143.480 ;
        RECT 31.770 143.140 32.850 143.480 ;
        RECT 33.290 143.240 34.230 143.580 ;
        RECT 33.290 142.600 33.630 143.240 ;
        RECT 27.810 142.260 28.890 142.600 ;
        RECT 29.190 142.260 33.630 142.600 ;
        RECT 25.650 141.820 27.510 142.160 ;
        RECT 25.650 140.060 26.730 140.400 ;
        RECT 25.650 138.300 26.730 138.640 ;
        RECT 25.010 136.540 26.730 136.880 ;
        RECT 27.170 136.440 27.510 141.820 ;
        RECT 27.810 141.380 28.890 141.720 ;
        RECT 28.180 140.840 28.520 141.380 ;
        RECT 27.810 140.500 28.890 140.840 ;
        RECT 27.810 139.620 28.890 139.960 ;
        RECT 28.180 139.080 28.520 139.620 ;
        RECT 27.810 138.740 28.890 139.080 ;
        RECT 29.190 138.200 29.530 142.260 ;
        RECT 33.930 141.820 35.010 142.160 ;
        RECT 31.770 141.380 32.850 141.720 ;
        RECT 31.770 140.500 32.850 140.840 ;
        RECT 33.930 140.060 35.010 140.400 ;
        RECT 27.810 137.860 29.530 138.200 ;
        RECT 31.130 139.620 32.850 139.960 ;
        RECT 31.130 139.080 31.470 139.620 ;
        RECT 31.130 138.740 32.850 139.080 ;
        RECT 31.130 137.320 31.470 138.740 ;
        RECT 35.310 138.640 35.650 148.860 ;
        RECT 33.930 138.300 35.650 138.640 ;
        RECT 31.770 137.860 32.850 138.200 ;
        RECT 27.810 136.980 28.890 137.320 ;
        RECT 31.130 136.980 32.850 137.320 ;
        RECT 33.930 136.540 35.010 136.880 ;
        RECT 27.170 136.100 32.850 136.440 ;
        RECT 27.170 135.220 28.890 135.560 ;
        RECT 31.770 135.220 33.630 135.560 ;
        RECT 27.170 135.120 27.510 135.220 ;
        RECT 20.550 134.780 27.510 135.120 ;
        RECT 20.550 134.680 20.890 134.780 ;
        RECT 14.430 134.340 16.290 134.680 ;
        RECT 19.170 134.340 20.890 134.680 ;
        RECT 23.490 133.850 24.570 134.780 ;
        RECT 27.170 134.680 27.510 134.780 ;
        RECT 33.290 135.120 33.630 135.220 ;
        RECT 36.090 135.120 37.170 186.700 ;
        RECT 39.630 186.600 39.970 186.700 ;
        RECT 45.750 187.040 46.090 187.140 ;
        RECT 48.690 187.040 49.770 187.970 ;
        RECT 52.370 187.140 54.090 187.480 ;
        RECT 56.970 187.140 58.830 187.480 ;
        RECT 52.370 187.040 52.710 187.140 ;
        RECT 45.750 186.700 52.710 187.040 ;
        RECT 45.750 186.600 46.090 186.700 ;
        RECT 39.630 186.260 41.490 186.600 ;
        RECT 44.370 186.260 46.090 186.600 ;
        RECT 44.370 185.720 45.290 185.890 ;
        RECT 40.410 185.380 45.450 185.720 ;
        RECT 38.250 184.940 39.970 185.280 ;
        RECT 46.530 184.940 47.610 185.280 ;
        RECT 38.250 183.180 39.330 183.520 ;
        RECT 39.630 183.080 39.970 184.940 ;
        RECT 40.410 184.500 41.490 184.840 ;
        RECT 44.370 184.500 45.450 184.840 ;
        RECT 40.410 183.620 41.490 183.960 ;
        RECT 41.790 183.620 45.450 183.960 ;
        RECT 41.790 183.080 42.130 183.620 ;
        RECT 46.530 183.180 47.610 183.520 ;
        RECT 39.630 182.740 42.130 183.080 ;
        RECT 44.370 182.740 45.450 183.080 ;
        RECT 38.250 182.300 39.330 182.640 ;
        RECT 46.530 182.300 47.610 182.640 ;
        RECT 39.030 181.960 39.970 182.300 ;
        RECT 39.630 181.320 39.970 181.960 ;
        RECT 40.410 181.860 41.490 182.200 ;
        RECT 44.370 181.860 45.450 182.200 ;
        RECT 39.630 180.980 45.450 181.320 ;
        RECT 38.250 180.540 39.330 180.880 ;
        RECT 46.530 180.540 47.610 180.880 ;
        RECT 39.030 180.200 39.970 180.540 ;
        RECT 39.630 179.560 39.970 180.200 ;
        RECT 40.410 180.100 41.490 180.440 ;
        RECT 44.370 180.100 45.450 180.440 ;
        RECT 39.630 179.220 42.130 179.560 ;
        RECT 44.370 179.220 45.450 179.560 ;
        RECT 38.250 178.780 39.330 179.120 ;
        RECT 41.790 178.680 42.130 179.220 ;
        RECT 46.530 178.780 47.610 179.120 ;
        RECT 40.410 178.340 41.490 178.680 ;
        RECT 41.790 178.340 45.450 178.680 ;
        RECT 38.250 177.900 39.330 178.240 ;
        RECT 46.530 177.900 47.610 178.240 ;
        RECT 38.620 176.480 38.960 177.900 ;
        RECT 40.410 177.460 41.490 177.800 ;
        RECT 44.370 177.460 45.450 177.800 ;
        RECT 40.410 176.580 45.450 176.920 ;
        RECT 38.250 176.140 39.970 176.480 ;
        RECT 46.530 176.140 47.610 176.480 ;
        RECT 39.630 175.160 39.970 176.140 ;
        RECT 40.410 175.700 41.490 176.040 ;
        RECT 44.370 175.700 45.450 176.040 ;
        RECT 39.630 174.820 45.450 175.160 ;
        RECT 38.250 174.380 39.330 174.720 ;
        RECT 46.530 174.380 47.610 174.720 ;
        RECT 40.410 173.940 41.490 174.280 ;
        RECT 44.370 173.940 45.450 174.280 ;
        RECT 40.410 173.060 45.450 173.400 ;
        RECT 38.250 172.620 39.330 172.960 ;
        RECT 38.620 172.080 38.960 172.620 ;
        RECT 40.410 172.180 41.490 172.520 ;
        RECT 38.250 171.740 39.330 172.080 ;
        RECT 38.620 171.200 38.960 171.740 ;
        RECT 40.410 171.300 41.490 171.640 ;
        RECT 38.250 170.860 39.330 171.200 ;
        RECT 38.620 170.320 38.960 170.860 ;
        RECT 40.410 170.420 41.490 170.760 ;
        RECT 38.250 169.980 39.330 170.320 ;
        RECT 41.790 169.880 42.130 173.060 ;
        RECT 46.530 172.620 47.610 172.960 ;
        RECT 44.370 172.180 45.450 172.520 ;
        RECT 46.900 172.080 47.240 172.620 ;
        RECT 46.530 171.740 47.610 172.080 ;
        RECT 44.370 171.300 45.450 171.640 ;
        RECT 46.530 170.860 47.610 171.200 ;
        RECT 44.370 170.420 45.450 170.760 ;
        RECT 46.900 170.320 47.240 170.860 ;
        RECT 45.750 169.980 47.610 170.320 ;
        RECT 40.410 169.540 41.490 169.880 ;
        RECT 41.790 169.540 45.450 169.880 ;
        RECT 40.410 168.660 41.490 169.000 ;
        RECT 44.370 168.660 45.450 169.000 ;
        RECT 38.250 168.220 39.330 168.560 ;
        RECT 38.620 167.680 38.960 168.220 ;
        RECT 40.410 167.780 45.450 168.120 ;
        RECT 38.250 167.340 39.330 167.680 ;
        RECT 38.620 166.800 38.960 167.340 ;
        RECT 40.410 166.900 41.490 167.240 ;
        RECT 38.250 166.460 39.330 166.800 ;
        RECT 38.620 165.920 38.960 166.460 ;
        RECT 41.790 166.360 42.130 167.780 ;
        RECT 44.370 166.900 45.450 167.240 ;
        RECT 43.360 166.360 43.700 166.650 ;
        RECT 45.750 166.360 46.090 169.980 ;
        RECT 46.530 168.220 47.610 168.560 ;
        RECT 46.900 167.680 47.240 168.220 ;
        RECT 46.530 167.340 47.610 167.680 ;
        RECT 46.900 166.800 47.240 167.340 ;
        RECT 46.530 166.460 47.610 166.800 ;
        RECT 40.410 166.020 46.090 166.360 ;
        RECT 38.250 165.580 39.970 165.920 ;
        RECT 43.360 165.730 43.700 166.020 ;
        RECT 46.900 165.920 47.240 166.460 ;
        RECT 46.530 165.580 47.610 165.920 ;
        RECT 38.250 163.820 39.330 164.160 ;
        RECT 38.620 163.280 38.960 163.820 ;
        RECT 38.250 162.940 39.330 163.280 ;
        RECT 38.620 162.400 38.960 162.940 ;
        RECT 38.250 162.060 39.330 162.400 ;
        RECT 38.620 161.520 38.960 162.060 ;
        RECT 39.630 161.960 39.970 165.580 ;
        RECT 40.410 165.140 41.490 165.480 ;
        RECT 44.370 165.140 45.450 165.480 ;
        RECT 40.410 164.260 41.490 164.600 ;
        RECT 44.370 164.260 45.450 164.600 ;
        RECT 46.530 163.820 47.610 164.160 ;
        RECT 40.410 163.380 45.450 163.720 ;
        RECT 40.410 162.500 41.490 162.840 ;
        RECT 41.790 161.960 42.130 163.380 ;
        RECT 46.900 163.280 47.240 163.820 ;
        RECT 46.530 162.940 47.610 163.280 ;
        RECT 44.370 162.500 45.450 162.840 ;
        RECT 46.900 162.400 47.240 162.940 ;
        RECT 42.575 161.960 42.915 162.250 ;
        RECT 46.530 162.060 47.610 162.400 ;
        RECT 39.630 161.620 45.450 161.960 ;
        RECT 38.250 161.180 39.330 161.520 ;
        RECT 42.575 161.330 42.915 161.620 ;
        RECT 46.900 161.520 47.240 162.060 ;
        RECT 46.530 161.180 47.610 161.520 ;
        RECT 40.410 160.740 41.490 161.080 ;
        RECT 44.370 160.740 45.450 161.080 ;
        RECT 40.410 159.860 41.490 160.200 ;
        RECT 44.370 159.860 45.450 160.200 ;
        RECT 38.250 159.420 39.330 159.760 ;
        RECT 46.530 159.420 47.610 159.760 ;
        RECT 38.620 158.880 38.960 159.420 ;
        RECT 40.410 158.980 45.450 159.320 ;
        RECT 38.250 158.540 39.330 158.880 ;
        RECT 38.620 158.000 38.960 158.540 ;
        RECT 40.410 158.100 41.490 158.440 ;
        RECT 38.250 157.660 39.330 158.000 ;
        RECT 41.790 157.850 42.130 158.980 ;
        RECT 46.900 158.880 47.240 159.420 ;
        RECT 46.530 158.540 47.610 158.880 ;
        RECT 44.370 158.100 45.450 158.440 ;
        RECT 46.900 158.000 47.240 158.540 ;
        RECT 38.620 157.120 38.960 157.660 ;
        RECT 41.790 157.560 42.200 157.850 ;
        RECT 46.530 157.660 47.610 158.000 ;
        RECT 40.410 157.220 45.450 157.560 ;
        RECT 38.250 156.780 39.970 157.120 ;
        RECT 41.860 156.930 42.200 157.220 ;
        RECT 46.900 157.120 47.240 157.660 ;
        RECT 46.530 156.780 47.610 157.120 ;
        RECT 38.250 155.020 39.330 155.360 ;
        RECT 38.620 154.480 38.960 155.020 ;
        RECT 38.250 154.140 39.330 154.480 ;
        RECT 38.620 153.600 38.960 154.140 ;
        RECT 38.250 153.260 39.330 153.600 ;
        RECT 38.620 152.720 38.960 153.260 ;
        RECT 39.630 153.160 39.970 156.780 ;
        RECT 40.410 156.340 41.490 156.680 ;
        RECT 44.370 156.340 45.450 156.680 ;
        RECT 40.410 155.460 41.490 155.800 ;
        RECT 44.370 155.460 45.450 155.800 ;
        RECT 46.530 155.020 47.610 155.360 ;
        RECT 40.410 154.580 45.450 154.920 ;
        RECT 40.410 153.700 41.490 154.040 ;
        RECT 41.790 153.160 42.130 154.580 ;
        RECT 46.900 154.480 47.240 155.020 ;
        RECT 46.530 154.140 47.610 154.480 ;
        RECT 44.370 153.700 45.450 154.040 ;
        RECT 46.900 153.600 47.240 154.140 ;
        RECT 46.530 153.260 47.610 153.600 ;
        RECT 39.630 152.820 45.450 153.160 ;
        RECT 46.900 152.720 47.240 153.260 ;
        RECT 38.250 152.380 39.330 152.720 ;
        RECT 45.890 152.380 47.610 152.720 ;
        RECT 40.410 151.940 41.490 152.280 ;
        RECT 44.370 151.940 45.450 152.280 ;
        RECT 45.890 151.400 46.230 152.380 ;
        RECT 40.410 151.060 46.230 151.400 ;
        RECT 38.250 150.620 39.330 150.960 ;
        RECT 46.530 150.620 48.250 150.960 ;
        RECT 40.410 150.180 41.490 150.520 ;
        RECT 44.370 150.180 45.450 150.520 ;
        RECT 46.900 150.080 47.240 150.620 ;
        RECT 38.250 149.740 39.970 150.080 ;
        RECT 46.530 149.740 47.610 150.080 ;
        RECT 37.610 148.860 39.330 149.200 ;
        RECT 37.610 138.640 37.950 148.860 ;
        RECT 38.250 147.100 39.330 147.440 ;
        RECT 39.630 146.560 39.970 149.740 ;
        RECT 40.410 149.300 41.490 149.640 ;
        RECT 44.370 149.300 45.450 149.640 ;
        RECT 46.900 149.200 47.240 149.740 ;
        RECT 46.530 148.860 47.610 149.200 ;
        RECT 40.410 148.420 41.490 148.760 ;
        RECT 44.370 148.420 45.450 148.760 ;
        RECT 40.410 147.540 45.450 147.880 ;
        RECT 47.910 147.440 48.250 150.620 ;
        RECT 46.530 147.100 48.250 147.440 ;
        RECT 40.410 146.660 41.490 147.000 ;
        RECT 44.370 146.660 45.450 147.000 ;
        RECT 46.900 146.560 47.240 147.100 ;
        RECT 38.250 146.220 39.970 146.560 ;
        RECT 46.530 146.220 47.610 146.560 ;
        RECT 38.250 145.340 39.330 145.680 ;
        RECT 39.630 144.360 39.970 146.220 ;
        RECT 40.410 145.780 41.490 146.120 ;
        RECT 44.370 145.780 45.450 146.120 ;
        RECT 46.900 145.680 47.240 146.220 ;
        RECT 46.530 145.340 47.610 145.680 ;
        RECT 40.410 144.900 41.490 145.240 ;
        RECT 44.370 144.900 45.450 145.240 ;
        RECT 39.630 144.020 45.450 144.360 ;
        RECT 38.250 143.580 39.330 143.920 ;
        RECT 46.530 143.580 47.610 143.920 ;
        RECT 39.030 143.240 39.970 143.580 ;
        RECT 39.630 142.600 39.970 143.240 ;
        RECT 40.410 143.140 41.490 143.480 ;
        RECT 44.370 143.140 45.450 143.480 ;
        RECT 39.630 142.260 44.070 142.600 ;
        RECT 44.370 142.260 45.450 142.600 ;
        RECT 38.250 141.820 39.330 142.160 ;
        RECT 40.410 141.380 41.490 141.720 ;
        RECT 40.410 140.500 41.490 140.840 ;
        RECT 38.250 140.060 39.330 140.400 ;
        RECT 40.410 139.620 42.130 139.960 ;
        RECT 41.790 139.080 42.130 139.620 ;
        RECT 40.410 138.740 42.130 139.080 ;
        RECT 37.610 138.300 39.330 138.640 ;
        RECT 40.410 137.860 41.490 138.200 ;
        RECT 41.790 137.320 42.130 138.740 ;
        RECT 43.730 138.200 44.070 142.260 ;
        RECT 45.750 141.820 47.610 142.160 ;
        RECT 44.370 141.380 45.450 141.720 ;
        RECT 44.740 140.840 45.080 141.380 ;
        RECT 44.370 140.500 45.450 140.840 ;
        RECT 44.370 139.620 45.450 139.960 ;
        RECT 44.740 139.080 45.080 139.620 ;
        RECT 44.370 138.740 45.450 139.080 ;
        RECT 43.730 137.860 45.450 138.200 ;
        RECT 40.410 136.980 42.130 137.320 ;
        RECT 44.370 136.980 45.450 137.320 ;
        RECT 38.250 136.540 39.330 136.880 ;
        RECT 45.750 136.440 46.090 141.820 ;
        RECT 46.530 140.060 47.610 140.400 ;
        RECT 46.530 138.300 47.610 138.640 ;
        RECT 47.910 136.880 48.250 147.100 ;
        RECT 46.530 136.540 48.250 136.880 ;
        RECT 40.410 136.100 46.090 136.440 ;
        RECT 39.630 135.220 41.490 135.560 ;
        RECT 44.370 135.220 46.090 135.560 ;
        RECT 39.630 135.120 39.970 135.220 ;
        RECT 33.290 134.780 39.970 135.120 ;
        RECT 33.290 134.680 33.630 134.780 ;
        RECT 27.170 134.340 28.890 134.680 ;
        RECT 31.770 134.340 33.630 134.680 ;
        RECT 36.090 133.850 37.170 134.780 ;
        RECT 39.630 134.680 39.970 134.780 ;
        RECT 45.750 135.120 46.090 135.220 ;
        RECT 48.690 135.120 49.770 186.700 ;
        RECT 52.370 186.600 52.710 186.700 ;
        RECT 58.490 187.040 58.830 187.140 ;
        RECT 61.290 187.040 62.370 187.970 ;
        RECT 64.830 187.140 66.690 187.480 ;
        RECT 69.570 187.140 71.290 187.480 ;
        RECT 64.830 187.040 65.170 187.140 ;
        RECT 58.490 186.700 65.170 187.040 ;
        RECT 58.490 186.600 58.830 186.700 ;
        RECT 52.370 186.260 54.090 186.600 ;
        RECT 56.970 186.260 58.830 186.600 ;
        RECT 53.010 185.380 58.050 185.720 ;
        RECT 50.850 184.940 51.930 185.280 ;
        RECT 58.490 184.940 60.210 185.280 ;
        RECT 53.010 184.500 54.090 184.840 ;
        RECT 56.970 184.500 58.050 184.840 ;
        RECT 53.010 183.620 56.670 183.960 ;
        RECT 56.970 183.620 58.050 183.960 ;
        RECT 50.850 183.180 51.930 183.520 ;
        RECT 56.330 183.080 56.670 183.620 ;
        RECT 58.490 183.080 58.830 184.940 ;
        RECT 59.130 183.180 60.210 183.520 ;
        RECT 53.010 182.740 54.090 183.080 ;
        RECT 56.330 182.740 58.830 183.080 ;
        RECT 50.850 182.300 51.930 182.640 ;
        RECT 59.130 182.300 60.210 182.640 ;
        RECT 53.010 181.860 54.090 182.200 ;
        RECT 56.970 181.860 58.050 182.200 ;
        RECT 58.490 181.960 59.430 182.300 ;
        RECT 58.490 181.320 58.830 181.960 ;
        RECT 53.010 180.980 58.830 181.320 ;
        RECT 50.850 180.540 51.930 180.880 ;
        RECT 59.130 180.540 60.210 180.880 ;
        RECT 53.010 180.100 54.090 180.440 ;
        RECT 56.970 180.100 58.050 180.440 ;
        RECT 58.490 180.200 59.430 180.540 ;
        RECT 58.490 179.560 58.830 180.200 ;
        RECT 53.010 179.220 54.090 179.560 ;
        RECT 56.330 179.220 58.830 179.560 ;
        RECT 50.850 178.780 51.930 179.120 ;
        RECT 56.330 178.680 56.670 179.220 ;
        RECT 59.130 178.780 60.210 179.120 ;
        RECT 53.010 178.340 56.670 178.680 ;
        RECT 56.970 178.340 58.050 178.680 ;
        RECT 50.850 177.900 51.930 178.240 ;
        RECT 59.130 177.900 60.210 178.240 ;
        RECT 53.010 177.460 54.090 177.800 ;
        RECT 56.970 177.460 58.050 177.800 ;
        RECT 53.010 176.580 58.050 176.920 ;
        RECT 59.500 176.480 59.840 177.900 ;
        RECT 50.850 176.140 51.930 176.480 ;
        RECT 58.490 176.140 60.210 176.480 ;
        RECT 53.010 175.700 54.090 176.040 ;
        RECT 56.970 175.700 58.050 176.040 ;
        RECT 58.490 175.160 58.830 176.140 ;
        RECT 53.010 174.820 58.830 175.160 ;
        RECT 50.850 174.380 51.930 174.720 ;
        RECT 59.130 174.380 60.210 174.720 ;
        RECT 53.010 173.940 54.090 174.280 ;
        RECT 56.970 173.940 58.050 174.280 ;
        RECT 53.010 173.060 58.050 173.400 ;
        RECT 50.850 172.620 51.930 172.960 ;
        RECT 51.220 172.080 51.560 172.620 ;
        RECT 53.010 172.180 54.090 172.520 ;
        RECT 50.850 171.740 51.930 172.080 ;
        RECT 53.010 171.300 54.090 171.640 ;
        RECT 50.850 170.860 51.930 171.200 ;
        RECT 51.220 170.320 51.560 170.860 ;
        RECT 53.010 170.420 54.090 170.760 ;
        RECT 50.850 169.980 52.710 170.320 ;
        RECT 50.850 168.220 51.930 168.560 ;
        RECT 51.220 167.680 51.560 168.220 ;
        RECT 50.850 167.340 51.930 167.680 ;
        RECT 51.220 166.800 51.560 167.340 ;
        RECT 50.850 166.460 51.930 166.800 ;
        RECT 51.220 165.920 51.560 166.460 ;
        RECT 52.370 166.360 52.710 169.980 ;
        RECT 56.330 169.880 56.670 173.060 ;
        RECT 59.130 172.620 60.210 172.960 ;
        RECT 56.970 172.180 58.050 172.520 ;
        RECT 59.500 172.080 59.840 172.620 ;
        RECT 59.130 171.740 60.210 172.080 ;
        RECT 56.970 171.300 58.050 171.640 ;
        RECT 59.500 171.200 59.840 171.740 ;
        RECT 59.130 170.860 60.210 171.200 ;
        RECT 56.970 170.420 58.050 170.760 ;
        RECT 59.500 170.320 59.840 170.860 ;
        RECT 59.130 169.980 60.210 170.320 ;
        RECT 53.010 169.540 56.670 169.880 ;
        RECT 56.970 169.540 58.050 169.880 ;
        RECT 53.010 168.660 54.090 169.000 ;
        RECT 56.970 168.660 58.050 169.000 ;
        RECT 59.130 168.220 60.210 168.560 ;
        RECT 53.010 167.780 58.050 168.120 ;
        RECT 53.010 166.900 54.090 167.240 ;
        RECT 54.760 166.360 55.100 166.650 ;
        RECT 56.330 166.360 56.670 167.780 ;
        RECT 59.500 167.680 59.840 168.220 ;
        RECT 59.130 167.340 60.210 167.680 ;
        RECT 56.970 166.900 58.050 167.240 ;
        RECT 59.500 166.800 59.840 167.340 ;
        RECT 59.130 166.460 60.210 166.800 ;
        RECT 52.370 166.020 58.050 166.360 ;
        RECT 50.850 165.580 51.930 165.920 ;
        RECT 54.760 165.730 55.100 166.020 ;
        RECT 59.500 165.920 59.840 166.460 ;
        RECT 58.490 165.580 60.210 165.920 ;
        RECT 53.010 165.140 54.090 165.480 ;
        RECT 56.970 165.140 58.050 165.480 ;
        RECT 53.010 164.260 54.090 164.600 ;
        RECT 56.970 164.260 58.050 164.600 ;
        RECT 50.850 163.820 51.930 164.160 ;
        RECT 51.220 163.280 51.560 163.820 ;
        RECT 53.010 163.380 58.050 163.720 ;
        RECT 50.850 162.940 51.930 163.280 ;
        RECT 51.220 162.400 51.560 162.940 ;
        RECT 53.010 162.500 54.090 162.840 ;
        RECT 50.850 162.060 51.930 162.400 ;
        RECT 51.220 161.520 51.560 162.060 ;
        RECT 55.545 161.960 55.885 162.250 ;
        RECT 56.330 161.960 56.670 163.380 ;
        RECT 56.970 162.500 58.050 162.840 ;
        RECT 58.490 161.960 58.830 165.580 ;
        RECT 59.130 163.820 60.210 164.160 ;
        RECT 59.500 163.280 59.840 163.820 ;
        RECT 59.130 162.940 60.210 163.280 ;
        RECT 59.500 162.400 59.840 162.940 ;
        RECT 59.130 162.060 60.210 162.400 ;
        RECT 53.010 161.620 58.830 161.960 ;
        RECT 50.850 161.180 51.930 161.520 ;
        RECT 55.545 161.330 55.885 161.620 ;
        RECT 59.500 161.520 59.840 162.060 ;
        RECT 59.130 161.180 60.210 161.520 ;
        RECT 53.010 160.740 54.090 161.080 ;
        RECT 56.970 160.740 58.050 161.080 ;
        RECT 53.010 159.860 54.090 160.200 ;
        RECT 56.970 159.860 58.050 160.200 ;
        RECT 50.850 159.420 51.930 159.760 ;
        RECT 59.130 159.420 60.210 159.760 ;
        RECT 51.220 158.880 51.560 159.420 ;
        RECT 53.010 158.980 58.050 159.320 ;
        RECT 50.850 158.540 51.930 158.880 ;
        RECT 51.220 158.000 51.560 158.540 ;
        RECT 53.010 158.100 54.090 158.440 ;
        RECT 50.850 157.660 51.930 158.000 ;
        RECT 56.330 157.850 56.670 158.980 ;
        RECT 59.500 158.880 59.840 159.420 ;
        RECT 59.130 158.540 60.210 158.880 ;
        RECT 56.970 158.100 58.050 158.440 ;
        RECT 59.500 158.000 59.840 158.540 ;
        RECT 51.220 157.120 51.560 157.660 ;
        RECT 56.260 157.560 56.670 157.850 ;
        RECT 59.130 157.660 60.210 158.000 ;
        RECT 53.010 157.220 58.050 157.560 ;
        RECT 50.850 156.780 51.930 157.120 ;
        RECT 56.260 156.930 56.600 157.220 ;
        RECT 59.500 157.120 59.840 157.660 ;
        RECT 58.490 156.780 60.210 157.120 ;
        RECT 53.010 156.340 54.090 156.680 ;
        RECT 56.970 156.340 58.050 156.680 ;
        RECT 53.010 155.460 54.090 155.800 ;
        RECT 56.970 155.460 58.050 155.800 ;
        RECT 50.850 155.020 51.930 155.360 ;
        RECT 51.220 154.480 51.560 155.020 ;
        RECT 53.010 154.580 58.050 154.920 ;
        RECT 50.850 154.140 51.930 154.480 ;
        RECT 51.220 153.600 51.560 154.140 ;
        RECT 53.010 153.700 54.090 154.040 ;
        RECT 50.850 153.260 51.930 153.600 ;
        RECT 51.220 152.720 51.560 153.260 ;
        RECT 56.330 153.160 56.670 154.580 ;
        RECT 56.970 153.700 58.050 154.040 ;
        RECT 58.490 153.160 58.830 156.780 ;
        RECT 59.130 155.020 60.210 155.360 ;
        RECT 59.500 154.480 59.840 155.020 ;
        RECT 59.130 154.140 60.210 154.480 ;
        RECT 59.500 153.600 59.840 154.140 ;
        RECT 59.130 153.260 60.210 153.600 ;
        RECT 53.010 152.820 58.830 153.160 ;
        RECT 59.500 152.720 59.840 153.260 ;
        RECT 50.850 152.380 52.570 152.720 ;
        RECT 59.130 152.380 60.210 152.720 ;
        RECT 52.230 151.400 52.570 152.380 ;
        RECT 53.010 151.940 54.090 152.280 ;
        RECT 56.970 151.940 58.050 152.280 ;
        RECT 52.230 151.060 58.050 151.400 ;
        RECT 50.210 150.620 51.930 150.960 ;
        RECT 59.130 150.620 60.210 150.960 ;
        RECT 50.210 147.440 50.550 150.620 ;
        RECT 51.220 150.080 51.560 150.620 ;
        RECT 53.010 150.180 54.090 150.520 ;
        RECT 56.970 150.180 58.050 150.520 ;
        RECT 50.850 149.740 51.930 150.080 ;
        RECT 58.490 149.740 60.210 150.080 ;
        RECT 51.220 149.200 51.560 149.740 ;
        RECT 53.010 149.300 54.090 149.640 ;
        RECT 56.970 149.300 58.050 149.640 ;
        RECT 50.850 148.860 51.930 149.200 ;
        RECT 53.010 148.420 54.090 148.760 ;
        RECT 56.970 148.420 58.050 148.760 ;
        RECT 53.010 147.540 58.050 147.880 ;
        RECT 50.210 147.100 51.930 147.440 ;
        RECT 50.210 136.880 50.550 147.100 ;
        RECT 51.220 146.560 51.560 147.100 ;
        RECT 53.010 146.660 54.090 147.000 ;
        RECT 56.970 146.660 58.050 147.000 ;
        RECT 58.490 146.560 58.830 149.740 ;
        RECT 59.130 148.860 60.850 149.200 ;
        RECT 59.130 147.100 60.210 147.440 ;
        RECT 50.850 146.220 51.930 146.560 ;
        RECT 58.490 146.220 60.210 146.560 ;
        RECT 51.220 145.680 51.560 146.220 ;
        RECT 53.010 145.780 54.090 146.120 ;
        RECT 56.970 145.780 58.050 146.120 ;
        RECT 50.850 145.340 51.930 145.680 ;
        RECT 53.010 144.900 54.090 145.240 ;
        RECT 56.970 144.900 58.050 145.240 ;
        RECT 58.490 144.360 58.830 146.220 ;
        RECT 59.130 145.340 60.210 145.680 ;
        RECT 53.010 144.020 58.830 144.360 ;
        RECT 50.850 143.580 51.930 143.920 ;
        RECT 59.130 143.580 60.210 143.920 ;
        RECT 53.010 143.140 54.090 143.480 ;
        RECT 56.970 143.140 58.050 143.480 ;
        RECT 58.490 143.240 59.430 143.580 ;
        RECT 58.490 142.600 58.830 143.240 ;
        RECT 53.010 142.260 54.090 142.600 ;
        RECT 54.390 142.260 58.830 142.600 ;
        RECT 50.850 141.820 52.710 142.160 ;
        RECT 50.850 140.060 51.930 140.400 ;
        RECT 50.850 138.300 51.930 138.640 ;
        RECT 50.210 136.540 51.930 136.880 ;
        RECT 52.370 136.440 52.710 141.820 ;
        RECT 53.010 141.380 54.090 141.720 ;
        RECT 53.380 140.840 53.720 141.380 ;
        RECT 53.010 140.500 54.090 140.840 ;
        RECT 53.010 139.620 54.090 139.960 ;
        RECT 53.380 139.080 53.720 139.620 ;
        RECT 53.010 138.740 54.090 139.080 ;
        RECT 54.390 138.200 54.730 142.260 ;
        RECT 59.130 141.820 60.210 142.160 ;
        RECT 56.970 141.380 58.050 141.720 ;
        RECT 56.970 140.500 58.050 140.840 ;
        RECT 59.130 140.060 60.210 140.400 ;
        RECT 53.010 137.860 54.730 138.200 ;
        RECT 56.330 139.620 58.050 139.960 ;
        RECT 56.330 139.080 56.670 139.620 ;
        RECT 56.330 138.740 58.050 139.080 ;
        RECT 56.330 137.320 56.670 138.740 ;
        RECT 60.510 138.640 60.850 148.860 ;
        RECT 59.130 138.300 60.850 138.640 ;
        RECT 56.970 137.860 58.050 138.200 ;
        RECT 53.010 136.980 54.090 137.320 ;
        RECT 56.330 136.980 58.050 137.320 ;
        RECT 59.130 136.540 60.210 136.880 ;
        RECT 52.370 136.100 58.050 136.440 ;
        RECT 52.370 135.220 54.090 135.560 ;
        RECT 56.970 135.220 58.830 135.560 ;
        RECT 52.370 135.120 52.710 135.220 ;
        RECT 45.750 134.780 52.710 135.120 ;
        RECT 45.750 134.680 46.090 134.780 ;
        RECT 39.630 134.340 41.490 134.680 ;
        RECT 44.370 134.340 46.090 134.680 ;
        RECT 48.690 133.850 49.770 134.780 ;
        RECT 52.370 134.680 52.710 134.780 ;
        RECT 58.490 135.120 58.830 135.220 ;
        RECT 61.290 135.120 62.370 186.700 ;
        RECT 64.830 186.600 65.170 186.700 ;
        RECT 70.950 187.040 71.290 187.140 ;
        RECT 73.890 187.040 74.970 187.970 ;
        RECT 77.570 187.140 79.290 187.480 ;
        RECT 82.170 187.140 84.030 187.480 ;
        RECT 77.570 187.040 77.910 187.140 ;
        RECT 70.950 186.700 77.910 187.040 ;
        RECT 70.950 186.600 71.290 186.700 ;
        RECT 64.830 186.260 66.690 186.600 ;
        RECT 69.570 186.260 71.290 186.600 ;
        RECT 69.570 185.720 70.490 185.890 ;
        RECT 65.610 185.380 70.650 185.720 ;
        RECT 63.450 184.940 65.170 185.280 ;
        RECT 71.730 184.940 72.810 185.280 ;
        RECT 63.450 183.180 64.530 183.520 ;
        RECT 64.830 183.080 65.170 184.940 ;
        RECT 65.610 184.500 66.690 184.840 ;
        RECT 69.570 184.500 70.650 184.840 ;
        RECT 65.610 183.620 66.690 183.960 ;
        RECT 66.990 183.620 70.650 183.960 ;
        RECT 66.990 183.080 67.330 183.620 ;
        RECT 71.730 183.180 72.810 183.520 ;
        RECT 64.830 182.740 67.330 183.080 ;
        RECT 69.570 182.740 70.650 183.080 ;
        RECT 63.450 182.300 64.530 182.640 ;
        RECT 71.730 182.300 72.810 182.640 ;
        RECT 64.230 181.960 65.170 182.300 ;
        RECT 64.830 181.320 65.170 181.960 ;
        RECT 65.610 181.860 66.690 182.200 ;
        RECT 69.570 181.860 70.650 182.200 ;
        RECT 64.830 180.980 70.650 181.320 ;
        RECT 63.450 180.540 64.530 180.880 ;
        RECT 71.730 180.540 72.810 180.880 ;
        RECT 64.230 180.200 65.170 180.540 ;
        RECT 64.830 179.560 65.170 180.200 ;
        RECT 65.610 180.100 66.690 180.440 ;
        RECT 69.570 180.100 70.650 180.440 ;
        RECT 64.830 179.220 67.330 179.560 ;
        RECT 69.570 179.220 70.650 179.560 ;
        RECT 63.450 178.780 64.530 179.120 ;
        RECT 66.990 178.680 67.330 179.220 ;
        RECT 71.730 178.780 72.810 179.120 ;
        RECT 65.610 178.340 66.690 178.680 ;
        RECT 66.990 178.340 70.650 178.680 ;
        RECT 63.450 177.900 64.530 178.240 ;
        RECT 71.730 177.900 72.810 178.240 ;
        RECT 63.820 176.480 64.160 177.900 ;
        RECT 65.610 177.460 66.690 177.800 ;
        RECT 69.570 177.460 70.650 177.800 ;
        RECT 65.610 176.580 70.650 176.920 ;
        RECT 63.450 176.140 65.170 176.480 ;
        RECT 71.730 176.140 72.810 176.480 ;
        RECT 64.830 175.160 65.170 176.140 ;
        RECT 65.610 175.700 66.690 176.040 ;
        RECT 69.570 175.700 70.650 176.040 ;
        RECT 64.830 174.820 70.650 175.160 ;
        RECT 63.450 174.380 64.530 174.720 ;
        RECT 71.730 174.380 72.810 174.720 ;
        RECT 65.610 173.940 66.690 174.280 ;
        RECT 69.570 173.940 70.650 174.280 ;
        RECT 65.610 173.060 70.650 173.400 ;
        RECT 63.450 172.620 64.530 172.960 ;
        RECT 63.820 172.080 64.160 172.620 ;
        RECT 65.610 172.180 66.690 172.520 ;
        RECT 63.450 171.740 64.530 172.080 ;
        RECT 63.820 171.200 64.160 171.740 ;
        RECT 65.610 171.300 66.690 171.640 ;
        RECT 63.450 170.860 64.530 171.200 ;
        RECT 63.820 170.320 64.160 170.860 ;
        RECT 65.610 170.420 66.690 170.760 ;
        RECT 63.450 169.980 64.530 170.320 ;
        RECT 66.990 169.880 67.330 173.060 ;
        RECT 71.730 172.620 72.810 172.960 ;
        RECT 69.570 172.180 70.650 172.520 ;
        RECT 72.100 172.080 72.440 172.620 ;
        RECT 71.730 171.740 72.810 172.080 ;
        RECT 69.570 171.300 70.650 171.640 ;
        RECT 71.730 170.860 72.810 171.200 ;
        RECT 69.570 170.420 70.650 170.760 ;
        RECT 72.100 170.320 72.440 170.860 ;
        RECT 70.950 169.980 72.810 170.320 ;
        RECT 65.610 169.540 66.690 169.880 ;
        RECT 66.990 169.540 70.650 169.880 ;
        RECT 65.610 168.660 66.690 169.000 ;
        RECT 69.570 168.660 70.650 169.000 ;
        RECT 63.450 168.220 64.530 168.560 ;
        RECT 63.820 167.680 64.160 168.220 ;
        RECT 65.610 167.780 70.650 168.120 ;
        RECT 63.450 167.340 64.530 167.680 ;
        RECT 63.820 166.800 64.160 167.340 ;
        RECT 65.610 166.900 66.690 167.240 ;
        RECT 63.450 166.460 64.530 166.800 ;
        RECT 63.820 165.920 64.160 166.460 ;
        RECT 66.990 166.360 67.330 167.780 ;
        RECT 69.570 166.900 70.650 167.240 ;
        RECT 68.560 166.360 68.900 166.650 ;
        RECT 70.950 166.360 71.290 169.980 ;
        RECT 71.730 168.220 72.810 168.560 ;
        RECT 72.100 167.680 72.440 168.220 ;
        RECT 71.730 167.340 72.810 167.680 ;
        RECT 72.100 166.800 72.440 167.340 ;
        RECT 71.730 166.460 72.810 166.800 ;
        RECT 65.610 166.020 71.290 166.360 ;
        RECT 63.450 165.580 65.170 165.920 ;
        RECT 68.560 165.730 68.900 166.020 ;
        RECT 72.100 165.920 72.440 166.460 ;
        RECT 71.730 165.580 72.810 165.920 ;
        RECT 63.450 163.820 64.530 164.160 ;
        RECT 63.820 163.280 64.160 163.820 ;
        RECT 63.450 162.940 64.530 163.280 ;
        RECT 63.820 162.400 64.160 162.940 ;
        RECT 63.450 162.060 64.530 162.400 ;
        RECT 63.820 161.520 64.160 162.060 ;
        RECT 64.830 161.960 65.170 165.580 ;
        RECT 65.610 165.140 66.690 165.480 ;
        RECT 69.570 165.140 70.650 165.480 ;
        RECT 65.610 164.260 66.690 164.600 ;
        RECT 69.570 164.260 70.650 164.600 ;
        RECT 71.730 163.820 72.810 164.160 ;
        RECT 65.610 163.380 70.650 163.720 ;
        RECT 65.610 162.500 66.690 162.840 ;
        RECT 66.990 161.960 67.330 163.380 ;
        RECT 72.100 163.280 72.440 163.820 ;
        RECT 71.730 162.940 72.810 163.280 ;
        RECT 69.570 162.500 70.650 162.840 ;
        RECT 72.100 162.400 72.440 162.940 ;
        RECT 67.775 161.960 68.115 162.250 ;
        RECT 71.730 162.060 72.810 162.400 ;
        RECT 64.830 161.620 70.650 161.960 ;
        RECT 63.450 161.180 64.530 161.520 ;
        RECT 67.775 161.330 68.115 161.620 ;
        RECT 72.100 161.520 72.440 162.060 ;
        RECT 71.730 161.180 72.810 161.520 ;
        RECT 65.610 160.740 66.690 161.080 ;
        RECT 69.570 160.740 70.650 161.080 ;
        RECT 65.610 159.860 66.690 160.200 ;
        RECT 69.570 159.860 70.650 160.200 ;
        RECT 63.450 159.420 64.530 159.760 ;
        RECT 71.730 159.420 72.810 159.760 ;
        RECT 63.820 158.880 64.160 159.420 ;
        RECT 65.610 158.980 70.650 159.320 ;
        RECT 63.450 158.540 64.530 158.880 ;
        RECT 63.820 158.000 64.160 158.540 ;
        RECT 65.610 158.100 66.690 158.440 ;
        RECT 63.450 157.660 64.530 158.000 ;
        RECT 66.990 157.850 67.330 158.980 ;
        RECT 72.100 158.880 72.440 159.420 ;
        RECT 71.730 158.540 72.810 158.880 ;
        RECT 69.570 158.100 70.650 158.440 ;
        RECT 72.100 158.000 72.440 158.540 ;
        RECT 63.820 157.120 64.160 157.660 ;
        RECT 66.990 157.560 67.400 157.850 ;
        RECT 71.730 157.660 72.810 158.000 ;
        RECT 65.610 157.220 70.650 157.560 ;
        RECT 63.450 156.780 65.170 157.120 ;
        RECT 67.060 156.930 67.400 157.220 ;
        RECT 72.100 157.120 72.440 157.660 ;
        RECT 71.730 156.780 72.810 157.120 ;
        RECT 63.450 155.020 64.530 155.360 ;
        RECT 63.820 154.480 64.160 155.020 ;
        RECT 63.450 154.140 64.530 154.480 ;
        RECT 63.820 153.600 64.160 154.140 ;
        RECT 63.450 153.260 64.530 153.600 ;
        RECT 63.820 152.720 64.160 153.260 ;
        RECT 64.830 153.160 65.170 156.780 ;
        RECT 65.610 156.340 66.690 156.680 ;
        RECT 69.570 156.340 70.650 156.680 ;
        RECT 65.610 155.460 66.690 155.800 ;
        RECT 69.570 155.460 70.650 155.800 ;
        RECT 71.730 155.020 72.810 155.360 ;
        RECT 65.610 154.580 70.650 154.920 ;
        RECT 65.610 153.700 66.690 154.040 ;
        RECT 66.990 153.160 67.330 154.580 ;
        RECT 72.100 154.480 72.440 155.020 ;
        RECT 71.730 154.140 72.810 154.480 ;
        RECT 69.570 153.700 70.650 154.040 ;
        RECT 72.100 153.600 72.440 154.140 ;
        RECT 71.730 153.260 72.810 153.600 ;
        RECT 64.830 152.820 70.650 153.160 ;
        RECT 72.100 152.720 72.440 153.260 ;
        RECT 63.450 152.380 64.530 152.720 ;
        RECT 71.090 152.380 72.810 152.720 ;
        RECT 65.610 151.940 66.690 152.280 ;
        RECT 69.570 151.940 70.650 152.280 ;
        RECT 71.090 151.400 71.430 152.380 ;
        RECT 65.610 151.060 71.430 151.400 ;
        RECT 63.450 150.620 64.530 150.960 ;
        RECT 71.730 150.620 73.450 150.960 ;
        RECT 65.610 150.180 66.690 150.520 ;
        RECT 69.570 150.180 70.650 150.520 ;
        RECT 72.100 150.080 72.440 150.620 ;
        RECT 63.450 149.740 65.170 150.080 ;
        RECT 71.730 149.740 72.810 150.080 ;
        RECT 62.810 148.860 64.530 149.200 ;
        RECT 62.810 138.640 63.150 148.860 ;
        RECT 63.450 147.100 64.530 147.440 ;
        RECT 64.830 146.560 65.170 149.740 ;
        RECT 65.610 149.300 66.690 149.640 ;
        RECT 69.570 149.300 70.650 149.640 ;
        RECT 72.100 149.200 72.440 149.740 ;
        RECT 71.730 148.860 72.810 149.200 ;
        RECT 65.610 148.420 66.690 148.760 ;
        RECT 69.570 148.420 70.650 148.760 ;
        RECT 65.610 147.540 70.650 147.880 ;
        RECT 73.110 147.440 73.450 150.620 ;
        RECT 71.730 147.100 73.450 147.440 ;
        RECT 65.610 146.660 66.690 147.000 ;
        RECT 69.570 146.660 70.650 147.000 ;
        RECT 72.100 146.560 72.440 147.100 ;
        RECT 63.450 146.220 65.170 146.560 ;
        RECT 71.730 146.220 72.810 146.560 ;
        RECT 63.450 145.340 64.530 145.680 ;
        RECT 64.830 144.360 65.170 146.220 ;
        RECT 65.610 145.780 66.690 146.120 ;
        RECT 69.570 145.780 70.650 146.120 ;
        RECT 72.100 145.680 72.440 146.220 ;
        RECT 71.730 145.340 72.810 145.680 ;
        RECT 65.610 144.900 66.690 145.240 ;
        RECT 69.570 144.900 70.650 145.240 ;
        RECT 64.830 144.020 70.650 144.360 ;
        RECT 63.450 143.580 64.530 143.920 ;
        RECT 71.730 143.580 72.810 143.920 ;
        RECT 64.230 143.240 65.170 143.580 ;
        RECT 64.830 142.600 65.170 143.240 ;
        RECT 65.610 143.140 66.690 143.480 ;
        RECT 69.570 143.140 70.650 143.480 ;
        RECT 64.830 142.260 69.270 142.600 ;
        RECT 69.570 142.260 70.650 142.600 ;
        RECT 63.450 141.820 64.530 142.160 ;
        RECT 65.610 141.380 66.690 141.720 ;
        RECT 65.610 140.500 66.690 140.840 ;
        RECT 63.450 140.060 64.530 140.400 ;
        RECT 65.610 139.620 67.330 139.960 ;
        RECT 66.990 139.080 67.330 139.620 ;
        RECT 65.610 138.740 67.330 139.080 ;
        RECT 62.810 138.300 64.530 138.640 ;
        RECT 65.610 137.860 66.690 138.200 ;
        RECT 66.990 137.320 67.330 138.740 ;
        RECT 68.930 138.200 69.270 142.260 ;
        RECT 70.950 141.820 72.810 142.160 ;
        RECT 69.570 141.380 70.650 141.720 ;
        RECT 69.940 140.840 70.280 141.380 ;
        RECT 69.570 140.500 70.650 140.840 ;
        RECT 69.570 139.620 70.650 139.960 ;
        RECT 69.940 139.080 70.280 139.620 ;
        RECT 69.570 138.740 70.650 139.080 ;
        RECT 68.930 137.860 70.650 138.200 ;
        RECT 65.610 136.980 67.330 137.320 ;
        RECT 69.570 136.980 70.650 137.320 ;
        RECT 63.450 136.540 64.530 136.880 ;
        RECT 70.950 136.440 71.290 141.820 ;
        RECT 71.730 140.060 72.810 140.400 ;
        RECT 71.730 138.300 72.810 138.640 ;
        RECT 73.110 136.880 73.450 147.100 ;
        RECT 71.730 136.540 73.450 136.880 ;
        RECT 65.610 136.100 71.290 136.440 ;
        RECT 64.830 135.220 66.690 135.560 ;
        RECT 69.570 135.220 71.290 135.560 ;
        RECT 64.830 135.120 65.170 135.220 ;
        RECT 58.490 134.780 65.170 135.120 ;
        RECT 58.490 134.680 58.830 134.780 ;
        RECT 52.370 134.340 54.090 134.680 ;
        RECT 56.970 134.340 58.830 134.680 ;
        RECT 61.290 133.850 62.370 134.780 ;
        RECT 64.830 134.680 65.170 134.780 ;
        RECT 70.950 135.120 71.290 135.220 ;
        RECT 73.890 135.120 74.970 186.700 ;
        RECT 77.570 186.600 77.910 186.700 ;
        RECT 83.690 187.040 84.030 187.140 ;
        RECT 86.490 187.040 87.570 187.970 ;
        RECT 90.030 187.140 91.890 187.480 ;
        RECT 94.770 187.140 96.490 187.480 ;
        RECT 90.030 187.040 90.370 187.140 ;
        RECT 83.690 186.700 90.370 187.040 ;
        RECT 83.690 186.600 84.030 186.700 ;
        RECT 77.570 186.260 79.290 186.600 ;
        RECT 82.170 186.260 84.030 186.600 ;
        RECT 78.210 185.380 83.250 185.720 ;
        RECT 76.050 184.940 77.130 185.280 ;
        RECT 83.690 184.940 85.410 185.280 ;
        RECT 78.210 184.500 79.290 184.840 ;
        RECT 82.170 184.500 83.250 184.840 ;
        RECT 78.210 183.620 81.870 183.960 ;
        RECT 82.170 183.620 83.250 183.960 ;
        RECT 76.050 183.180 77.130 183.520 ;
        RECT 81.530 183.080 81.870 183.620 ;
        RECT 83.690 183.080 84.030 184.940 ;
        RECT 84.330 183.180 85.410 183.520 ;
        RECT 78.210 182.740 79.290 183.080 ;
        RECT 81.530 182.740 84.030 183.080 ;
        RECT 76.050 182.300 77.130 182.640 ;
        RECT 84.330 182.300 85.410 182.640 ;
        RECT 78.210 181.860 79.290 182.200 ;
        RECT 82.170 181.860 83.250 182.200 ;
        RECT 83.690 181.960 84.630 182.300 ;
        RECT 83.690 181.320 84.030 181.960 ;
        RECT 78.210 180.980 84.030 181.320 ;
        RECT 76.050 180.540 77.130 180.880 ;
        RECT 84.330 180.540 85.410 180.880 ;
        RECT 78.210 180.100 79.290 180.440 ;
        RECT 82.170 180.100 83.250 180.440 ;
        RECT 83.690 180.200 84.630 180.540 ;
        RECT 83.690 179.560 84.030 180.200 ;
        RECT 78.210 179.220 79.290 179.560 ;
        RECT 81.530 179.220 84.030 179.560 ;
        RECT 76.050 178.780 77.130 179.120 ;
        RECT 81.530 178.680 81.870 179.220 ;
        RECT 84.330 178.780 85.410 179.120 ;
        RECT 78.210 178.340 81.870 178.680 ;
        RECT 82.170 178.340 83.250 178.680 ;
        RECT 76.050 177.900 77.130 178.240 ;
        RECT 84.330 177.900 85.410 178.240 ;
        RECT 78.210 177.460 79.290 177.800 ;
        RECT 82.170 177.460 83.250 177.800 ;
        RECT 78.210 176.580 83.250 176.920 ;
        RECT 84.700 176.480 85.040 177.900 ;
        RECT 76.050 176.140 77.130 176.480 ;
        RECT 83.690 176.140 85.410 176.480 ;
        RECT 78.210 175.700 79.290 176.040 ;
        RECT 82.170 175.700 83.250 176.040 ;
        RECT 83.690 175.160 84.030 176.140 ;
        RECT 78.210 174.820 84.030 175.160 ;
        RECT 76.050 174.380 77.130 174.720 ;
        RECT 84.330 174.380 85.410 174.720 ;
        RECT 78.210 173.940 79.290 174.280 ;
        RECT 82.170 173.940 83.250 174.280 ;
        RECT 78.210 173.060 83.250 173.400 ;
        RECT 76.050 172.620 77.130 172.960 ;
        RECT 76.420 172.080 76.760 172.620 ;
        RECT 78.210 172.180 79.290 172.520 ;
        RECT 76.050 171.740 77.130 172.080 ;
        RECT 78.210 171.300 79.290 171.640 ;
        RECT 76.050 170.860 77.130 171.200 ;
        RECT 76.420 170.320 76.760 170.860 ;
        RECT 78.210 170.420 79.290 170.760 ;
        RECT 76.050 169.980 77.910 170.320 ;
        RECT 76.050 168.220 77.130 168.560 ;
        RECT 76.420 167.680 76.760 168.220 ;
        RECT 76.050 167.340 77.130 167.680 ;
        RECT 76.420 166.800 76.760 167.340 ;
        RECT 76.050 166.460 77.130 166.800 ;
        RECT 76.420 165.920 76.760 166.460 ;
        RECT 77.570 166.360 77.910 169.980 ;
        RECT 81.530 169.880 81.870 173.060 ;
        RECT 84.330 172.620 85.410 172.960 ;
        RECT 82.170 172.180 83.250 172.520 ;
        RECT 84.700 172.080 85.040 172.620 ;
        RECT 84.330 171.740 85.410 172.080 ;
        RECT 82.170 171.300 83.250 171.640 ;
        RECT 84.700 171.200 85.040 171.740 ;
        RECT 84.330 170.860 85.410 171.200 ;
        RECT 82.170 170.420 83.250 170.760 ;
        RECT 84.700 170.320 85.040 170.860 ;
        RECT 84.330 169.980 85.410 170.320 ;
        RECT 78.210 169.540 81.870 169.880 ;
        RECT 82.170 169.540 83.250 169.880 ;
        RECT 78.210 168.660 79.290 169.000 ;
        RECT 82.170 168.660 83.250 169.000 ;
        RECT 84.330 168.220 85.410 168.560 ;
        RECT 78.210 167.780 83.250 168.120 ;
        RECT 78.210 166.900 79.290 167.240 ;
        RECT 79.960 166.360 80.300 166.650 ;
        RECT 81.530 166.360 81.870 167.780 ;
        RECT 84.700 167.680 85.040 168.220 ;
        RECT 84.330 167.340 85.410 167.680 ;
        RECT 82.170 166.900 83.250 167.240 ;
        RECT 84.700 166.800 85.040 167.340 ;
        RECT 84.330 166.460 85.410 166.800 ;
        RECT 77.570 166.020 83.250 166.360 ;
        RECT 76.050 165.580 77.130 165.920 ;
        RECT 79.960 165.730 80.300 166.020 ;
        RECT 84.700 165.920 85.040 166.460 ;
        RECT 83.690 165.580 85.410 165.920 ;
        RECT 78.210 165.140 79.290 165.480 ;
        RECT 82.170 165.140 83.250 165.480 ;
        RECT 78.210 164.260 79.290 164.600 ;
        RECT 82.170 164.260 83.250 164.600 ;
        RECT 76.050 163.820 77.130 164.160 ;
        RECT 76.420 163.280 76.760 163.820 ;
        RECT 78.210 163.380 83.250 163.720 ;
        RECT 76.050 162.940 77.130 163.280 ;
        RECT 76.420 162.400 76.760 162.940 ;
        RECT 78.210 162.500 79.290 162.840 ;
        RECT 76.050 162.060 77.130 162.400 ;
        RECT 76.420 161.520 76.760 162.060 ;
        RECT 80.745 161.960 81.085 162.250 ;
        RECT 81.530 161.960 81.870 163.380 ;
        RECT 82.170 162.500 83.250 162.840 ;
        RECT 83.690 161.960 84.030 165.580 ;
        RECT 84.330 163.820 85.410 164.160 ;
        RECT 84.700 163.280 85.040 163.820 ;
        RECT 84.330 162.940 85.410 163.280 ;
        RECT 84.700 162.400 85.040 162.940 ;
        RECT 84.330 162.060 85.410 162.400 ;
        RECT 78.210 161.620 84.030 161.960 ;
        RECT 76.050 161.180 77.130 161.520 ;
        RECT 80.745 161.330 81.085 161.620 ;
        RECT 84.700 161.520 85.040 162.060 ;
        RECT 84.330 161.180 85.410 161.520 ;
        RECT 78.210 160.740 79.290 161.080 ;
        RECT 82.170 160.740 83.250 161.080 ;
        RECT 78.210 159.860 79.290 160.200 ;
        RECT 82.170 159.860 83.250 160.200 ;
        RECT 76.050 159.420 77.130 159.760 ;
        RECT 84.330 159.420 85.410 159.760 ;
        RECT 76.420 158.880 76.760 159.420 ;
        RECT 78.210 158.980 83.250 159.320 ;
        RECT 76.050 158.540 77.130 158.880 ;
        RECT 76.420 158.000 76.760 158.540 ;
        RECT 78.210 158.100 79.290 158.440 ;
        RECT 76.050 157.660 77.130 158.000 ;
        RECT 81.530 157.850 81.870 158.980 ;
        RECT 84.700 158.880 85.040 159.420 ;
        RECT 84.330 158.540 85.410 158.880 ;
        RECT 82.170 158.100 83.250 158.440 ;
        RECT 84.700 158.000 85.040 158.540 ;
        RECT 76.420 157.120 76.760 157.660 ;
        RECT 81.460 157.560 81.870 157.850 ;
        RECT 84.330 157.660 85.410 158.000 ;
        RECT 78.210 157.220 83.250 157.560 ;
        RECT 76.050 156.780 77.130 157.120 ;
        RECT 81.460 156.930 81.800 157.220 ;
        RECT 84.700 157.120 85.040 157.660 ;
        RECT 83.690 156.780 85.410 157.120 ;
        RECT 78.210 156.340 79.290 156.680 ;
        RECT 82.170 156.340 83.250 156.680 ;
        RECT 78.210 155.460 79.290 155.800 ;
        RECT 82.170 155.460 83.250 155.800 ;
        RECT 76.050 155.020 77.130 155.360 ;
        RECT 76.420 154.480 76.760 155.020 ;
        RECT 78.210 154.580 83.250 154.920 ;
        RECT 76.050 154.140 77.130 154.480 ;
        RECT 76.420 153.600 76.760 154.140 ;
        RECT 78.210 153.700 79.290 154.040 ;
        RECT 76.050 153.260 77.130 153.600 ;
        RECT 76.420 152.720 76.760 153.260 ;
        RECT 81.530 153.160 81.870 154.580 ;
        RECT 82.170 153.700 83.250 154.040 ;
        RECT 83.690 153.160 84.030 156.780 ;
        RECT 84.330 155.020 85.410 155.360 ;
        RECT 84.700 154.480 85.040 155.020 ;
        RECT 84.330 154.140 85.410 154.480 ;
        RECT 84.700 153.600 85.040 154.140 ;
        RECT 84.330 153.260 85.410 153.600 ;
        RECT 78.210 152.820 84.030 153.160 ;
        RECT 84.700 152.720 85.040 153.260 ;
        RECT 76.050 152.380 77.770 152.720 ;
        RECT 84.330 152.380 85.410 152.720 ;
        RECT 77.430 151.400 77.770 152.380 ;
        RECT 78.210 151.940 79.290 152.280 ;
        RECT 82.170 151.940 83.250 152.280 ;
        RECT 77.430 151.060 83.250 151.400 ;
        RECT 75.410 150.620 77.130 150.960 ;
        RECT 84.330 150.620 85.410 150.960 ;
        RECT 75.410 147.440 75.750 150.620 ;
        RECT 76.420 150.080 76.760 150.620 ;
        RECT 78.210 150.180 79.290 150.520 ;
        RECT 82.170 150.180 83.250 150.520 ;
        RECT 76.050 149.740 77.130 150.080 ;
        RECT 83.690 149.740 85.410 150.080 ;
        RECT 76.420 149.200 76.760 149.740 ;
        RECT 78.210 149.300 79.290 149.640 ;
        RECT 82.170 149.300 83.250 149.640 ;
        RECT 76.050 148.860 77.130 149.200 ;
        RECT 78.210 148.420 79.290 148.760 ;
        RECT 82.170 148.420 83.250 148.760 ;
        RECT 78.210 147.540 83.250 147.880 ;
        RECT 75.410 147.100 77.130 147.440 ;
        RECT 75.410 136.880 75.750 147.100 ;
        RECT 76.420 146.560 76.760 147.100 ;
        RECT 78.210 146.660 79.290 147.000 ;
        RECT 82.170 146.660 83.250 147.000 ;
        RECT 83.690 146.560 84.030 149.740 ;
        RECT 84.330 148.860 86.050 149.200 ;
        RECT 84.330 147.100 85.410 147.440 ;
        RECT 76.050 146.220 77.130 146.560 ;
        RECT 83.690 146.220 85.410 146.560 ;
        RECT 76.420 145.680 76.760 146.220 ;
        RECT 78.210 145.780 79.290 146.120 ;
        RECT 82.170 145.780 83.250 146.120 ;
        RECT 76.050 145.340 77.130 145.680 ;
        RECT 78.210 144.900 79.290 145.240 ;
        RECT 82.170 144.900 83.250 145.240 ;
        RECT 83.690 144.360 84.030 146.220 ;
        RECT 84.330 145.340 85.410 145.680 ;
        RECT 78.210 144.020 84.030 144.360 ;
        RECT 76.050 143.580 77.130 143.920 ;
        RECT 84.330 143.580 85.410 143.920 ;
        RECT 78.210 143.140 79.290 143.480 ;
        RECT 82.170 143.140 83.250 143.480 ;
        RECT 83.690 143.240 84.630 143.580 ;
        RECT 83.690 142.600 84.030 143.240 ;
        RECT 78.210 142.260 79.290 142.600 ;
        RECT 79.590 142.260 84.030 142.600 ;
        RECT 76.050 141.820 77.910 142.160 ;
        RECT 76.050 140.060 77.130 140.400 ;
        RECT 76.050 138.300 77.130 138.640 ;
        RECT 75.410 136.540 77.130 136.880 ;
        RECT 77.570 136.440 77.910 141.820 ;
        RECT 78.210 141.380 79.290 141.720 ;
        RECT 78.580 140.840 78.920 141.380 ;
        RECT 78.210 140.500 79.290 140.840 ;
        RECT 78.210 139.620 79.290 139.960 ;
        RECT 78.580 139.080 78.920 139.620 ;
        RECT 78.210 138.740 79.290 139.080 ;
        RECT 79.590 138.200 79.930 142.260 ;
        RECT 84.330 141.820 85.410 142.160 ;
        RECT 82.170 141.380 83.250 141.720 ;
        RECT 82.170 140.500 83.250 140.840 ;
        RECT 84.330 140.060 85.410 140.400 ;
        RECT 78.210 137.860 79.930 138.200 ;
        RECT 81.530 139.620 83.250 139.960 ;
        RECT 81.530 139.080 81.870 139.620 ;
        RECT 81.530 138.740 83.250 139.080 ;
        RECT 81.530 137.320 81.870 138.740 ;
        RECT 85.710 138.640 86.050 148.860 ;
        RECT 84.330 138.300 86.050 138.640 ;
        RECT 82.170 137.860 83.250 138.200 ;
        RECT 78.210 136.980 79.290 137.320 ;
        RECT 81.530 136.980 83.250 137.320 ;
        RECT 84.330 136.540 85.410 136.880 ;
        RECT 77.570 136.100 83.250 136.440 ;
        RECT 77.570 135.220 79.290 135.560 ;
        RECT 82.170 135.220 84.030 135.560 ;
        RECT 77.570 135.120 77.910 135.220 ;
        RECT 70.950 134.780 77.910 135.120 ;
        RECT 70.950 134.680 71.290 134.780 ;
        RECT 64.830 134.340 66.690 134.680 ;
        RECT 69.570 134.340 71.290 134.680 ;
        RECT 73.890 133.850 74.970 134.780 ;
        RECT 77.570 134.680 77.910 134.780 ;
        RECT 83.690 135.120 84.030 135.220 ;
        RECT 86.490 135.120 87.570 186.700 ;
        RECT 90.030 186.600 90.370 186.700 ;
        RECT 96.150 187.040 96.490 187.140 ;
        RECT 99.090 187.040 100.170 187.970 ;
        RECT 102.770 187.140 104.490 187.480 ;
        RECT 107.370 187.140 109.230 187.480 ;
        RECT 102.770 187.040 103.110 187.140 ;
        RECT 96.150 186.700 103.110 187.040 ;
        RECT 96.150 186.600 96.490 186.700 ;
        RECT 90.030 186.260 91.890 186.600 ;
        RECT 94.770 186.260 96.490 186.600 ;
        RECT 94.770 185.720 95.690 185.890 ;
        RECT 90.810 185.380 95.850 185.720 ;
        RECT 88.650 184.940 90.370 185.280 ;
        RECT 96.930 184.940 98.010 185.280 ;
        RECT 88.650 183.180 89.730 183.520 ;
        RECT 90.030 183.080 90.370 184.940 ;
        RECT 90.810 184.500 91.890 184.840 ;
        RECT 94.770 184.500 95.850 184.840 ;
        RECT 90.810 183.620 91.890 183.960 ;
        RECT 92.190 183.620 95.850 183.960 ;
        RECT 92.190 183.080 92.530 183.620 ;
        RECT 96.930 183.180 98.010 183.520 ;
        RECT 90.030 182.740 92.530 183.080 ;
        RECT 94.770 182.740 95.850 183.080 ;
        RECT 88.650 182.300 89.730 182.640 ;
        RECT 96.930 182.300 98.010 182.640 ;
        RECT 89.430 181.960 90.370 182.300 ;
        RECT 90.030 181.320 90.370 181.960 ;
        RECT 90.810 181.860 91.890 182.200 ;
        RECT 94.770 181.860 95.850 182.200 ;
        RECT 90.030 180.980 95.850 181.320 ;
        RECT 88.650 180.540 89.730 180.880 ;
        RECT 96.930 180.540 98.010 180.880 ;
        RECT 89.430 180.200 90.370 180.540 ;
        RECT 90.030 179.560 90.370 180.200 ;
        RECT 90.810 180.100 91.890 180.440 ;
        RECT 94.770 180.100 95.850 180.440 ;
        RECT 90.030 179.220 92.530 179.560 ;
        RECT 94.770 179.220 95.850 179.560 ;
        RECT 88.650 178.780 89.730 179.120 ;
        RECT 92.190 178.680 92.530 179.220 ;
        RECT 96.930 178.780 98.010 179.120 ;
        RECT 90.810 178.340 91.890 178.680 ;
        RECT 92.190 178.340 95.850 178.680 ;
        RECT 88.650 177.900 89.730 178.240 ;
        RECT 96.930 177.900 98.010 178.240 ;
        RECT 89.020 176.480 89.360 177.900 ;
        RECT 90.810 177.460 91.890 177.800 ;
        RECT 94.770 177.460 95.850 177.800 ;
        RECT 90.810 176.580 95.850 176.920 ;
        RECT 88.650 176.140 90.370 176.480 ;
        RECT 96.930 176.140 98.010 176.480 ;
        RECT 90.030 175.160 90.370 176.140 ;
        RECT 90.810 175.700 91.890 176.040 ;
        RECT 94.770 175.700 95.850 176.040 ;
        RECT 90.030 174.820 95.850 175.160 ;
        RECT 88.650 174.380 89.730 174.720 ;
        RECT 96.930 174.380 98.010 174.720 ;
        RECT 90.810 173.940 91.890 174.280 ;
        RECT 94.770 173.940 95.850 174.280 ;
        RECT 90.810 173.060 95.850 173.400 ;
        RECT 88.650 172.620 89.730 172.960 ;
        RECT 89.020 172.080 89.360 172.620 ;
        RECT 90.810 172.180 91.890 172.520 ;
        RECT 88.650 171.740 89.730 172.080 ;
        RECT 89.020 171.200 89.360 171.740 ;
        RECT 90.810 171.300 91.890 171.640 ;
        RECT 88.650 170.860 89.730 171.200 ;
        RECT 89.020 170.320 89.360 170.860 ;
        RECT 90.810 170.420 91.890 170.760 ;
        RECT 88.650 169.980 89.730 170.320 ;
        RECT 92.190 169.880 92.530 173.060 ;
        RECT 96.930 172.620 98.010 172.960 ;
        RECT 94.770 172.180 95.850 172.520 ;
        RECT 97.300 172.080 97.640 172.620 ;
        RECT 96.930 171.740 98.010 172.080 ;
        RECT 94.770 171.300 95.850 171.640 ;
        RECT 96.930 170.860 98.010 171.200 ;
        RECT 94.770 170.420 95.850 170.760 ;
        RECT 97.300 170.320 97.640 170.860 ;
        RECT 96.150 169.980 98.010 170.320 ;
        RECT 90.810 169.540 91.890 169.880 ;
        RECT 92.190 169.540 95.850 169.880 ;
        RECT 90.810 168.660 91.890 169.000 ;
        RECT 94.770 168.660 95.850 169.000 ;
        RECT 88.650 168.220 89.730 168.560 ;
        RECT 89.020 167.680 89.360 168.220 ;
        RECT 90.810 167.780 95.850 168.120 ;
        RECT 88.650 167.340 89.730 167.680 ;
        RECT 89.020 166.800 89.360 167.340 ;
        RECT 90.810 166.900 91.890 167.240 ;
        RECT 88.650 166.460 89.730 166.800 ;
        RECT 89.020 165.920 89.360 166.460 ;
        RECT 92.190 166.360 92.530 167.780 ;
        RECT 94.770 166.900 95.850 167.240 ;
        RECT 93.760 166.360 94.100 166.650 ;
        RECT 96.150 166.360 96.490 169.980 ;
        RECT 96.930 168.220 98.010 168.560 ;
        RECT 97.300 167.680 97.640 168.220 ;
        RECT 96.930 167.340 98.010 167.680 ;
        RECT 97.300 166.800 97.640 167.340 ;
        RECT 96.930 166.460 98.010 166.800 ;
        RECT 90.810 166.020 96.490 166.360 ;
        RECT 88.650 165.580 90.370 165.920 ;
        RECT 93.760 165.730 94.100 166.020 ;
        RECT 97.300 165.920 97.640 166.460 ;
        RECT 96.930 165.580 98.010 165.920 ;
        RECT 88.650 163.820 89.730 164.160 ;
        RECT 89.020 163.280 89.360 163.820 ;
        RECT 88.650 162.940 89.730 163.280 ;
        RECT 89.020 162.400 89.360 162.940 ;
        RECT 88.650 162.060 89.730 162.400 ;
        RECT 89.020 161.520 89.360 162.060 ;
        RECT 90.030 161.960 90.370 165.580 ;
        RECT 90.810 165.140 91.890 165.480 ;
        RECT 94.770 165.140 95.850 165.480 ;
        RECT 90.810 164.260 91.890 164.600 ;
        RECT 94.770 164.260 95.850 164.600 ;
        RECT 96.930 163.820 98.010 164.160 ;
        RECT 90.810 163.380 95.850 163.720 ;
        RECT 90.810 162.500 91.890 162.840 ;
        RECT 92.190 161.960 92.530 163.380 ;
        RECT 97.300 163.280 97.640 163.820 ;
        RECT 96.930 162.940 98.010 163.280 ;
        RECT 94.770 162.500 95.850 162.840 ;
        RECT 97.300 162.400 97.640 162.940 ;
        RECT 92.975 161.960 93.315 162.250 ;
        RECT 96.930 162.060 98.010 162.400 ;
        RECT 90.030 161.620 95.850 161.960 ;
        RECT 88.650 161.180 89.730 161.520 ;
        RECT 92.975 161.330 93.315 161.620 ;
        RECT 97.300 161.520 97.640 162.060 ;
        RECT 96.930 161.180 98.010 161.520 ;
        RECT 90.810 160.740 91.890 161.080 ;
        RECT 94.770 160.740 95.850 161.080 ;
        RECT 90.810 159.860 91.890 160.200 ;
        RECT 94.770 159.860 95.850 160.200 ;
        RECT 88.650 159.420 89.730 159.760 ;
        RECT 96.930 159.420 98.010 159.760 ;
        RECT 89.020 158.880 89.360 159.420 ;
        RECT 90.810 158.980 95.850 159.320 ;
        RECT 88.650 158.540 89.730 158.880 ;
        RECT 89.020 158.000 89.360 158.540 ;
        RECT 90.810 158.100 91.890 158.440 ;
        RECT 88.650 157.660 89.730 158.000 ;
        RECT 92.190 157.850 92.530 158.980 ;
        RECT 97.300 158.880 97.640 159.420 ;
        RECT 96.930 158.540 98.010 158.880 ;
        RECT 94.770 158.100 95.850 158.440 ;
        RECT 97.300 158.000 97.640 158.540 ;
        RECT 89.020 157.120 89.360 157.660 ;
        RECT 92.190 157.560 92.600 157.850 ;
        RECT 96.930 157.660 98.010 158.000 ;
        RECT 90.810 157.220 95.850 157.560 ;
        RECT 88.650 156.780 90.370 157.120 ;
        RECT 92.260 156.930 92.600 157.220 ;
        RECT 97.300 157.120 97.640 157.660 ;
        RECT 96.930 156.780 98.010 157.120 ;
        RECT 88.650 155.020 89.730 155.360 ;
        RECT 89.020 154.480 89.360 155.020 ;
        RECT 88.650 154.140 89.730 154.480 ;
        RECT 89.020 153.600 89.360 154.140 ;
        RECT 88.650 153.260 89.730 153.600 ;
        RECT 89.020 152.720 89.360 153.260 ;
        RECT 90.030 153.160 90.370 156.780 ;
        RECT 90.810 156.340 91.890 156.680 ;
        RECT 94.770 156.340 95.850 156.680 ;
        RECT 90.810 155.460 91.890 155.800 ;
        RECT 94.770 155.460 95.850 155.800 ;
        RECT 96.930 155.020 98.010 155.360 ;
        RECT 90.810 154.580 95.850 154.920 ;
        RECT 90.810 153.700 91.890 154.040 ;
        RECT 92.190 153.160 92.530 154.580 ;
        RECT 97.300 154.480 97.640 155.020 ;
        RECT 96.930 154.140 98.010 154.480 ;
        RECT 94.770 153.700 95.850 154.040 ;
        RECT 97.300 153.600 97.640 154.140 ;
        RECT 96.930 153.260 98.010 153.600 ;
        RECT 90.030 152.820 95.850 153.160 ;
        RECT 97.300 152.720 97.640 153.260 ;
        RECT 88.650 152.380 89.730 152.720 ;
        RECT 96.290 152.380 98.010 152.720 ;
        RECT 90.810 151.940 91.890 152.280 ;
        RECT 94.770 151.940 95.850 152.280 ;
        RECT 96.290 151.400 96.630 152.380 ;
        RECT 90.810 151.060 96.630 151.400 ;
        RECT 88.650 150.620 89.730 150.960 ;
        RECT 96.930 150.620 98.650 150.960 ;
        RECT 90.810 150.180 91.890 150.520 ;
        RECT 94.770 150.180 95.850 150.520 ;
        RECT 97.300 150.080 97.640 150.620 ;
        RECT 88.650 149.740 90.370 150.080 ;
        RECT 96.930 149.740 98.010 150.080 ;
        RECT 88.010 148.860 89.730 149.200 ;
        RECT 88.010 138.640 88.350 148.860 ;
        RECT 88.650 147.100 89.730 147.440 ;
        RECT 90.030 146.560 90.370 149.740 ;
        RECT 90.810 149.300 91.890 149.640 ;
        RECT 94.770 149.300 95.850 149.640 ;
        RECT 97.300 149.200 97.640 149.740 ;
        RECT 96.930 148.860 98.010 149.200 ;
        RECT 90.810 148.420 91.890 148.760 ;
        RECT 94.770 148.420 95.850 148.760 ;
        RECT 90.810 147.540 95.850 147.880 ;
        RECT 98.310 147.440 98.650 150.620 ;
        RECT 96.930 147.100 98.650 147.440 ;
        RECT 90.810 146.660 91.890 147.000 ;
        RECT 94.770 146.660 95.850 147.000 ;
        RECT 97.300 146.560 97.640 147.100 ;
        RECT 88.650 146.220 90.370 146.560 ;
        RECT 96.930 146.220 98.010 146.560 ;
        RECT 88.650 145.340 89.730 145.680 ;
        RECT 90.030 144.360 90.370 146.220 ;
        RECT 90.810 145.780 91.890 146.120 ;
        RECT 94.770 145.780 95.850 146.120 ;
        RECT 97.300 145.680 97.640 146.220 ;
        RECT 96.930 145.340 98.010 145.680 ;
        RECT 90.810 144.900 91.890 145.240 ;
        RECT 94.770 144.900 95.850 145.240 ;
        RECT 90.030 144.020 95.850 144.360 ;
        RECT 88.650 143.580 89.730 143.920 ;
        RECT 96.930 143.580 98.010 143.920 ;
        RECT 89.430 143.240 90.370 143.580 ;
        RECT 90.030 142.600 90.370 143.240 ;
        RECT 90.810 143.140 91.890 143.480 ;
        RECT 94.770 143.140 95.850 143.480 ;
        RECT 90.030 142.260 94.470 142.600 ;
        RECT 94.770 142.260 95.850 142.600 ;
        RECT 88.650 141.820 89.730 142.160 ;
        RECT 90.810 141.380 91.890 141.720 ;
        RECT 90.810 140.500 91.890 140.840 ;
        RECT 88.650 140.060 89.730 140.400 ;
        RECT 90.810 139.620 92.530 139.960 ;
        RECT 92.190 139.080 92.530 139.620 ;
        RECT 90.810 138.740 92.530 139.080 ;
        RECT 88.010 138.300 89.730 138.640 ;
        RECT 90.810 137.860 91.890 138.200 ;
        RECT 92.190 137.320 92.530 138.740 ;
        RECT 94.130 138.200 94.470 142.260 ;
        RECT 96.150 141.820 98.010 142.160 ;
        RECT 94.770 141.380 95.850 141.720 ;
        RECT 95.140 140.840 95.480 141.380 ;
        RECT 94.770 140.500 95.850 140.840 ;
        RECT 94.770 139.620 95.850 139.960 ;
        RECT 95.140 139.080 95.480 139.620 ;
        RECT 94.770 138.740 95.850 139.080 ;
        RECT 94.130 137.860 95.850 138.200 ;
        RECT 90.810 136.980 92.530 137.320 ;
        RECT 94.770 136.980 95.850 137.320 ;
        RECT 88.650 136.540 89.730 136.880 ;
        RECT 96.150 136.440 96.490 141.820 ;
        RECT 96.930 140.060 98.010 140.400 ;
        RECT 96.930 138.300 98.010 138.640 ;
        RECT 98.310 136.880 98.650 147.100 ;
        RECT 96.930 136.540 98.650 136.880 ;
        RECT 90.810 136.100 96.490 136.440 ;
        RECT 90.030 135.220 91.890 135.560 ;
        RECT 94.770 135.220 96.490 135.560 ;
        RECT 90.030 135.120 90.370 135.220 ;
        RECT 83.690 134.780 90.370 135.120 ;
        RECT 83.690 134.680 84.030 134.780 ;
        RECT 77.570 134.340 79.290 134.680 ;
        RECT 82.170 134.340 84.030 134.680 ;
        RECT 86.490 133.850 87.570 134.780 ;
        RECT 90.030 134.680 90.370 134.780 ;
        RECT 96.150 135.120 96.490 135.220 ;
        RECT 99.090 135.120 100.170 186.700 ;
        RECT 102.770 186.600 103.110 186.700 ;
        RECT 108.890 187.040 109.230 187.140 ;
        RECT 111.690 187.040 112.770 187.970 ;
        RECT 108.890 186.700 112.770 187.040 ;
        RECT 108.890 186.600 109.230 186.700 ;
        RECT 102.770 186.260 104.490 186.600 ;
        RECT 107.370 186.260 109.230 186.600 ;
        RECT 103.410 185.380 108.450 185.720 ;
        RECT 101.250 184.940 102.330 185.280 ;
        RECT 108.890 184.940 110.610 185.280 ;
        RECT 103.410 184.500 104.490 184.840 ;
        RECT 107.370 184.500 108.450 184.840 ;
        RECT 103.410 183.620 107.070 183.960 ;
        RECT 107.370 183.620 108.450 183.960 ;
        RECT 101.250 183.180 102.330 183.520 ;
        RECT 106.730 183.080 107.070 183.620 ;
        RECT 108.890 183.080 109.230 184.940 ;
        RECT 109.530 183.180 110.610 183.520 ;
        RECT 103.410 182.740 104.490 183.080 ;
        RECT 106.730 182.740 109.230 183.080 ;
        RECT 111.690 182.640 112.770 186.700 ;
        RECT 115.230 182.740 117.090 183.080 ;
        RECT 119.970 182.740 121.690 183.080 ;
        RECT 115.230 182.640 115.570 182.740 ;
        RECT 101.250 182.300 102.330 182.640 ;
        RECT 109.530 182.300 110.610 182.640 ;
        RECT 111.690 182.300 115.570 182.640 ;
        RECT 103.410 181.860 104.490 182.200 ;
        RECT 107.370 181.860 108.450 182.200 ;
        RECT 108.890 181.960 109.830 182.300 ;
        RECT 108.890 181.320 109.230 181.960 ;
        RECT 103.410 180.980 109.230 181.320 ;
        RECT 101.250 180.540 102.330 180.880 ;
        RECT 109.530 180.540 110.610 180.880 ;
        RECT 103.410 180.100 104.490 180.440 ;
        RECT 107.370 180.100 108.450 180.440 ;
        RECT 108.890 180.200 109.830 180.540 ;
        RECT 108.890 179.560 109.230 180.200 ;
        RECT 103.410 179.220 104.490 179.560 ;
        RECT 106.730 179.220 109.230 179.560 ;
        RECT 101.250 178.780 102.330 179.120 ;
        RECT 106.730 178.680 107.070 179.220 ;
        RECT 109.530 178.780 110.610 179.120 ;
        RECT 103.410 178.340 107.070 178.680 ;
        RECT 107.370 178.340 108.450 178.680 ;
        RECT 101.250 177.900 102.330 178.240 ;
        RECT 109.530 177.900 110.610 178.240 ;
        RECT 103.410 177.460 104.490 177.800 ;
        RECT 107.370 177.460 108.450 177.800 ;
        RECT 103.410 176.580 108.450 176.920 ;
        RECT 109.900 176.480 110.240 177.900 ;
        RECT 101.250 176.140 102.330 176.480 ;
        RECT 108.890 176.140 110.610 176.480 ;
        RECT 103.410 175.700 104.490 176.040 ;
        RECT 107.370 175.700 108.450 176.040 ;
        RECT 108.890 175.160 109.230 176.140 ;
        RECT 103.410 174.820 109.230 175.160 ;
        RECT 101.250 174.380 102.330 174.720 ;
        RECT 109.530 174.380 110.610 174.720 ;
        RECT 103.410 173.940 104.490 174.280 ;
        RECT 107.370 173.940 108.450 174.280 ;
        RECT 103.410 173.060 108.450 173.400 ;
        RECT 101.250 172.620 102.330 172.960 ;
        RECT 101.620 172.080 101.960 172.620 ;
        RECT 103.410 172.180 104.490 172.520 ;
        RECT 101.250 171.740 102.330 172.080 ;
        RECT 103.410 171.300 104.490 171.640 ;
        RECT 101.250 170.860 102.330 171.200 ;
        RECT 101.620 170.320 101.960 170.860 ;
        RECT 103.410 170.420 104.490 170.760 ;
        RECT 101.250 169.980 103.110 170.320 ;
        RECT 101.250 168.220 102.330 168.560 ;
        RECT 101.620 167.680 101.960 168.220 ;
        RECT 101.250 167.340 102.330 167.680 ;
        RECT 101.620 166.800 101.960 167.340 ;
        RECT 101.250 166.460 102.330 166.800 ;
        RECT 101.620 165.920 101.960 166.460 ;
        RECT 102.770 166.360 103.110 169.980 ;
        RECT 106.730 169.880 107.070 173.060 ;
        RECT 109.530 172.620 110.610 172.960 ;
        RECT 107.370 172.180 108.450 172.520 ;
        RECT 109.900 172.080 110.240 172.620 ;
        RECT 109.530 171.740 110.610 172.080 ;
        RECT 107.370 171.300 108.450 171.640 ;
        RECT 109.900 171.200 110.240 171.740 ;
        RECT 109.530 170.860 110.610 171.200 ;
        RECT 107.370 170.420 108.450 170.760 ;
        RECT 109.900 170.320 110.240 170.860 ;
        RECT 109.530 169.980 110.610 170.320 ;
        RECT 103.410 169.540 107.070 169.880 ;
        RECT 107.370 169.540 108.450 169.880 ;
        RECT 103.410 168.660 104.490 169.000 ;
        RECT 107.370 168.660 108.450 169.000 ;
        RECT 109.530 168.220 110.610 168.560 ;
        RECT 103.410 167.780 108.450 168.120 ;
        RECT 103.410 166.900 104.490 167.240 ;
        RECT 105.160 166.360 105.500 166.650 ;
        RECT 106.730 166.360 107.070 167.780 ;
        RECT 109.900 167.680 110.240 168.220 ;
        RECT 109.530 167.340 110.610 167.680 ;
        RECT 107.370 166.900 108.450 167.240 ;
        RECT 109.900 166.800 110.240 167.340 ;
        RECT 109.530 166.460 110.610 166.800 ;
        RECT 102.770 166.020 108.450 166.360 ;
        RECT 101.250 165.580 102.330 165.920 ;
        RECT 105.160 165.730 105.500 166.020 ;
        RECT 109.900 165.920 110.240 166.460 ;
        RECT 108.890 165.580 110.610 165.920 ;
        RECT 103.410 165.140 104.490 165.480 ;
        RECT 107.370 165.140 108.450 165.480 ;
        RECT 103.410 164.260 104.490 164.600 ;
        RECT 107.370 164.260 108.450 164.600 ;
        RECT 101.250 163.820 102.330 164.160 ;
        RECT 101.620 163.280 101.960 163.820 ;
        RECT 103.410 163.380 108.450 163.720 ;
        RECT 101.250 162.940 102.330 163.280 ;
        RECT 101.620 162.400 101.960 162.940 ;
        RECT 103.410 162.500 104.490 162.840 ;
        RECT 101.250 162.060 102.330 162.400 ;
        RECT 101.620 161.520 101.960 162.060 ;
        RECT 105.945 161.960 106.285 162.250 ;
        RECT 106.730 161.960 107.070 163.380 ;
        RECT 107.370 162.500 108.450 162.840 ;
        RECT 108.890 161.960 109.230 165.580 ;
        RECT 109.530 163.820 110.610 164.160 ;
        RECT 109.900 163.280 110.240 163.820 ;
        RECT 109.530 162.940 110.610 163.280 ;
        RECT 109.900 162.400 110.240 162.940 ;
        RECT 109.530 162.060 110.610 162.400 ;
        RECT 103.410 161.620 109.230 161.960 ;
        RECT 101.250 161.180 102.330 161.520 ;
        RECT 105.945 161.330 106.285 161.620 ;
        RECT 109.900 161.520 110.240 162.060 ;
        RECT 109.530 161.180 110.610 161.520 ;
        RECT 103.410 160.740 104.490 161.080 ;
        RECT 107.370 160.740 108.450 161.080 ;
        RECT 103.410 159.860 104.490 160.200 ;
        RECT 107.370 159.860 108.450 160.200 ;
        RECT 101.250 159.420 102.330 159.760 ;
        RECT 109.530 159.420 110.610 159.760 ;
        RECT 101.620 158.880 101.960 159.420 ;
        RECT 103.410 158.980 108.450 159.320 ;
        RECT 101.250 158.540 102.330 158.880 ;
        RECT 101.620 158.000 101.960 158.540 ;
        RECT 103.410 158.100 104.490 158.440 ;
        RECT 101.250 157.660 102.330 158.000 ;
        RECT 106.730 157.850 107.070 158.980 ;
        RECT 109.900 158.880 110.240 159.420 ;
        RECT 109.530 158.540 110.610 158.880 ;
        RECT 107.370 158.100 108.450 158.440 ;
        RECT 109.900 158.000 110.240 158.540 ;
        RECT 101.620 157.120 101.960 157.660 ;
        RECT 106.660 157.560 107.070 157.850 ;
        RECT 109.530 157.660 110.610 158.000 ;
        RECT 103.410 157.220 108.450 157.560 ;
        RECT 101.250 156.780 102.330 157.120 ;
        RECT 106.660 156.930 107.000 157.220 ;
        RECT 109.900 157.120 110.240 157.660 ;
        RECT 108.890 156.780 110.610 157.120 ;
        RECT 103.410 156.340 104.490 156.680 ;
        RECT 107.370 156.340 108.450 156.680 ;
        RECT 103.410 155.460 104.490 155.800 ;
        RECT 107.370 155.460 108.450 155.800 ;
        RECT 101.250 155.020 102.330 155.360 ;
        RECT 101.620 154.480 101.960 155.020 ;
        RECT 103.410 154.580 108.450 154.920 ;
        RECT 101.250 154.140 102.330 154.480 ;
        RECT 101.620 153.600 101.960 154.140 ;
        RECT 103.410 153.700 104.490 154.040 ;
        RECT 101.250 153.260 102.330 153.600 ;
        RECT 101.620 152.720 101.960 153.260 ;
        RECT 106.730 153.160 107.070 154.580 ;
        RECT 107.370 153.700 108.450 154.040 ;
        RECT 108.890 153.160 109.230 156.780 ;
        RECT 109.530 155.020 110.610 155.360 ;
        RECT 109.900 154.480 110.240 155.020 ;
        RECT 109.530 154.140 110.610 154.480 ;
        RECT 109.900 153.600 110.240 154.140 ;
        RECT 109.530 153.260 110.610 153.600 ;
        RECT 103.410 152.820 109.230 153.160 ;
        RECT 109.900 152.720 110.240 153.260 ;
        RECT 101.250 152.380 102.970 152.720 ;
        RECT 109.530 152.380 110.610 152.720 ;
        RECT 102.630 151.400 102.970 152.380 ;
        RECT 103.410 151.940 104.490 152.280 ;
        RECT 107.370 151.940 108.450 152.280 ;
        RECT 102.630 151.060 108.450 151.400 ;
        RECT 100.610 150.620 102.330 150.960 ;
        RECT 109.530 150.620 110.610 150.960 ;
        RECT 100.610 147.440 100.950 150.620 ;
        RECT 101.620 150.080 101.960 150.620 ;
        RECT 103.410 150.180 104.490 150.520 ;
        RECT 107.370 150.180 108.450 150.520 ;
        RECT 101.250 149.740 102.330 150.080 ;
        RECT 108.890 149.740 110.610 150.080 ;
        RECT 101.620 149.200 101.960 149.740 ;
        RECT 103.410 149.300 104.490 149.640 ;
        RECT 107.370 149.300 108.450 149.640 ;
        RECT 101.250 148.860 102.330 149.200 ;
        RECT 103.410 148.420 104.490 148.760 ;
        RECT 107.370 148.420 108.450 148.760 ;
        RECT 103.410 147.540 108.450 147.880 ;
        RECT 100.610 147.100 102.330 147.440 ;
        RECT 100.610 136.880 100.950 147.100 ;
        RECT 101.620 146.560 101.960 147.100 ;
        RECT 103.410 146.660 104.490 147.000 ;
        RECT 107.370 146.660 108.450 147.000 ;
        RECT 108.890 146.560 109.230 149.740 ;
        RECT 109.530 148.860 111.250 149.200 ;
        RECT 109.530 147.100 110.610 147.440 ;
        RECT 101.250 146.220 102.330 146.560 ;
        RECT 108.890 146.220 110.610 146.560 ;
        RECT 101.620 145.680 101.960 146.220 ;
        RECT 103.410 145.780 104.490 146.120 ;
        RECT 107.370 145.780 108.450 146.120 ;
        RECT 101.250 145.340 102.330 145.680 ;
        RECT 103.410 144.900 104.490 145.240 ;
        RECT 107.370 144.900 108.450 145.240 ;
        RECT 108.890 144.360 109.230 146.220 ;
        RECT 109.530 145.340 110.610 145.680 ;
        RECT 103.410 144.020 109.230 144.360 ;
        RECT 101.250 143.580 102.330 143.920 ;
        RECT 109.530 143.580 110.610 143.920 ;
        RECT 103.410 143.140 104.490 143.480 ;
        RECT 107.370 143.140 108.450 143.480 ;
        RECT 108.890 143.240 109.830 143.580 ;
        RECT 108.890 142.600 109.230 143.240 ;
        RECT 103.410 142.260 104.490 142.600 ;
        RECT 104.790 142.260 109.230 142.600 ;
        RECT 101.250 141.820 103.110 142.160 ;
        RECT 101.250 140.060 102.330 140.400 ;
        RECT 101.250 138.300 102.330 138.640 ;
        RECT 100.610 136.540 102.330 136.880 ;
        RECT 102.770 136.440 103.110 141.820 ;
        RECT 103.410 141.380 104.490 141.720 ;
        RECT 103.780 140.840 104.120 141.380 ;
        RECT 103.410 140.500 104.490 140.840 ;
        RECT 103.410 139.620 104.490 139.960 ;
        RECT 103.780 139.080 104.120 139.620 ;
        RECT 103.410 138.740 104.490 139.080 ;
        RECT 104.790 138.200 105.130 142.260 ;
        RECT 109.530 141.820 110.610 142.160 ;
        RECT 107.370 141.380 108.450 141.720 ;
        RECT 107.370 140.500 108.450 140.840 ;
        RECT 109.530 140.060 110.610 140.400 ;
        RECT 103.410 137.860 105.130 138.200 ;
        RECT 106.730 139.620 108.450 139.960 ;
        RECT 106.730 139.080 107.070 139.620 ;
        RECT 106.730 138.740 108.450 139.080 ;
        RECT 106.730 137.320 107.070 138.740 ;
        RECT 110.910 138.640 111.250 148.860 ;
        RECT 109.530 138.300 111.250 138.640 ;
        RECT 107.370 137.860 108.450 138.200 ;
        RECT 103.410 136.980 104.490 137.320 ;
        RECT 106.730 136.980 108.450 137.320 ;
        RECT 109.530 136.540 110.610 136.880 ;
        RECT 102.770 136.100 108.450 136.440 ;
        RECT 102.770 135.220 104.490 135.560 ;
        RECT 107.370 135.220 109.230 135.560 ;
        RECT 102.770 135.120 103.110 135.220 ;
        RECT 96.150 134.780 103.110 135.120 ;
        RECT 96.150 134.680 96.490 134.780 ;
        RECT 90.030 134.340 91.890 134.680 ;
        RECT 94.770 134.340 96.490 134.680 ;
        RECT 99.090 133.850 100.170 134.780 ;
        RECT 102.770 134.680 103.110 134.780 ;
        RECT 108.890 135.120 109.230 135.220 ;
        RECT 111.690 135.120 112.770 182.300 ;
        RECT 115.230 182.200 115.570 182.300 ;
        RECT 121.350 182.640 121.690 182.740 ;
        RECT 124.290 182.640 125.370 183.570 ;
        RECT 121.350 182.300 125.370 182.640 ;
        RECT 121.350 182.200 121.690 182.300 ;
        RECT 115.230 181.860 117.090 182.200 ;
        RECT 119.970 181.860 121.690 182.200 ;
        RECT 113.850 180.880 114.770 181.050 ;
        RECT 116.010 180.980 121.690 181.320 ;
        RECT 113.850 180.540 114.930 180.880 ;
        RECT 116.010 180.100 117.090 180.440 ;
        RECT 119.970 180.100 121.050 180.440 ;
        RECT 116.010 179.220 117.090 179.560 ;
        RECT 117.390 179.220 121.050 179.560 ;
        RECT 113.850 178.780 114.930 179.120 ;
        RECT 117.390 178.680 117.730 179.220 ;
        RECT 115.370 178.340 117.730 178.680 ;
        RECT 119.970 178.340 121.050 178.680 ;
        RECT 113.850 177.900 114.930 178.240 ;
        RECT 113.850 176.140 114.930 176.480 ;
        RECT 115.370 175.600 115.710 178.340 ;
        RECT 116.010 177.460 117.090 177.800 ;
        RECT 119.970 177.460 121.050 177.800 ;
        RECT 116.010 176.580 117.730 176.920 ;
        RECT 119.970 176.580 121.050 176.920 ;
        RECT 117.390 176.040 117.730 176.580 ;
        RECT 121.350 176.480 121.690 180.980 ;
        RECT 122.130 180.540 123.210 180.880 ;
        RECT 122.130 178.780 123.210 179.120 ;
        RECT 122.130 177.900 123.210 178.240 ;
        RECT 121.350 176.140 123.210 176.480 ;
        RECT 116.010 175.700 117.090 176.040 ;
        RECT 117.390 175.700 121.050 176.040 ;
        RECT 113.850 175.260 115.710 175.600 ;
        RECT 122.130 175.260 123.210 175.600 ;
        RECT 116.010 174.820 117.090 175.160 ;
        RECT 119.970 174.820 121.050 175.160 ;
        RECT 115.230 173.940 121.050 174.280 ;
        RECT 113.850 173.500 114.930 173.840 ;
        RECT 115.230 172.080 115.570 173.940 ;
        RECT 122.130 173.500 123.210 173.840 ;
        RECT 116.010 173.060 117.090 173.400 ;
        RECT 119.970 173.060 121.050 173.400 ;
        RECT 116.010 172.180 121.690 172.520 ;
        RECT 113.210 171.740 115.570 172.080 ;
        RECT 113.210 159.760 113.550 171.740 ;
        RECT 120.340 171.640 120.680 172.180 ;
        RECT 121.350 172.080 121.690 172.180 ;
        RECT 121.350 171.740 123.210 172.080 ;
        RECT 116.010 171.300 117.090 171.640 ;
        RECT 119.970 171.300 121.050 171.640 ;
        RECT 113.850 170.860 114.930 171.200 ;
        RECT 114.220 170.320 114.560 170.860 ;
        RECT 116.380 170.760 116.720 171.300 ;
        RECT 120.340 170.760 120.680 171.300 ;
        RECT 122.500 171.200 122.840 171.740 ;
        RECT 122.130 170.860 123.210 171.200 ;
        RECT 116.010 170.420 117.090 170.760 ;
        RECT 119.970 170.420 121.050 170.760 ;
        RECT 113.850 169.980 114.930 170.320 ;
        RECT 114.220 169.440 114.560 169.980 ;
        RECT 116.380 169.880 116.720 170.420 ;
        RECT 120.340 169.880 120.680 170.420 ;
        RECT 122.500 170.320 122.840 170.860 ;
        RECT 122.130 169.980 123.210 170.320 ;
        RECT 116.010 169.540 117.090 169.880 ;
        RECT 119.970 169.540 121.050 169.880 ;
        RECT 113.850 169.100 114.930 169.440 ;
        RECT 114.220 168.560 114.560 169.100 ;
        RECT 116.380 169.000 116.720 169.540 ;
        RECT 120.340 169.000 120.680 169.540 ;
        RECT 122.500 169.440 122.840 169.980 ;
        RECT 122.130 169.100 123.210 169.440 ;
        RECT 116.010 168.660 117.090 169.000 ;
        RECT 119.970 168.660 121.050 169.000 ;
        RECT 113.850 168.220 114.930 168.560 ;
        RECT 114.220 167.680 114.560 168.220 ;
        RECT 116.380 168.120 116.720 168.660 ;
        RECT 120.340 168.120 120.680 168.660 ;
        RECT 122.500 168.560 122.840 169.100 ;
        RECT 122.130 168.220 123.210 168.560 ;
        RECT 116.010 167.780 117.090 168.120 ;
        RECT 119.970 167.780 121.050 168.120 ;
        RECT 113.850 167.340 114.930 167.680 ;
        RECT 116.380 167.240 116.720 167.780 ;
        RECT 120.340 167.240 120.680 167.780 ;
        RECT 122.500 167.680 122.840 168.220 ;
        RECT 122.130 167.340 123.210 167.680 ;
        RECT 116.010 166.900 117.730 167.240 ;
        RECT 119.970 166.900 121.050 167.240 ;
        RECT 113.850 166.460 114.930 166.800 ;
        RECT 117.390 166.360 117.730 166.900 ;
        RECT 122.130 166.460 123.210 166.800 ;
        RECT 116.010 166.020 117.090 166.360 ;
        RECT 117.390 166.020 121.050 166.360 ;
        RECT 116.010 165.140 119.670 165.480 ;
        RECT 119.970 165.140 121.050 165.480 ;
        RECT 113.850 164.700 114.930 165.040 ;
        RECT 119.330 164.600 119.670 165.140 ;
        RECT 122.130 164.700 123.210 165.040 ;
        RECT 116.010 164.260 117.730 164.600 ;
        RECT 113.850 163.820 114.930 164.160 ;
        RECT 114.220 163.280 114.560 163.820 ;
        RECT 115.370 163.380 117.090 163.720 ;
        RECT 113.850 162.940 114.930 163.280 ;
        RECT 114.220 162.400 114.560 162.940 ;
        RECT 113.850 162.060 114.930 162.400 ;
        RECT 114.220 161.520 114.560 162.060 ;
        RECT 115.370 161.960 115.710 163.380 ;
        RECT 117.390 162.840 117.730 164.260 ;
        RECT 116.010 162.500 117.730 162.840 ;
        RECT 119.330 164.260 121.050 164.600 ;
        RECT 119.330 162.840 119.670 164.260 ;
        RECT 122.500 164.160 122.840 164.700 ;
        RECT 122.130 163.820 123.210 164.160 ;
        RECT 119.970 163.380 121.050 163.720 ;
        RECT 122.500 163.280 122.840 163.820 ;
        RECT 121.350 162.940 123.210 163.280 ;
        RECT 119.330 162.500 121.050 162.840 ;
        RECT 115.370 161.620 117.090 161.960 ;
        RECT 113.850 161.180 114.930 161.520 ;
        RECT 114.220 160.640 114.560 161.180 ;
        RECT 113.850 160.300 114.930 160.640 ;
        RECT 115.370 160.200 115.710 161.620 ;
        RECT 117.390 161.080 117.730 162.500 ;
        RECT 119.970 161.620 121.050 161.960 ;
        RECT 116.010 160.740 121.050 161.080 ;
        RECT 115.370 159.860 117.730 160.200 ;
        RECT 119.970 159.860 121.050 160.200 ;
        RECT 113.210 159.420 114.930 159.760 ;
        RECT 113.210 143.920 113.550 159.420 ;
        RECT 113.850 157.660 114.930 158.000 ;
        RECT 114.220 157.120 114.560 157.660 ;
        RECT 113.850 156.780 114.930 157.120 ;
        RECT 114.220 156.240 114.560 156.780 ;
        RECT 113.850 155.900 114.930 156.240 ;
        RECT 114.220 155.360 114.560 155.900 ;
        RECT 113.850 155.020 114.930 155.360 ;
        RECT 113.850 153.260 114.930 153.600 ;
        RECT 114.220 152.720 114.560 153.260 ;
        RECT 113.850 152.380 114.930 152.720 ;
        RECT 114.220 151.840 114.560 152.380 ;
        RECT 113.850 151.500 114.930 151.840 ;
        RECT 114.220 150.960 114.560 151.500 ;
        RECT 113.850 150.620 114.930 150.960 ;
        RECT 113.850 148.860 114.930 149.200 ;
        RECT 113.850 147.980 114.930 148.320 ;
        RECT 114.220 147.440 114.560 147.980 ;
        RECT 115.370 147.880 115.710 159.860 ;
        RECT 117.390 159.320 117.730 159.860 ;
        RECT 116.010 158.980 117.090 159.320 ;
        RECT 117.390 158.980 121.050 159.320 ;
        RECT 116.010 158.100 117.090 158.440 ;
        RECT 119.970 158.100 121.050 158.440 ;
        RECT 116.010 157.220 121.050 157.560 ;
        RECT 116.010 156.340 117.090 156.680 ;
        RECT 117.390 155.800 117.730 157.220 ;
        RECT 119.970 156.340 121.050 156.680 ;
        RECT 116.010 155.460 121.050 155.800 ;
        RECT 121.350 155.360 121.690 162.940 ;
        RECT 122.130 162.060 123.850 162.400 ;
        RECT 122.130 161.180 123.210 161.520 ;
        RECT 123.510 160.640 123.850 162.060 ;
        RECT 122.130 160.300 123.850 160.640 ;
        RECT 123.510 159.760 123.850 160.300 ;
        RECT 122.130 159.420 123.850 159.760 ;
        RECT 122.130 157.660 123.210 158.000 ;
        RECT 122.500 157.120 122.840 157.660 ;
        RECT 122.130 156.780 123.210 157.120 ;
        RECT 122.500 156.240 122.840 156.780 ;
        RECT 122.130 155.900 123.210 156.240 ;
        RECT 122.500 155.360 122.840 155.900 ;
        RECT 121.350 155.020 123.210 155.360 ;
        RECT 116.010 154.580 117.090 154.920 ;
        RECT 119.970 154.580 121.050 154.920 ;
        RECT 116.010 153.700 117.090 154.040 ;
        RECT 119.970 153.700 121.050 154.040 ;
        RECT 116.010 152.820 121.050 153.160 ;
        RECT 116.010 151.940 117.090 152.280 ;
        RECT 116.170 151.400 117.090 151.570 ;
        RECT 117.390 151.400 117.730 152.820 ;
        RECT 119.970 151.940 121.050 152.280 ;
        RECT 116.010 151.060 121.050 151.400 ;
        RECT 116.010 150.180 117.090 150.520 ;
        RECT 119.970 150.180 121.050 150.520 ;
        RECT 116.010 149.300 119.670 149.640 ;
        RECT 119.970 149.300 121.050 149.640 ;
        RECT 119.330 148.760 119.670 149.300 ;
        RECT 121.350 148.760 121.690 155.020 ;
        RECT 122.130 153.260 123.210 153.600 ;
        RECT 122.500 152.720 122.840 153.260 ;
        RECT 122.130 152.380 123.210 152.720 ;
        RECT 122.500 151.840 122.840 152.380 ;
        RECT 122.130 151.500 123.210 151.840 ;
        RECT 122.500 150.960 122.840 151.500 ;
        RECT 122.130 150.620 123.210 150.960 ;
        RECT 122.130 148.860 123.210 149.200 ;
        RECT 116.010 148.420 117.730 148.760 ;
        RECT 115.370 147.540 117.090 147.880 ;
        RECT 113.850 147.100 114.930 147.440 ;
        RECT 114.220 146.560 114.560 147.100 ;
        RECT 113.850 146.220 114.930 146.560 ;
        RECT 114.220 145.680 114.560 146.220 ;
        RECT 115.370 146.120 115.710 147.540 ;
        RECT 117.390 147.000 117.730 148.420 ;
        RECT 116.010 146.660 117.730 147.000 ;
        RECT 119.330 148.420 121.690 148.760 ;
        RECT 119.330 147.000 119.670 148.420 ;
        RECT 122.500 148.320 122.840 148.860 ;
        RECT 122.130 147.980 123.210 148.320 ;
        RECT 119.970 147.540 121.050 147.880 ;
        RECT 122.500 147.440 122.840 147.980 ;
        RECT 122.130 147.100 123.210 147.440 ;
        RECT 119.330 146.660 121.050 147.000 ;
        RECT 115.370 145.780 117.090 146.120 ;
        RECT 113.850 145.340 114.930 145.680 ;
        RECT 114.220 144.800 114.560 145.340 ;
        RECT 113.850 144.460 114.930 144.800 ;
        RECT 115.370 144.360 115.710 145.780 ;
        RECT 117.390 145.240 117.730 146.660 ;
        RECT 122.130 146.220 123.850 146.560 ;
        RECT 119.970 145.780 121.050 146.120 ;
        RECT 122.130 145.340 123.210 145.680 ;
        RECT 116.010 144.900 121.050 145.240 ;
        RECT 123.510 144.800 123.850 146.220 ;
        RECT 122.130 144.460 123.850 144.800 ;
        RECT 115.370 144.020 117.730 144.360 ;
        RECT 119.970 144.020 121.050 144.360 ;
        RECT 113.210 143.580 114.930 143.920 ;
        RECT 113.210 142.160 113.550 143.580 ;
        RECT 117.390 143.480 117.730 144.020 ;
        RECT 123.510 143.920 123.850 144.460 ;
        RECT 122.130 143.580 123.850 143.920 ;
        RECT 116.010 143.140 117.090 143.480 ;
        RECT 117.390 143.140 121.050 143.480 ;
        RECT 116.010 142.260 121.690 142.600 ;
        RECT 113.210 141.820 114.930 142.160 ;
        RECT 120.340 141.720 120.680 142.260 ;
        RECT 121.350 142.160 121.690 142.260 ;
        RECT 121.350 141.820 123.210 142.160 ;
        RECT 116.010 141.380 117.090 141.720 ;
        RECT 119.970 141.380 121.050 141.720 ;
        RECT 113.850 140.940 114.930 141.280 ;
        RECT 114.220 140.400 114.560 140.940 ;
        RECT 116.380 140.840 116.720 141.380 ;
        RECT 120.340 140.840 120.680 141.380 ;
        RECT 122.500 141.280 122.840 141.820 ;
        RECT 122.130 140.940 123.210 141.280 ;
        RECT 116.010 140.500 117.090 140.840 ;
        RECT 119.970 140.500 121.050 140.840 ;
        RECT 113.850 140.060 114.930 140.400 ;
        RECT 114.220 139.520 114.560 140.060 ;
        RECT 116.380 139.960 116.720 140.500 ;
        RECT 120.340 139.960 120.680 140.500 ;
        RECT 122.500 140.400 122.840 140.940 ;
        RECT 122.130 140.060 123.210 140.400 ;
        RECT 116.010 139.620 117.090 139.960 ;
        RECT 119.970 139.620 121.050 139.960 ;
        RECT 113.850 139.180 114.930 139.520 ;
        RECT 114.220 138.640 114.560 139.180 ;
        RECT 116.380 139.080 116.720 139.620 ;
        RECT 120.340 139.080 120.680 139.620 ;
        RECT 122.500 139.520 122.840 140.060 ;
        RECT 122.130 139.180 123.210 139.520 ;
        RECT 116.010 138.740 117.090 139.080 ;
        RECT 119.970 138.740 121.050 139.080 ;
        RECT 113.850 138.300 114.930 138.640 ;
        RECT 114.220 137.760 114.560 138.300 ;
        RECT 116.380 138.200 116.720 138.740 ;
        RECT 120.340 138.200 120.680 138.740 ;
        RECT 122.500 138.640 122.840 139.180 ;
        RECT 122.130 138.300 123.210 138.640 ;
        RECT 116.010 137.860 117.090 138.200 ;
        RECT 119.970 137.860 121.050 138.200 ;
        RECT 113.850 137.420 114.930 137.760 ;
        RECT 116.380 137.320 116.720 137.860 ;
        RECT 120.340 137.320 120.680 137.860 ;
        RECT 122.500 137.760 122.840 138.300 ;
        RECT 122.130 137.420 123.210 137.760 ;
        RECT 116.010 136.980 117.730 137.320 ;
        RECT 119.970 136.980 121.050 137.320 ;
        RECT 113.850 136.540 114.930 136.880 ;
        RECT 117.390 136.440 117.730 136.980 ;
        RECT 122.130 136.540 123.210 136.880 ;
        RECT 116.010 136.100 117.090 136.440 ;
        RECT 117.390 136.100 121.050 136.440 ;
        RECT 115.230 135.220 117.090 135.560 ;
        RECT 119.970 135.220 121.690 135.560 ;
        RECT 115.230 135.120 115.570 135.220 ;
        RECT 108.890 134.780 115.570 135.120 ;
        RECT 108.890 134.680 109.230 134.780 ;
        RECT 102.770 134.340 104.490 134.680 ;
        RECT 107.370 134.340 109.230 134.680 ;
        RECT 111.690 133.850 112.770 134.780 ;
        RECT 115.230 134.680 115.570 134.780 ;
        RECT 121.350 135.120 121.690 135.220 ;
        RECT 124.290 135.120 125.370 182.300 ;
        RECT 121.350 134.780 125.370 135.120 ;
        RECT 121.350 134.680 121.690 134.780 ;
        RECT 115.230 134.340 117.090 134.680 ;
        RECT 119.970 134.340 121.690 134.680 ;
        RECT 124.290 133.850 125.370 134.780 ;
        RECT 22.800 105.560 23.140 105.850 ;
        RECT 113.120 105.560 113.460 105.850 ;
        RECT 13.240 105.220 55.440 105.560 ;
        RECT 55.780 105.220 57.040 105.560 ;
        RECT 79.220 105.220 80.480 105.560 ;
        RECT 80.820 105.220 123.020 105.560 ;
        RECT 22.800 104.930 23.140 105.220 ;
        RECT 113.120 104.930 113.460 105.220 ;
        RECT 21.480 102.540 21.820 102.830 ;
        RECT 25.440 102.540 25.780 102.830 ;
        RECT 42.600 102.540 42.940 102.830 ;
        RECT 46.560 102.540 46.900 102.830 ;
        RECT 89.360 102.540 89.700 102.830 ;
        RECT 93.320 102.540 93.660 102.830 ;
        RECT 110.480 102.540 110.820 102.830 ;
        RECT 114.440 102.540 114.780 102.830 ;
        RECT 13.240 102.200 55.440 102.540 ;
        RECT 55.780 102.200 57.040 102.540 ;
        RECT 79.220 102.200 80.480 102.540 ;
        RECT 80.820 102.200 123.020 102.540 ;
        RECT 21.480 101.910 21.820 102.200 ;
        RECT 25.440 101.910 25.780 102.200 ;
        RECT 42.600 101.910 42.940 102.200 ;
        RECT 46.560 101.910 46.900 102.200 ;
        RECT 89.360 101.910 89.700 102.200 ;
        RECT 93.320 101.910 93.660 102.200 ;
        RECT 110.480 101.910 110.820 102.200 ;
        RECT 114.440 101.910 114.780 102.200 ;
        RECT 18.840 99.520 19.180 99.810 ;
        RECT 20.160 99.520 20.500 99.810 ;
        RECT 26.760 99.520 27.100 99.810 ;
        RECT 28.080 99.520 28.420 99.810 ;
        RECT 39.960 99.520 40.300 99.810 ;
        RECT 41.280 99.520 41.620 99.810 ;
        RECT 47.880 99.520 48.220 99.810 ;
        RECT 49.200 99.520 49.540 99.810 ;
        RECT 86.720 99.520 87.060 99.810 ;
        RECT 88.040 99.520 88.380 99.810 ;
        RECT 94.640 99.520 94.980 99.810 ;
        RECT 95.960 99.520 96.300 99.810 ;
        RECT 107.840 99.520 108.180 99.810 ;
        RECT 109.160 99.520 109.500 99.810 ;
        RECT 115.760 99.520 116.100 99.810 ;
        RECT 117.080 99.520 117.420 99.810 ;
        RECT 13.240 99.180 55.440 99.520 ;
        RECT 55.780 99.180 57.040 99.520 ;
        RECT 79.220 99.180 80.480 99.520 ;
        RECT 80.820 99.180 123.020 99.520 ;
        RECT 18.840 98.890 19.180 99.180 ;
        RECT 20.160 98.890 20.500 99.180 ;
        RECT 26.760 98.890 27.100 99.180 ;
        RECT 28.080 98.890 28.420 99.180 ;
        RECT 39.960 98.890 40.300 99.180 ;
        RECT 41.280 98.890 41.620 99.180 ;
        RECT 47.880 98.890 48.220 99.180 ;
        RECT 49.200 98.890 49.540 99.180 ;
        RECT 86.720 98.890 87.060 99.180 ;
        RECT 88.040 98.890 88.380 99.180 ;
        RECT 94.640 98.890 94.980 99.180 ;
        RECT 95.960 98.890 96.300 99.180 ;
        RECT 107.840 98.890 108.180 99.180 ;
        RECT 109.160 98.890 109.500 99.180 ;
        RECT 115.760 98.890 116.100 99.180 ;
        RECT 117.080 98.890 117.420 99.180 ;
        RECT 24.120 96.500 24.460 96.790 ;
        RECT 43.920 96.500 44.260 96.790 ;
        RECT 92.000 96.500 92.340 96.790 ;
        RECT 111.800 96.500 112.140 96.790 ;
        RECT 13.240 96.160 55.440 96.500 ;
        RECT 55.780 96.160 57.040 96.500 ;
        RECT 79.220 96.160 80.480 96.500 ;
        RECT 80.820 96.160 123.020 96.500 ;
        RECT 24.120 95.870 24.460 96.160 ;
        RECT 43.920 95.870 44.260 96.160 ;
        RECT 92.000 95.870 92.340 96.160 ;
        RECT 111.800 95.870 112.140 96.160 ;
        RECT 13.560 93.480 13.900 93.770 ;
        RECT 14.880 93.480 15.220 93.770 ;
        RECT 16.200 93.480 16.540 93.770 ;
        RECT 17.520 93.480 17.860 93.770 ;
        RECT 29.400 93.480 29.740 93.770 ;
        RECT 30.720 93.480 31.060 93.770 ;
        RECT 32.040 93.480 32.380 93.770 ;
        RECT 33.360 93.480 33.700 93.770 ;
        RECT 34.680 93.480 35.020 93.770 ;
        RECT 36.000 93.480 36.340 93.770 ;
        RECT 37.320 93.480 37.660 93.770 ;
        RECT 38.640 93.480 38.980 93.770 ;
        RECT 50.520 93.480 50.860 93.770 ;
        RECT 51.840 93.480 52.180 93.770 ;
        RECT 53.160 93.480 53.500 93.770 ;
        RECT 54.480 93.480 54.820 93.770 ;
        RECT 81.440 93.480 81.780 93.770 ;
        RECT 82.760 93.480 83.100 93.770 ;
        RECT 84.080 93.480 84.420 93.770 ;
        RECT 85.400 93.480 85.740 93.770 ;
        RECT 97.280 93.480 97.620 93.770 ;
        RECT 98.600 93.480 98.940 93.770 ;
        RECT 99.920 93.480 100.260 93.770 ;
        RECT 101.240 93.480 101.580 93.770 ;
        RECT 102.560 93.480 102.900 93.770 ;
        RECT 103.880 93.480 104.220 93.770 ;
        RECT 105.200 93.480 105.540 93.770 ;
        RECT 106.520 93.480 106.860 93.770 ;
        RECT 118.400 93.480 118.740 93.770 ;
        RECT 119.720 93.480 120.060 93.770 ;
        RECT 121.040 93.480 121.380 93.770 ;
        RECT 122.360 93.480 122.700 93.770 ;
        RECT 13.240 93.140 55.440 93.480 ;
        RECT 55.780 93.140 57.040 93.480 ;
        RECT 79.220 93.140 80.480 93.480 ;
        RECT 80.820 93.140 123.020 93.480 ;
        RECT 13.560 92.850 13.900 93.140 ;
        RECT 14.880 92.850 15.220 93.140 ;
        RECT 16.200 92.850 16.540 93.140 ;
        RECT 17.520 92.850 17.860 93.140 ;
        RECT 29.400 92.850 29.740 93.140 ;
        RECT 30.720 92.850 31.060 93.140 ;
        RECT 32.040 92.850 32.380 93.140 ;
        RECT 33.360 92.850 33.700 93.140 ;
        RECT 34.680 92.850 35.020 93.140 ;
        RECT 36.000 92.850 36.340 93.140 ;
        RECT 37.320 92.850 37.660 93.140 ;
        RECT 38.640 92.850 38.980 93.140 ;
        RECT 50.520 92.850 50.860 93.140 ;
        RECT 51.840 92.850 52.180 93.140 ;
        RECT 53.160 92.850 53.500 93.140 ;
        RECT 54.480 92.850 54.820 93.140 ;
        RECT 81.440 92.850 81.780 93.140 ;
        RECT 82.760 92.850 83.100 93.140 ;
        RECT 84.080 92.850 84.420 93.140 ;
        RECT 85.400 92.850 85.740 93.140 ;
        RECT 97.280 92.850 97.620 93.140 ;
        RECT 98.600 92.850 98.940 93.140 ;
        RECT 99.920 92.850 100.260 93.140 ;
        RECT 101.240 92.850 101.580 93.140 ;
        RECT 102.560 92.850 102.900 93.140 ;
        RECT 103.880 92.850 104.220 93.140 ;
        RECT 105.200 92.850 105.540 93.140 ;
        RECT 106.520 92.850 106.860 93.140 ;
        RECT 118.400 92.850 118.740 93.140 ;
        RECT 119.720 92.850 120.060 93.140 ;
        RECT 121.040 92.850 121.380 93.140 ;
        RECT 122.360 92.850 122.700 93.140 ;
        RECT 45.240 90.460 45.580 90.750 ;
        RECT 90.680 90.460 91.020 90.750 ;
        RECT 13.240 90.120 55.440 90.460 ;
        RECT 55.780 90.120 57.040 90.460 ;
        RECT 79.220 90.120 80.480 90.460 ;
        RECT 80.820 90.120 123.020 90.460 ;
        RECT 45.240 89.830 45.580 90.120 ;
        RECT 90.680 89.830 91.020 90.120 ;
        RECT 22.800 88.560 23.140 88.850 ;
        RECT 113.120 88.560 113.460 88.850 ;
        RECT 13.240 88.220 55.440 88.560 ;
        RECT 55.780 88.220 57.040 88.560 ;
        RECT 79.220 88.220 80.480 88.560 ;
        RECT 80.820 88.220 123.020 88.560 ;
        RECT 22.800 87.930 23.140 88.220 ;
        RECT 113.120 87.930 113.460 88.220 ;
        RECT 21.480 85.540 21.820 85.830 ;
        RECT 25.440 85.540 25.780 85.830 ;
        RECT 42.600 85.540 42.940 85.830 ;
        RECT 46.560 85.540 46.900 85.830 ;
        RECT 89.360 85.540 89.700 85.830 ;
        RECT 93.320 85.540 93.660 85.830 ;
        RECT 110.480 85.540 110.820 85.830 ;
        RECT 114.440 85.540 114.780 85.830 ;
        RECT 13.240 85.200 55.440 85.540 ;
        RECT 55.780 85.200 57.040 85.540 ;
        RECT 79.220 85.200 80.480 85.540 ;
        RECT 80.820 85.200 123.020 85.540 ;
        RECT 21.480 84.910 21.820 85.200 ;
        RECT 25.440 84.910 25.780 85.200 ;
        RECT 42.600 84.910 42.940 85.200 ;
        RECT 46.560 84.910 46.900 85.200 ;
        RECT 89.360 84.910 89.700 85.200 ;
        RECT 93.320 84.910 93.660 85.200 ;
        RECT 110.480 84.910 110.820 85.200 ;
        RECT 114.440 84.910 114.780 85.200 ;
        RECT 18.840 82.520 19.180 82.810 ;
        RECT 20.160 82.520 20.500 82.810 ;
        RECT 26.760 82.520 27.100 82.810 ;
        RECT 28.080 82.520 28.420 82.810 ;
        RECT 39.960 82.520 40.300 82.810 ;
        RECT 41.280 82.520 41.620 82.810 ;
        RECT 47.880 82.520 48.220 82.810 ;
        RECT 49.200 82.520 49.540 82.810 ;
        RECT 86.720 82.520 87.060 82.810 ;
        RECT 88.040 82.520 88.380 82.810 ;
        RECT 94.640 82.520 94.980 82.810 ;
        RECT 95.960 82.520 96.300 82.810 ;
        RECT 107.840 82.520 108.180 82.810 ;
        RECT 109.160 82.520 109.500 82.810 ;
        RECT 115.760 82.520 116.100 82.810 ;
        RECT 117.080 82.520 117.420 82.810 ;
        RECT 13.240 82.180 55.440 82.520 ;
        RECT 55.780 82.180 57.040 82.520 ;
        RECT 79.220 82.180 80.480 82.520 ;
        RECT 80.820 82.180 123.020 82.520 ;
        RECT 18.840 81.890 19.180 82.180 ;
        RECT 20.160 81.890 20.500 82.180 ;
        RECT 26.760 81.890 27.100 82.180 ;
        RECT 28.080 81.890 28.420 82.180 ;
        RECT 39.960 81.890 40.300 82.180 ;
        RECT 41.280 81.890 41.620 82.180 ;
        RECT 47.880 81.890 48.220 82.180 ;
        RECT 49.200 81.890 49.540 82.180 ;
        RECT 86.720 81.890 87.060 82.180 ;
        RECT 88.040 81.890 88.380 82.180 ;
        RECT 94.640 81.890 94.980 82.180 ;
        RECT 95.960 81.890 96.300 82.180 ;
        RECT 107.840 81.890 108.180 82.180 ;
        RECT 109.160 81.890 109.500 82.180 ;
        RECT 115.760 81.890 116.100 82.180 ;
        RECT 117.080 81.890 117.420 82.180 ;
        RECT 24.120 79.500 24.460 79.790 ;
        RECT 43.920 79.500 44.260 79.790 ;
        RECT 92.000 79.500 92.340 79.790 ;
        RECT 111.800 79.500 112.140 79.790 ;
        RECT 13.240 79.160 55.440 79.500 ;
        RECT 55.780 79.160 57.040 79.500 ;
        RECT 79.220 79.160 80.480 79.500 ;
        RECT 80.820 79.160 123.020 79.500 ;
        RECT 24.120 78.870 24.460 79.160 ;
        RECT 43.920 78.870 44.260 79.160 ;
        RECT 92.000 78.870 92.340 79.160 ;
        RECT 111.800 78.870 112.140 79.160 ;
        RECT 13.560 76.480 13.900 76.770 ;
        RECT 14.880 76.480 15.220 76.770 ;
        RECT 16.200 76.480 16.540 76.770 ;
        RECT 17.520 76.480 17.860 76.770 ;
        RECT 29.400 76.480 29.740 76.770 ;
        RECT 30.720 76.480 31.060 76.770 ;
        RECT 32.040 76.480 32.380 76.770 ;
        RECT 33.360 76.480 33.700 76.770 ;
        RECT 34.680 76.480 35.020 76.770 ;
        RECT 36.000 76.480 36.340 76.770 ;
        RECT 37.320 76.480 37.660 76.770 ;
        RECT 38.640 76.480 38.980 76.770 ;
        RECT 50.520 76.480 50.860 76.770 ;
        RECT 51.840 76.480 52.180 76.770 ;
        RECT 53.160 76.480 53.500 76.770 ;
        RECT 54.480 76.480 54.820 76.770 ;
        RECT 81.440 76.480 81.780 76.770 ;
        RECT 82.760 76.480 83.100 76.770 ;
        RECT 84.080 76.480 84.420 76.770 ;
        RECT 85.400 76.480 85.740 76.770 ;
        RECT 97.280 76.480 97.620 76.770 ;
        RECT 98.600 76.480 98.940 76.770 ;
        RECT 99.920 76.480 100.260 76.770 ;
        RECT 101.240 76.480 101.580 76.770 ;
        RECT 102.560 76.480 102.900 76.770 ;
        RECT 103.880 76.480 104.220 76.770 ;
        RECT 105.200 76.480 105.540 76.770 ;
        RECT 106.520 76.480 106.860 76.770 ;
        RECT 118.400 76.480 118.740 76.770 ;
        RECT 119.720 76.480 120.060 76.770 ;
        RECT 121.040 76.480 121.380 76.770 ;
        RECT 122.360 76.480 122.700 76.770 ;
        RECT 13.240 76.140 55.440 76.480 ;
        RECT 55.780 76.140 57.040 76.480 ;
        RECT 79.220 76.140 80.480 76.480 ;
        RECT 80.820 76.140 123.020 76.480 ;
        RECT 13.560 75.850 13.900 76.140 ;
        RECT 14.880 75.850 15.220 76.140 ;
        RECT 16.200 75.850 16.540 76.140 ;
        RECT 17.520 75.850 17.860 76.140 ;
        RECT 29.400 75.850 29.740 76.140 ;
        RECT 30.720 75.850 31.060 76.140 ;
        RECT 32.040 75.850 32.380 76.140 ;
        RECT 33.360 75.850 33.700 76.140 ;
        RECT 34.680 75.850 35.020 76.140 ;
        RECT 36.000 75.850 36.340 76.140 ;
        RECT 37.320 75.850 37.660 76.140 ;
        RECT 38.640 75.850 38.980 76.140 ;
        RECT 50.520 75.850 50.860 76.140 ;
        RECT 51.840 75.850 52.180 76.140 ;
        RECT 53.160 75.850 53.500 76.140 ;
        RECT 54.480 75.850 54.820 76.140 ;
        RECT 81.440 75.850 81.780 76.140 ;
        RECT 82.760 75.850 83.100 76.140 ;
        RECT 84.080 75.850 84.420 76.140 ;
        RECT 85.400 75.850 85.740 76.140 ;
        RECT 97.280 75.850 97.620 76.140 ;
        RECT 98.600 75.850 98.940 76.140 ;
        RECT 99.920 75.850 100.260 76.140 ;
        RECT 101.240 75.850 101.580 76.140 ;
        RECT 102.560 75.850 102.900 76.140 ;
        RECT 103.880 75.850 104.220 76.140 ;
        RECT 105.200 75.850 105.540 76.140 ;
        RECT 106.520 75.850 106.860 76.140 ;
        RECT 118.400 75.850 118.740 76.140 ;
        RECT 119.720 75.850 120.060 76.140 ;
        RECT 121.040 75.850 121.380 76.140 ;
        RECT 122.360 75.850 122.700 76.140 ;
        RECT 45.240 73.460 45.580 73.750 ;
        RECT 90.680 73.460 91.020 73.750 ;
        RECT 13.240 73.120 55.440 73.460 ;
        RECT 55.780 73.120 57.040 73.460 ;
        RECT 79.220 73.120 80.480 73.460 ;
        RECT 80.820 73.120 123.020 73.460 ;
        RECT 45.240 72.830 45.580 73.120 ;
        RECT 90.680 72.830 91.020 73.120 ;
        RECT 22.800 71.560 23.140 71.850 ;
        RECT 113.120 71.560 113.460 71.850 ;
        RECT 13.240 71.220 55.440 71.560 ;
        RECT 55.780 71.220 57.040 71.560 ;
        RECT 79.220 71.220 80.480 71.560 ;
        RECT 80.820 71.220 123.020 71.560 ;
        RECT 22.800 70.930 23.140 71.220 ;
        RECT 113.120 70.930 113.460 71.220 ;
        RECT 21.480 68.540 21.820 68.830 ;
        RECT 25.440 68.540 25.780 68.830 ;
        RECT 42.600 68.540 42.940 68.830 ;
        RECT 46.560 68.540 46.900 68.830 ;
        RECT 89.360 68.540 89.700 68.830 ;
        RECT 93.320 68.540 93.660 68.830 ;
        RECT 110.480 68.540 110.820 68.830 ;
        RECT 114.440 68.540 114.780 68.830 ;
        RECT 13.240 68.200 55.440 68.540 ;
        RECT 55.780 68.200 57.040 68.540 ;
        RECT 79.220 68.200 80.480 68.540 ;
        RECT 80.820 68.200 123.020 68.540 ;
        RECT 21.480 67.910 21.820 68.200 ;
        RECT 25.440 67.910 25.780 68.200 ;
        RECT 42.600 67.910 42.940 68.200 ;
        RECT 46.560 67.910 46.900 68.200 ;
        RECT 89.360 67.910 89.700 68.200 ;
        RECT 93.320 67.910 93.660 68.200 ;
        RECT 110.480 67.910 110.820 68.200 ;
        RECT 114.440 67.910 114.780 68.200 ;
        RECT 18.840 65.520 19.180 65.810 ;
        RECT 20.160 65.520 20.500 65.810 ;
        RECT 26.760 65.520 27.100 65.810 ;
        RECT 28.080 65.520 28.420 65.810 ;
        RECT 39.960 65.520 40.300 65.810 ;
        RECT 41.280 65.520 41.620 65.810 ;
        RECT 47.880 65.520 48.220 65.810 ;
        RECT 49.200 65.520 49.540 65.810 ;
        RECT 86.720 65.520 87.060 65.810 ;
        RECT 88.040 65.520 88.380 65.810 ;
        RECT 94.640 65.520 94.980 65.810 ;
        RECT 95.960 65.520 96.300 65.810 ;
        RECT 107.840 65.520 108.180 65.810 ;
        RECT 109.160 65.520 109.500 65.810 ;
        RECT 115.760 65.520 116.100 65.810 ;
        RECT 117.080 65.520 117.420 65.810 ;
        RECT 13.240 65.180 55.440 65.520 ;
        RECT 55.780 65.180 57.040 65.520 ;
        RECT 79.220 65.180 80.480 65.520 ;
        RECT 80.820 65.180 123.020 65.520 ;
        RECT 18.840 64.890 19.180 65.180 ;
        RECT 20.160 64.890 20.500 65.180 ;
        RECT 26.760 64.890 27.100 65.180 ;
        RECT 28.080 64.890 28.420 65.180 ;
        RECT 39.960 64.890 40.300 65.180 ;
        RECT 41.280 64.890 41.620 65.180 ;
        RECT 47.880 64.890 48.220 65.180 ;
        RECT 49.200 64.890 49.540 65.180 ;
        RECT 86.720 64.890 87.060 65.180 ;
        RECT 88.040 64.890 88.380 65.180 ;
        RECT 94.640 64.890 94.980 65.180 ;
        RECT 95.960 64.890 96.300 65.180 ;
        RECT 107.840 64.890 108.180 65.180 ;
        RECT 109.160 64.890 109.500 65.180 ;
        RECT 115.760 64.890 116.100 65.180 ;
        RECT 117.080 64.890 117.420 65.180 ;
        RECT 24.120 62.500 24.460 62.790 ;
        RECT 43.920 62.500 44.260 62.790 ;
        RECT 92.000 62.500 92.340 62.790 ;
        RECT 111.800 62.500 112.140 62.790 ;
        RECT 13.240 62.160 55.440 62.500 ;
        RECT 55.780 62.160 57.040 62.500 ;
        RECT 79.220 62.160 80.480 62.500 ;
        RECT 80.820 62.160 123.020 62.500 ;
        RECT 24.120 61.870 24.460 62.160 ;
        RECT 43.920 61.870 44.260 62.160 ;
        RECT 92.000 61.870 92.340 62.160 ;
        RECT 111.800 61.870 112.140 62.160 ;
        RECT 13.560 59.480 13.900 59.770 ;
        RECT 14.880 59.480 15.220 59.770 ;
        RECT 16.200 59.480 16.540 59.770 ;
        RECT 17.520 59.480 17.860 59.770 ;
        RECT 29.400 59.480 29.740 59.770 ;
        RECT 30.720 59.480 31.060 59.770 ;
        RECT 32.040 59.480 32.380 59.770 ;
        RECT 33.360 59.480 33.700 59.770 ;
        RECT 34.680 59.480 35.020 59.770 ;
        RECT 36.000 59.480 36.340 59.770 ;
        RECT 37.320 59.480 37.660 59.770 ;
        RECT 38.640 59.480 38.980 59.770 ;
        RECT 50.520 59.480 50.860 59.770 ;
        RECT 51.840 59.480 52.180 59.770 ;
        RECT 53.160 59.480 53.500 59.770 ;
        RECT 54.480 59.480 54.820 59.770 ;
        RECT 81.440 59.480 81.780 59.770 ;
        RECT 82.760 59.480 83.100 59.770 ;
        RECT 84.080 59.480 84.420 59.770 ;
        RECT 85.400 59.480 85.740 59.770 ;
        RECT 97.280 59.480 97.620 59.770 ;
        RECT 98.600 59.480 98.940 59.770 ;
        RECT 99.920 59.480 100.260 59.770 ;
        RECT 101.240 59.480 101.580 59.770 ;
        RECT 102.560 59.480 102.900 59.770 ;
        RECT 103.880 59.480 104.220 59.770 ;
        RECT 105.200 59.480 105.540 59.770 ;
        RECT 106.520 59.480 106.860 59.770 ;
        RECT 118.400 59.480 118.740 59.770 ;
        RECT 119.720 59.480 120.060 59.770 ;
        RECT 121.040 59.480 121.380 59.770 ;
        RECT 122.360 59.480 122.700 59.770 ;
        RECT 13.240 59.140 55.440 59.480 ;
        RECT 55.780 59.140 57.040 59.480 ;
        RECT 79.220 59.140 80.480 59.480 ;
        RECT 80.820 59.140 123.020 59.480 ;
        RECT 13.560 58.850 13.900 59.140 ;
        RECT 14.880 58.850 15.220 59.140 ;
        RECT 16.200 58.850 16.540 59.140 ;
        RECT 17.520 58.850 17.860 59.140 ;
        RECT 29.400 58.850 29.740 59.140 ;
        RECT 30.720 58.850 31.060 59.140 ;
        RECT 32.040 58.850 32.380 59.140 ;
        RECT 33.360 58.850 33.700 59.140 ;
        RECT 34.680 58.850 35.020 59.140 ;
        RECT 36.000 58.850 36.340 59.140 ;
        RECT 37.320 58.850 37.660 59.140 ;
        RECT 38.640 58.850 38.980 59.140 ;
        RECT 50.520 58.850 50.860 59.140 ;
        RECT 51.840 58.850 52.180 59.140 ;
        RECT 53.160 58.850 53.500 59.140 ;
        RECT 54.480 58.850 54.820 59.140 ;
        RECT 81.440 58.850 81.780 59.140 ;
        RECT 82.760 58.850 83.100 59.140 ;
        RECT 84.080 58.850 84.420 59.140 ;
        RECT 85.400 58.850 85.740 59.140 ;
        RECT 97.280 58.850 97.620 59.140 ;
        RECT 98.600 58.850 98.940 59.140 ;
        RECT 99.920 58.850 100.260 59.140 ;
        RECT 101.240 58.850 101.580 59.140 ;
        RECT 102.560 58.850 102.900 59.140 ;
        RECT 103.880 58.850 104.220 59.140 ;
        RECT 105.200 58.850 105.540 59.140 ;
        RECT 106.520 58.850 106.860 59.140 ;
        RECT 118.400 58.850 118.740 59.140 ;
        RECT 119.720 58.850 120.060 59.140 ;
        RECT 121.040 58.850 121.380 59.140 ;
        RECT 122.360 58.850 122.700 59.140 ;
        RECT 45.240 56.460 45.580 56.750 ;
        RECT 56.700 56.460 57.040 56.750 ;
        RECT 13.240 56.120 55.440 56.460 ;
        RECT 55.780 56.120 57.040 56.460 ;
        RECT 45.240 55.830 45.580 56.120 ;
        RECT 56.700 55.830 57.040 56.120 ;
        RECT 79.220 56.460 79.560 56.750 ;
        RECT 90.680 56.460 91.020 56.750 ;
        RECT 79.220 56.120 80.480 56.460 ;
        RECT 80.820 56.120 123.020 56.460 ;
        RECT 79.220 55.830 79.560 56.120 ;
        RECT 90.680 55.830 91.020 56.120 ;
        RECT 22.800 54.560 23.140 54.850 ;
        RECT 113.120 54.560 113.460 54.850 ;
        RECT 13.240 54.220 55.440 54.560 ;
        RECT 55.780 54.220 57.040 54.560 ;
        RECT 79.220 54.220 80.480 54.560 ;
        RECT 80.820 54.220 123.020 54.560 ;
        RECT 22.800 53.930 23.140 54.220 ;
        RECT 113.120 53.930 113.460 54.220 ;
        RECT 21.480 51.540 21.820 51.830 ;
        RECT 25.440 51.540 25.780 51.830 ;
        RECT 42.600 51.540 42.940 51.830 ;
        RECT 46.560 51.540 46.900 51.830 ;
        RECT 89.360 51.540 89.700 51.830 ;
        RECT 93.320 51.540 93.660 51.830 ;
        RECT 110.480 51.540 110.820 51.830 ;
        RECT 114.440 51.540 114.780 51.830 ;
        RECT 13.240 51.200 55.440 51.540 ;
        RECT 55.780 51.200 57.040 51.540 ;
        RECT 79.220 51.200 80.480 51.540 ;
        RECT 80.820 51.200 123.020 51.540 ;
        RECT 21.480 50.910 21.820 51.200 ;
        RECT 25.440 50.910 25.780 51.200 ;
        RECT 42.600 50.910 42.940 51.200 ;
        RECT 46.560 50.910 46.900 51.200 ;
        RECT 89.360 50.910 89.700 51.200 ;
        RECT 93.320 50.910 93.660 51.200 ;
        RECT 110.480 50.910 110.820 51.200 ;
        RECT 114.440 50.910 114.780 51.200 ;
        RECT 18.840 48.520 19.180 48.810 ;
        RECT 20.160 48.520 20.500 48.810 ;
        RECT 26.760 48.520 27.100 48.810 ;
        RECT 28.080 48.520 28.420 48.810 ;
        RECT 39.960 48.520 40.300 48.810 ;
        RECT 41.280 48.520 41.620 48.810 ;
        RECT 47.880 48.520 48.220 48.810 ;
        RECT 49.200 48.520 49.540 48.810 ;
        RECT 86.720 48.520 87.060 48.810 ;
        RECT 88.040 48.520 88.380 48.810 ;
        RECT 94.640 48.520 94.980 48.810 ;
        RECT 95.960 48.520 96.300 48.810 ;
        RECT 107.840 48.520 108.180 48.810 ;
        RECT 109.160 48.520 109.500 48.810 ;
        RECT 115.760 48.520 116.100 48.810 ;
        RECT 117.080 48.520 117.420 48.810 ;
        RECT 13.240 48.180 55.440 48.520 ;
        RECT 55.780 48.180 57.040 48.520 ;
        RECT 79.220 48.180 80.480 48.520 ;
        RECT 80.820 48.180 123.020 48.520 ;
        RECT 18.840 47.890 19.180 48.180 ;
        RECT 20.160 47.890 20.500 48.180 ;
        RECT 26.760 47.890 27.100 48.180 ;
        RECT 28.080 47.890 28.420 48.180 ;
        RECT 39.960 47.890 40.300 48.180 ;
        RECT 41.280 47.890 41.620 48.180 ;
        RECT 47.880 47.890 48.220 48.180 ;
        RECT 49.200 47.890 49.540 48.180 ;
        RECT 86.720 47.890 87.060 48.180 ;
        RECT 88.040 47.890 88.380 48.180 ;
        RECT 94.640 47.890 94.980 48.180 ;
        RECT 95.960 47.890 96.300 48.180 ;
        RECT 107.840 47.890 108.180 48.180 ;
        RECT 109.160 47.890 109.500 48.180 ;
        RECT 115.760 47.890 116.100 48.180 ;
        RECT 117.080 47.890 117.420 48.180 ;
        RECT 24.120 45.500 24.460 45.790 ;
        RECT 43.920 45.500 44.260 45.790 ;
        RECT 92.000 45.500 92.340 45.790 ;
        RECT 111.800 45.500 112.140 45.790 ;
        RECT 13.240 45.160 55.440 45.500 ;
        RECT 55.780 45.160 57.040 45.500 ;
        RECT 79.220 45.160 80.480 45.500 ;
        RECT 80.820 45.160 123.020 45.500 ;
        RECT 24.120 44.870 24.460 45.160 ;
        RECT 43.920 44.870 44.260 45.160 ;
        RECT 92.000 44.870 92.340 45.160 ;
        RECT 111.800 44.870 112.140 45.160 ;
        RECT 13.560 42.480 13.900 42.770 ;
        RECT 14.880 42.480 15.220 42.770 ;
        RECT 16.200 42.480 16.540 42.770 ;
        RECT 17.520 42.480 17.860 42.770 ;
        RECT 29.400 42.480 29.740 42.770 ;
        RECT 30.720 42.480 31.060 42.770 ;
        RECT 32.040 42.480 32.380 42.770 ;
        RECT 33.360 42.480 33.700 42.770 ;
        RECT 34.680 42.480 35.020 42.770 ;
        RECT 36.000 42.480 36.340 42.770 ;
        RECT 37.320 42.480 37.660 42.770 ;
        RECT 38.640 42.480 38.980 42.770 ;
        RECT 50.520 42.480 50.860 42.770 ;
        RECT 51.840 42.480 52.180 42.770 ;
        RECT 53.160 42.480 53.500 42.770 ;
        RECT 54.480 42.480 54.820 42.770 ;
        RECT 81.440 42.480 81.780 42.770 ;
        RECT 82.760 42.480 83.100 42.770 ;
        RECT 84.080 42.480 84.420 42.770 ;
        RECT 85.400 42.480 85.740 42.770 ;
        RECT 97.280 42.480 97.620 42.770 ;
        RECT 98.600 42.480 98.940 42.770 ;
        RECT 99.920 42.480 100.260 42.770 ;
        RECT 101.240 42.480 101.580 42.770 ;
        RECT 102.560 42.480 102.900 42.770 ;
        RECT 103.880 42.480 104.220 42.770 ;
        RECT 105.200 42.480 105.540 42.770 ;
        RECT 106.520 42.480 106.860 42.770 ;
        RECT 118.400 42.480 118.740 42.770 ;
        RECT 119.720 42.480 120.060 42.770 ;
        RECT 121.040 42.480 121.380 42.770 ;
        RECT 122.360 42.480 122.700 42.770 ;
        RECT 13.240 42.140 55.440 42.480 ;
        RECT 55.780 42.140 57.040 42.480 ;
        RECT 79.220 42.140 80.480 42.480 ;
        RECT 80.820 42.140 123.020 42.480 ;
        RECT 13.560 41.850 13.900 42.140 ;
        RECT 14.880 41.850 15.220 42.140 ;
        RECT 16.200 41.850 16.540 42.140 ;
        RECT 17.520 41.850 17.860 42.140 ;
        RECT 29.400 41.850 29.740 42.140 ;
        RECT 30.720 41.850 31.060 42.140 ;
        RECT 32.040 41.850 32.380 42.140 ;
        RECT 33.360 41.850 33.700 42.140 ;
        RECT 34.680 41.850 35.020 42.140 ;
        RECT 36.000 41.850 36.340 42.140 ;
        RECT 37.320 41.850 37.660 42.140 ;
        RECT 38.640 41.850 38.980 42.140 ;
        RECT 50.520 41.850 50.860 42.140 ;
        RECT 51.840 41.850 52.180 42.140 ;
        RECT 53.160 41.850 53.500 42.140 ;
        RECT 54.480 41.850 54.820 42.140 ;
        RECT 81.440 41.850 81.780 42.140 ;
        RECT 82.760 41.850 83.100 42.140 ;
        RECT 84.080 41.850 84.420 42.140 ;
        RECT 85.400 41.850 85.740 42.140 ;
        RECT 97.280 41.850 97.620 42.140 ;
        RECT 98.600 41.850 98.940 42.140 ;
        RECT 99.920 41.850 100.260 42.140 ;
        RECT 101.240 41.850 101.580 42.140 ;
        RECT 102.560 41.850 102.900 42.140 ;
        RECT 103.880 41.850 104.220 42.140 ;
        RECT 105.200 41.850 105.540 42.140 ;
        RECT 106.520 41.850 106.860 42.140 ;
        RECT 118.400 41.850 118.740 42.140 ;
        RECT 119.720 41.850 120.060 42.140 ;
        RECT 121.040 41.850 121.380 42.140 ;
        RECT 122.360 41.850 122.700 42.140 ;
        RECT 45.240 39.460 45.580 39.750 ;
        RECT 90.680 39.460 91.020 39.750 ;
        RECT 13.240 39.120 55.440 39.460 ;
        RECT 55.780 39.120 57.040 39.460 ;
        RECT 79.220 39.120 80.480 39.460 ;
        RECT 80.820 39.120 123.020 39.460 ;
        RECT 45.240 38.830 45.580 39.120 ;
        RECT 90.680 38.830 91.020 39.120 ;
        RECT 11.070 36.240 46.710 36.640 ;
        RECT 11.070 35.440 45.990 35.840 ;
        RECT 11.070 34.240 11.430 35.440 ;
        RECT 46.350 35.040 46.710 36.240 ;
        RECT 11.790 34.640 46.710 35.040 ;
        RECT 11.070 33.840 45.990 34.240 ;
        RECT 11.070 32.640 11.430 33.840 ;
        RECT 46.350 33.440 46.710 34.640 ;
        RECT 11.790 33.040 46.710 33.440 ;
        RECT 89.550 36.240 125.190 36.640 ;
        RECT 89.550 35.040 89.910 36.240 ;
        RECT 90.270 35.440 125.190 35.840 ;
        RECT 89.550 34.640 124.470 35.040 ;
        RECT 89.550 33.440 89.910 34.640 ;
        RECT 124.830 34.240 125.190 35.440 ;
        RECT 90.270 33.840 125.190 34.240 ;
        RECT 89.550 33.040 124.470 33.440 ;
        RECT 124.830 32.640 125.190 33.840 ;
        RECT 11.070 32.240 46.710 32.640 ;
        RECT 89.550 32.240 125.190 32.640 ;
        RECT 11.070 31.440 46.710 31.840 ;
        RECT 11.070 30.640 45.990 31.040 ;
        RECT 11.070 29.440 11.430 30.640 ;
        RECT 46.350 30.240 46.710 31.440 ;
        RECT 11.790 29.840 46.710 30.240 ;
        RECT 89.550 31.440 125.190 31.840 ;
        RECT 89.550 30.240 89.910 31.440 ;
        RECT 90.270 30.640 125.190 31.040 ;
        RECT 11.070 29.040 45.990 29.440 ;
        RECT 11.070 27.840 11.430 29.040 ;
        RECT 46.350 28.640 46.710 29.840 ;
        RECT 11.790 28.240 46.710 28.640 ;
        RECT 47.790 29.250 48.870 30.180 ;
        RECT 51.470 29.350 53.190 29.690 ;
        RECT 56.070 29.350 57.930 29.690 ;
        RECT 51.470 29.250 51.810 29.350 ;
        RECT 47.790 28.910 51.810 29.250 ;
        RECT 11.070 27.440 46.710 27.840 ;
        RECT 11.070 26.640 46.710 27.040 ;
        RECT 11.070 25.840 45.990 26.240 ;
        RECT 11.070 24.640 11.430 25.840 ;
        RECT 46.350 25.440 46.710 26.640 ;
        RECT 11.790 25.040 46.710 25.440 ;
        RECT 11.070 24.240 45.990 24.640 ;
        RECT 11.070 23.040 11.430 24.240 ;
        RECT 46.350 23.840 46.710 25.040 ;
        RECT 11.790 23.440 46.710 23.840 ;
        RECT 47.790 25.730 48.870 28.910 ;
        RECT 51.470 28.810 51.810 28.910 ;
        RECT 57.590 29.250 57.930 29.350 ;
        RECT 60.390 29.250 61.470 30.180 ;
        RECT 57.590 29.200 61.470 29.250 ;
        RECT 74.790 29.250 75.870 30.180 ;
        RECT 78.330 29.350 80.190 29.690 ;
        RECT 83.070 29.350 84.790 29.690 ;
        RECT 78.330 29.250 78.670 29.350 ;
        RECT 74.790 29.200 78.670 29.250 ;
        RECT 57.590 28.910 67.290 29.200 ;
        RECT 57.590 28.810 57.930 28.910 ;
        RECT 51.470 28.470 53.190 28.810 ;
        RECT 56.070 28.470 57.930 28.810 ;
        RECT 60.390 28.860 67.290 28.910 ;
        RECT 51.470 27.590 53.190 27.930 ;
        RECT 56.070 27.590 57.150 27.930 ;
        RECT 51.470 27.490 51.810 27.590 ;
        RECT 49.950 27.150 51.810 27.490 ;
        RECT 58.230 27.150 59.310 27.490 ;
        RECT 52.110 26.710 53.190 27.050 ;
        RECT 56.070 26.710 57.150 27.050 ;
        RECT 51.470 25.830 53.190 26.170 ;
        RECT 56.070 25.830 57.930 26.170 ;
        RECT 51.470 25.730 51.810 25.830 ;
        RECT 47.790 25.390 51.810 25.730 ;
        RECT 11.070 22.640 46.710 23.040 ;
        RECT 11.070 21.840 46.710 22.240 ;
        RECT 11.070 21.040 45.990 21.440 ;
        RECT 11.070 19.840 11.430 21.040 ;
        RECT 46.350 20.640 46.710 21.840 ;
        RECT 11.790 20.240 46.710 20.640 ;
        RECT 11.070 19.440 45.990 19.840 ;
        RECT 11.070 18.240 11.430 19.440 ;
        RECT 46.350 19.040 46.710 20.240 ;
        RECT 11.790 18.640 46.710 19.040 ;
        RECT 11.070 17.840 46.710 18.240 ;
        RECT 11.070 17.040 46.710 17.440 ;
        RECT 11.070 16.240 45.990 16.640 ;
        RECT 11.070 15.040 11.430 16.240 ;
        RECT 46.350 15.840 46.710 17.040 ;
        RECT 11.790 15.440 46.710 15.840 ;
        RECT 11.070 14.640 45.990 15.040 ;
        RECT 11.070 13.440 11.430 14.640 ;
        RECT 46.350 14.240 46.710 15.440 ;
        RECT 11.790 13.840 46.710 14.240 ;
        RECT 47.790 14.290 48.870 25.390 ;
        RECT 51.470 25.290 51.810 25.390 ;
        RECT 57.590 25.730 57.930 25.830 ;
        RECT 60.390 25.730 61.470 28.860 ;
        RECT 63.270 26.710 64.990 27.050 ;
        RECT 57.590 25.390 61.470 25.730 ;
        RECT 57.590 25.290 57.930 25.390 ;
        RECT 51.470 24.950 53.190 25.290 ;
        RECT 56.070 24.950 57.930 25.290 ;
        RECT 52.270 24.410 53.190 24.580 ;
        RECT 52.110 24.070 53.190 24.410 ;
        RECT 56.070 24.070 57.930 24.410 ;
        RECT 57.590 23.970 57.930 24.070 ;
        RECT 49.950 23.630 51.030 23.970 ;
        RECT 57.590 23.630 59.310 23.970 ;
        RECT 52.110 23.190 53.190 23.530 ;
        RECT 56.070 23.190 57.150 23.530 ;
        RECT 52.110 22.310 53.190 22.650 ;
        RECT 55.430 22.310 57.150 22.650 ;
        RECT 49.950 21.870 51.810 22.210 ;
        RECT 49.950 20.990 51.030 21.330 ;
        RECT 51.470 20.890 51.810 21.870 ;
        RECT 52.110 21.430 53.190 21.770 ;
        RECT 55.430 20.890 55.770 22.310 ;
        RECT 58.230 21.870 59.310 22.210 ;
        RECT 56.070 21.430 57.150 21.770 ;
        RECT 58.230 20.990 59.310 21.330 ;
        RECT 51.470 20.550 55.770 20.890 ;
        RECT 56.070 20.550 57.150 20.890 ;
        RECT 52.110 19.670 57.150 20.010 ;
        RECT 49.310 19.230 51.030 19.570 ;
        RECT 57.590 19.230 59.310 19.570 ;
        RECT 49.310 17.810 49.650 19.230 ;
        RECT 52.110 18.790 57.150 19.130 ;
        RECT 49.950 18.350 51.030 18.690 ;
        RECT 52.110 17.910 53.190 18.250 ;
        RECT 56.070 17.910 57.150 18.250 ;
        RECT 49.310 17.470 51.030 17.810 ;
        RECT 57.590 17.370 57.930 19.230 ;
        RECT 58.230 18.350 59.310 18.690 ;
        RECT 58.600 17.810 58.940 18.350 ;
        RECT 58.230 17.470 59.310 17.810 ;
        RECT 52.110 17.030 57.930 17.370 ;
        RECT 56.230 16.490 57.150 16.660 ;
        RECT 52.110 16.150 57.150 16.490 ;
        RECT 49.950 15.710 51.030 16.050 ;
        RECT 58.230 15.710 59.310 16.050 ;
        RECT 52.110 15.270 53.190 15.610 ;
        RECT 56.070 15.270 57.150 15.610 ;
        RECT 51.470 14.390 53.190 14.730 ;
        RECT 56.070 14.390 57.930 14.730 ;
        RECT 51.470 14.290 51.810 14.390 ;
        RECT 47.790 13.950 51.810 14.290 ;
        RECT 11.070 13.040 46.710 13.440 ;
        RECT 47.790 13.020 48.870 13.950 ;
        RECT 51.470 13.850 51.810 13.950 ;
        RECT 57.590 14.290 57.930 14.390 ;
        RECT 60.390 14.290 61.470 25.390 ;
        RECT 62.630 25.830 64.350 26.170 ;
        RECT 62.630 24.410 62.970 25.830 ;
        RECT 64.650 25.290 64.990 26.710 ;
        RECT 65.430 26.270 66.510 26.610 ;
        RECT 66.950 26.560 67.290 28.860 ;
        RECT 68.970 28.910 78.670 29.200 ;
        RECT 68.970 28.860 75.870 28.910 ;
        RECT 67.590 26.560 68.670 27.540 ;
        RECT 68.970 26.560 69.310 28.860 ;
        RECT 71.270 26.710 72.990 27.050 ;
        RECT 63.270 24.950 64.990 25.290 ;
        RECT 62.630 24.070 64.350 24.410 ;
        RECT 62.630 22.650 62.970 24.070 ;
        RECT 64.650 23.530 64.990 24.950 ;
        RECT 65.800 24.850 66.140 26.270 ;
        RECT 66.950 26.220 69.310 26.560 ;
        RECT 69.750 26.270 70.830 26.610 ;
        RECT 65.430 24.510 66.510 24.850 ;
        RECT 63.270 23.190 64.990 23.530 ;
        RECT 62.630 22.310 64.350 22.650 ;
        RECT 62.630 20.890 62.970 22.310 ;
        RECT 64.650 21.770 64.990 23.190 ;
        RECT 65.800 23.090 66.140 24.510 ;
        RECT 65.430 22.750 66.510 23.090 ;
        RECT 63.270 21.430 64.990 21.770 ;
        RECT 62.630 20.550 64.350 20.890 ;
        RECT 64.650 20.010 64.990 21.430 ;
        RECT 65.800 21.330 66.140 22.750 ;
        RECT 65.430 20.990 66.510 21.330 ;
        RECT 63.270 19.670 64.990 20.010 ;
        RECT 57.590 13.950 61.470 14.290 ;
        RECT 57.590 13.850 57.930 13.950 ;
        RECT 51.470 13.510 53.190 13.850 ;
        RECT 56.070 13.510 57.930 13.850 ;
        RECT 60.390 13.020 61.470 13.950 ;
        RECT 62.630 18.790 64.350 19.130 ;
        RECT 62.630 17.370 62.970 18.790 ;
        RECT 64.650 18.250 64.990 19.670 ;
        RECT 65.430 19.230 66.510 19.570 ;
        RECT 63.270 17.910 64.990 18.250 ;
        RECT 62.630 17.030 64.350 17.370 ;
        RECT 62.630 15.610 62.970 17.030 ;
        RECT 64.650 16.490 64.990 17.910 ;
        RECT 65.800 17.810 66.140 19.230 ;
        RECT 65.430 17.470 66.510 17.810 ;
        RECT 63.270 16.150 64.990 16.490 ;
        RECT 62.630 15.270 64.350 15.610 ;
        RECT 62.630 13.850 62.970 15.270 ;
        RECT 64.650 14.730 64.990 16.150 ;
        RECT 65.800 16.050 66.140 17.470 ;
        RECT 65.430 15.710 66.510 16.050 ;
        RECT 63.270 14.390 64.990 14.730 ;
        RECT 65.800 14.290 66.140 15.710 ;
        RECT 65.430 13.950 66.510 14.290 ;
        RECT 62.630 13.510 64.350 13.850 ;
        RECT 67.590 13.020 68.670 26.220 ;
        RECT 70.120 24.850 70.460 26.270 ;
        RECT 71.270 25.290 71.610 26.710 ;
        RECT 71.910 25.830 73.630 26.170 ;
        RECT 71.270 24.950 72.990 25.290 ;
        RECT 69.750 24.510 70.830 24.850 ;
        RECT 70.120 23.090 70.460 24.510 ;
        RECT 71.270 23.530 71.610 24.950 ;
        RECT 73.290 24.410 73.630 25.830 ;
        RECT 71.910 24.070 73.630 24.410 ;
        RECT 71.270 23.190 72.990 23.530 ;
        RECT 69.750 22.750 70.830 23.090 ;
        RECT 70.120 21.330 70.460 22.750 ;
        RECT 71.270 21.770 71.610 23.190 ;
        RECT 73.290 22.650 73.630 24.070 ;
        RECT 71.910 22.310 73.630 22.650 ;
        RECT 71.270 21.430 72.990 21.770 ;
        RECT 69.750 20.990 70.830 21.330 ;
        RECT 71.270 20.010 71.610 21.430 ;
        RECT 73.290 20.890 73.630 22.310 ;
        RECT 71.910 20.550 73.630 20.890 ;
        RECT 74.790 25.730 75.870 28.860 ;
        RECT 78.330 28.810 78.670 28.910 ;
        RECT 84.450 29.250 84.790 29.350 ;
        RECT 87.390 29.250 88.470 30.180 ;
        RECT 84.450 28.910 88.470 29.250 ;
        RECT 84.450 28.810 84.790 28.910 ;
        RECT 78.330 28.470 80.190 28.810 ;
        RECT 83.070 28.470 84.790 28.810 ;
        RECT 79.110 27.590 80.190 27.930 ;
        RECT 83.070 27.590 84.790 27.930 ;
        RECT 84.450 27.490 84.790 27.590 ;
        RECT 76.950 27.150 78.030 27.490 ;
        RECT 84.450 27.150 86.310 27.490 ;
        RECT 79.110 26.710 80.190 27.050 ;
        RECT 83.070 26.710 84.150 27.050 ;
        RECT 78.330 25.830 80.190 26.170 ;
        RECT 83.070 25.830 84.790 26.170 ;
        RECT 78.330 25.730 78.670 25.830 ;
        RECT 74.790 25.390 78.670 25.730 ;
        RECT 71.270 19.670 72.990 20.010 ;
        RECT 69.750 19.230 70.830 19.570 ;
        RECT 70.120 17.810 70.460 19.230 ;
        RECT 71.270 18.250 71.610 19.670 ;
        RECT 71.910 18.790 73.630 19.130 ;
        RECT 71.270 17.910 72.990 18.250 ;
        RECT 69.750 17.470 70.830 17.810 ;
        RECT 70.120 16.050 70.460 17.470 ;
        RECT 71.270 16.490 71.610 17.910 ;
        RECT 73.290 17.370 73.630 18.790 ;
        RECT 71.910 17.030 73.630 17.370 ;
        RECT 71.270 16.150 72.990 16.490 ;
        RECT 69.750 15.710 70.830 16.050 ;
        RECT 70.120 14.290 70.460 15.710 ;
        RECT 71.270 14.730 71.610 16.150 ;
        RECT 73.290 15.610 73.630 17.030 ;
        RECT 71.910 15.270 73.630 15.610 ;
        RECT 71.270 14.390 72.990 14.730 ;
        RECT 69.750 13.950 70.830 14.290 ;
        RECT 73.290 13.850 73.630 15.270 ;
        RECT 71.910 13.510 73.630 13.850 ;
        RECT 74.790 14.290 75.870 25.390 ;
        RECT 78.330 25.290 78.670 25.390 ;
        RECT 84.450 25.730 84.790 25.830 ;
        RECT 87.390 25.730 88.470 28.910 ;
        RECT 89.550 29.840 124.470 30.240 ;
        RECT 89.550 28.640 89.910 29.840 ;
        RECT 124.830 29.440 125.190 30.640 ;
        RECT 90.270 29.040 125.190 29.440 ;
        RECT 89.550 28.240 124.470 28.640 ;
        RECT 124.830 27.840 125.190 29.040 ;
        RECT 89.550 27.440 125.190 27.840 ;
        RECT 84.450 25.390 88.470 25.730 ;
        RECT 84.450 25.290 84.790 25.390 ;
        RECT 78.330 24.950 80.190 25.290 ;
        RECT 83.070 24.950 84.790 25.290 ;
        RECT 83.070 24.410 83.990 24.580 ;
        RECT 78.330 24.070 80.190 24.410 ;
        RECT 83.070 24.070 84.150 24.410 ;
        RECT 78.330 23.970 78.670 24.070 ;
        RECT 76.950 23.630 78.670 23.970 ;
        RECT 85.230 23.630 86.310 23.970 ;
        RECT 79.110 23.190 80.190 23.530 ;
        RECT 83.070 23.190 84.150 23.530 ;
        RECT 79.110 22.310 80.830 22.650 ;
        RECT 83.070 22.310 84.150 22.650 ;
        RECT 76.950 21.870 78.030 22.210 ;
        RECT 79.110 21.430 80.190 21.770 ;
        RECT 76.950 20.990 78.030 21.330 ;
        RECT 80.490 20.890 80.830 22.310 ;
        RECT 84.450 21.870 86.310 22.210 ;
        RECT 83.070 21.430 84.150 21.770 ;
        RECT 84.450 20.890 84.790 21.870 ;
        RECT 85.230 20.990 86.310 21.330 ;
        RECT 79.110 20.550 80.190 20.890 ;
        RECT 80.490 20.550 84.790 20.890 ;
        RECT 79.110 19.670 84.150 20.010 ;
        RECT 76.950 19.230 78.670 19.570 ;
        RECT 85.230 19.230 86.950 19.570 ;
        RECT 76.950 18.350 78.030 18.690 ;
        RECT 77.320 17.810 77.660 18.350 ;
        RECT 76.950 17.470 78.030 17.810 ;
        RECT 78.330 17.370 78.670 19.230 ;
        RECT 79.110 18.790 84.150 19.130 ;
        RECT 85.230 18.350 86.310 18.690 ;
        RECT 79.110 17.910 80.190 18.250 ;
        RECT 83.070 17.910 84.150 18.250 ;
        RECT 86.610 17.810 86.950 19.230 ;
        RECT 85.230 17.470 86.950 17.810 ;
        RECT 78.330 17.030 84.150 17.370 ;
        RECT 79.110 16.490 80.030 16.660 ;
        RECT 79.110 16.150 84.150 16.490 ;
        RECT 76.950 15.710 78.030 16.050 ;
        RECT 85.230 15.710 86.310 16.050 ;
        RECT 79.110 15.270 80.190 15.610 ;
        RECT 83.070 15.270 84.150 15.610 ;
        RECT 78.330 14.390 80.190 14.730 ;
        RECT 83.070 14.390 84.790 14.730 ;
        RECT 78.330 14.290 78.670 14.390 ;
        RECT 74.790 13.950 78.670 14.290 ;
        RECT 74.790 13.020 75.870 13.950 ;
        RECT 78.330 13.850 78.670 13.950 ;
        RECT 84.450 14.290 84.790 14.390 ;
        RECT 87.390 14.290 88.470 25.390 ;
        RECT 89.550 26.640 125.190 27.040 ;
        RECT 89.550 25.440 89.910 26.640 ;
        RECT 90.270 25.840 125.190 26.240 ;
        RECT 89.550 25.040 124.470 25.440 ;
        RECT 89.550 23.840 89.910 25.040 ;
        RECT 124.830 24.640 125.190 25.840 ;
        RECT 90.270 24.240 125.190 24.640 ;
        RECT 89.550 23.440 124.470 23.840 ;
        RECT 124.830 23.040 125.190 24.240 ;
        RECT 89.550 22.640 125.190 23.040 ;
        RECT 89.550 21.840 125.190 22.240 ;
        RECT 89.550 20.640 89.910 21.840 ;
        RECT 90.270 21.040 125.190 21.440 ;
        RECT 89.550 20.240 124.470 20.640 ;
        RECT 89.550 19.040 89.910 20.240 ;
        RECT 124.830 19.840 125.190 21.040 ;
        RECT 90.270 19.440 125.190 19.840 ;
        RECT 89.550 18.640 124.470 19.040 ;
        RECT 124.830 18.240 125.190 19.440 ;
        RECT 89.550 17.840 125.190 18.240 ;
        RECT 84.450 13.950 88.470 14.290 ;
        RECT 84.450 13.850 84.790 13.950 ;
        RECT 78.330 13.510 80.190 13.850 ;
        RECT 83.070 13.510 84.790 13.850 ;
        RECT 87.390 13.020 88.470 13.950 ;
        RECT 89.550 17.040 125.190 17.440 ;
        RECT 89.550 15.840 89.910 17.040 ;
        RECT 90.270 16.240 125.190 16.640 ;
        RECT 89.550 15.440 124.470 15.840 ;
        RECT 89.550 14.240 89.910 15.440 ;
        RECT 124.830 15.040 125.190 16.240 ;
        RECT 90.270 14.640 125.190 15.040 ;
        RECT 89.550 13.840 124.470 14.240 ;
        RECT 124.830 13.440 125.190 14.640 ;
        RECT 89.550 13.040 125.190 13.440 ;
        RECT 128.050 10.560 128.970 190.430 ;
        RECT 7.290 9.640 128.970 10.560 ;
        RECT 131.650 6.960 132.570 194.030 ;
        RECT 3.690 6.040 132.570 6.960 ;
        RECT 133.290 5.320 133.630 219.770 ;
        RECT 135.210 208.085 146.850 208.385 ;
        RECT 135.715 206.175 136.795 207.125 ;
        RECT 140.035 206.615 140.955 206.655 ;
        RECT 143.995 206.615 144.915 206.655 ;
        RECT 139.255 206.315 141.115 206.615 ;
        RECT 143.995 206.315 145.675 206.615 ;
        RECT 139.255 206.175 139.555 206.315 ;
        RECT 135.715 205.875 139.555 206.175 ;
        RECT 135.715 199.645 136.795 205.875 ;
        RECT 139.255 205.735 139.555 205.875 ;
        RECT 145.375 206.175 145.675 206.315 ;
        RECT 148.315 206.175 149.395 207.125 ;
        RECT 145.375 205.875 149.395 206.175 ;
        RECT 140.035 205.735 140.955 205.775 ;
        RECT 143.995 205.735 144.915 205.775 ;
        RECT 145.375 205.735 145.675 205.875 ;
        RECT 139.255 205.435 141.115 205.735 ;
        RECT 143.995 205.435 145.675 205.735 ;
        RECT 144.155 204.855 145.075 204.895 ;
        RECT 139.255 204.555 141.115 204.855 ;
        RECT 143.995 204.555 145.075 204.855 ;
        RECT 139.255 204.415 139.555 204.555 ;
        RECT 137.875 204.115 139.555 204.415 ;
        RECT 146.155 204.115 147.235 204.415 ;
        RECT 140.035 203.975 140.955 204.015 ;
        RECT 143.995 203.975 144.915 204.015 ;
        RECT 140.035 203.675 141.115 203.975 ;
        RECT 143.995 203.675 145.075 203.975 ;
        RECT 140.195 203.095 141.115 203.135 ;
        RECT 140.035 202.795 145.075 203.095 ;
        RECT 137.875 202.355 139.555 202.655 ;
        RECT 146.155 202.355 147.235 202.655 ;
        RECT 138.035 200.895 138.955 200.935 ;
        RECT 137.875 200.595 138.955 200.895 ;
        RECT 139.255 200.455 139.555 202.355 ;
        RECT 140.035 202.215 140.955 202.255 ;
        RECT 143.995 202.215 144.915 202.255 ;
        RECT 140.035 201.915 141.115 202.215 ;
        RECT 143.995 201.915 145.075 202.215 ;
        RECT 140.035 201.335 140.955 201.375 ;
        RECT 143.995 201.335 144.915 201.375 ;
        RECT 140.035 201.035 141.115 201.335 ;
        RECT 143.995 201.035 145.075 201.335 ;
        RECT 146.155 200.595 147.235 200.895 ;
        RECT 139.255 200.155 145.075 200.455 ;
        RECT 148.315 199.645 149.395 205.875 ;
        RECT 3.690 4.980 133.630 5.320 ;
        RECT 2.630 3.920 133.630 4.260 ;
      LAYER mcon ;
        RECT 60.150 224.050 60.390 224.290 ;
        RECT 136.440 224.020 136.740 224.320 ;
        RECT 112.670 223.050 112.910 223.290 ;
        RECT 135.210 223.020 135.510 223.320 ;
        RECT 15.450 220.350 15.730 220.630 ;
        RECT 15.970 220.350 16.250 220.630 ;
        RECT 19.330 220.350 19.610 220.630 ;
        RECT 19.850 220.350 20.130 220.630 ;
        RECT 15.370 219.470 15.650 219.750 ;
        RECT 15.890 219.470 16.170 219.750 ;
        RECT 19.330 219.470 19.610 219.750 ;
        RECT 19.850 219.470 20.130 219.750 ;
        RECT 13.210 218.150 13.490 218.430 ;
        RECT 13.730 218.150 14.010 218.430 ;
        RECT 15.370 216.830 15.650 217.110 ;
        RECT 15.890 216.830 16.170 217.110 ;
        RECT 19.330 216.830 19.610 217.110 ;
        RECT 19.850 216.830 20.130 217.110 ;
        RECT 13.210 212.870 13.490 213.150 ;
        RECT 13.730 212.870 14.010 213.150 ;
        RECT 15.370 214.190 15.650 214.470 ;
        RECT 15.890 214.190 16.170 214.470 ;
        RECT 19.330 214.190 19.610 214.470 ;
        RECT 19.850 214.190 20.130 214.470 ;
        RECT 19.330 213.310 19.610 213.590 ;
        RECT 19.850 213.310 20.130 213.590 ;
        RECT 15.370 212.430 15.650 212.710 ;
        RECT 15.890 212.430 16.170 212.710 ;
        RECT 19.330 212.430 19.610 212.710 ;
        RECT 19.850 212.430 20.130 212.710 ;
        RECT 15.370 211.550 15.650 211.830 ;
        RECT 15.890 211.550 16.170 211.830 ;
        RECT 13.210 208.470 13.490 208.750 ;
        RECT 13.730 208.470 14.010 208.750 ;
        RECT 13.290 207.590 13.570 207.870 ;
        RECT 13.810 207.590 14.090 207.870 ;
        RECT 15.370 209.790 15.650 210.070 ;
        RECT 15.890 209.790 16.170 210.070 ;
        RECT 19.330 209.790 19.610 210.070 ;
        RECT 19.850 209.790 20.130 210.070 ;
        RECT 21.490 217.270 21.770 217.550 ;
        RECT 22.010 217.270 22.290 217.550 ;
        RECT 21.490 215.510 21.770 215.790 ;
        RECT 22.010 215.510 22.290 215.790 ;
        RECT 21.490 214.630 21.770 214.910 ;
        RECT 22.010 214.630 22.290 214.910 ;
        RECT 21.490 211.110 21.770 211.390 ;
        RECT 22.010 211.110 22.290 211.390 ;
        RECT 21.490 210.230 21.770 210.510 ;
        RECT 22.010 210.230 22.290 210.510 ;
        RECT 15.370 207.150 15.650 207.430 ;
        RECT 15.890 207.150 16.170 207.430 ;
        RECT 19.330 207.150 19.610 207.430 ;
        RECT 19.850 207.150 20.130 207.430 ;
        RECT 15.370 205.390 15.650 205.670 ;
        RECT 15.890 205.390 16.170 205.670 ;
        RECT 19.330 205.390 19.610 205.670 ;
        RECT 19.850 205.390 20.130 205.670 ;
        RECT 15.370 204.510 15.650 204.790 ;
        RECT 15.890 204.510 16.170 204.790 ;
        RECT 19.330 204.510 19.610 204.790 ;
        RECT 19.850 204.510 20.130 204.790 ;
        RECT 13.290 204.070 13.570 204.350 ;
        RECT 13.810 204.070 14.090 204.350 ;
        RECT 15.370 203.630 15.650 203.910 ;
        RECT 15.890 203.630 16.170 203.910 ;
        RECT 19.330 203.630 19.610 203.910 ;
        RECT 19.850 203.630 20.130 203.910 ;
        RECT 15.370 202.750 15.650 203.030 ;
        RECT 15.890 202.750 16.170 203.030 ;
        RECT 19.330 202.750 19.610 203.030 ;
        RECT 19.850 202.750 20.130 203.030 ;
        RECT 28.130 220.350 28.410 220.630 ;
        RECT 28.650 220.350 28.930 220.630 ;
        RECT 32.010 220.350 32.290 220.630 ;
        RECT 32.530 220.350 32.810 220.630 ;
        RECT 28.130 219.470 28.410 219.750 ;
        RECT 28.650 219.470 28.930 219.750 ;
        RECT 32.090 219.470 32.370 219.750 ;
        RECT 32.610 219.470 32.890 219.750 ;
        RECT 25.970 217.270 26.250 217.550 ;
        RECT 26.490 217.270 26.770 217.550 ;
        RECT 25.970 215.510 26.250 215.790 ;
        RECT 26.490 215.510 26.770 215.790 ;
        RECT 25.970 214.630 26.250 214.910 ;
        RECT 26.490 214.630 26.770 214.910 ;
        RECT 25.970 211.110 26.250 211.390 ;
        RECT 26.490 211.110 26.770 211.390 ;
        RECT 25.970 210.230 26.250 210.510 ;
        RECT 26.490 210.230 26.770 210.510 ;
        RECT 28.130 216.830 28.410 217.110 ;
        RECT 28.650 216.830 28.930 217.110 ;
        RECT 34.250 218.150 34.530 218.430 ;
        RECT 34.770 218.150 35.050 218.430 ;
        RECT 32.090 216.830 32.370 217.110 ;
        RECT 32.610 216.830 32.890 217.110 ;
        RECT 28.130 214.190 28.410 214.470 ;
        RECT 28.650 214.190 28.930 214.470 ;
        RECT 32.090 214.190 32.370 214.470 ;
        RECT 32.610 214.190 32.890 214.470 ;
        RECT 28.130 213.310 28.410 213.590 ;
        RECT 28.650 213.310 28.930 213.590 ;
        RECT 28.130 212.430 28.410 212.710 ;
        RECT 28.650 212.430 28.930 212.710 ;
        RECT 32.090 212.430 32.370 212.710 ;
        RECT 32.610 212.430 32.890 212.710 ;
        RECT 32.090 211.550 32.370 211.830 ;
        RECT 32.610 211.550 32.890 211.830 ;
        RECT 28.130 209.790 28.410 210.070 ;
        RECT 28.650 209.790 28.930 210.070 ;
        RECT 34.250 212.870 34.530 213.150 ;
        RECT 34.770 212.870 35.050 213.150 ;
        RECT 32.090 209.790 32.370 210.070 ;
        RECT 32.610 209.790 32.890 210.070 ;
        RECT 28.130 207.150 28.410 207.430 ;
        RECT 28.650 207.150 28.930 207.430 ;
        RECT 32.090 207.150 32.370 207.430 ;
        RECT 32.610 207.150 32.890 207.430 ;
        RECT 34.250 208.470 34.530 208.750 ;
        RECT 34.770 208.470 35.050 208.750 ;
        RECT 34.170 207.590 34.450 207.870 ;
        RECT 34.690 207.590 34.970 207.870 ;
        RECT 28.130 205.390 28.410 205.670 ;
        RECT 28.650 205.390 28.930 205.670 ;
        RECT 32.090 205.390 32.370 205.670 ;
        RECT 32.610 205.390 32.890 205.670 ;
        RECT 28.130 204.510 28.410 204.790 ;
        RECT 28.650 204.510 28.930 204.790 ;
        RECT 32.090 204.510 32.370 204.790 ;
        RECT 32.610 204.510 32.890 204.790 ;
        RECT 34.170 204.070 34.450 204.350 ;
        RECT 34.690 204.070 34.970 204.350 ;
        RECT 28.130 203.630 28.410 203.910 ;
        RECT 28.650 203.630 28.930 203.910 ;
        RECT 32.090 203.630 32.370 203.910 ;
        RECT 32.610 203.630 32.890 203.910 ;
        RECT 28.130 202.750 28.410 203.030 ;
        RECT 28.650 202.750 28.930 203.030 ;
        RECT 32.090 202.750 32.370 203.030 ;
        RECT 32.610 202.750 32.890 203.030 ;
        RECT 15.370 201.870 15.650 202.150 ;
        RECT 15.890 201.870 16.170 202.150 ;
        RECT 19.330 201.870 19.610 202.150 ;
        RECT 19.850 201.870 20.130 202.150 ;
        RECT 40.650 220.350 40.930 220.630 ;
        RECT 41.170 220.350 41.450 220.630 ;
        RECT 44.530 220.350 44.810 220.630 ;
        RECT 45.050 220.350 45.330 220.630 ;
        RECT 40.570 219.470 40.850 219.750 ;
        RECT 41.090 219.470 41.370 219.750 ;
        RECT 44.530 219.470 44.810 219.750 ;
        RECT 45.050 219.470 45.330 219.750 ;
        RECT 38.410 218.150 38.690 218.430 ;
        RECT 38.930 218.150 39.210 218.430 ;
        RECT 40.570 216.830 40.850 217.110 ;
        RECT 41.090 216.830 41.370 217.110 ;
        RECT 44.530 216.830 44.810 217.110 ;
        RECT 45.050 216.830 45.330 217.110 ;
        RECT 38.410 212.870 38.690 213.150 ;
        RECT 38.930 212.870 39.210 213.150 ;
        RECT 40.570 214.190 40.850 214.470 ;
        RECT 41.090 214.190 41.370 214.470 ;
        RECT 44.530 214.190 44.810 214.470 ;
        RECT 45.050 214.190 45.330 214.470 ;
        RECT 44.530 213.310 44.810 213.590 ;
        RECT 45.050 213.310 45.330 213.590 ;
        RECT 40.570 212.430 40.850 212.710 ;
        RECT 41.090 212.430 41.370 212.710 ;
        RECT 44.530 212.430 44.810 212.710 ;
        RECT 45.050 212.430 45.330 212.710 ;
        RECT 40.570 211.550 40.850 211.830 ;
        RECT 41.090 211.550 41.370 211.830 ;
        RECT 38.410 208.470 38.690 208.750 ;
        RECT 38.930 208.470 39.210 208.750 ;
        RECT 38.490 207.590 38.770 207.870 ;
        RECT 39.010 207.590 39.290 207.870 ;
        RECT 40.570 209.790 40.850 210.070 ;
        RECT 41.090 209.790 41.370 210.070 ;
        RECT 44.530 209.790 44.810 210.070 ;
        RECT 45.050 209.790 45.330 210.070 ;
        RECT 46.690 217.270 46.970 217.550 ;
        RECT 47.210 217.270 47.490 217.550 ;
        RECT 46.690 215.510 46.970 215.790 ;
        RECT 47.210 215.510 47.490 215.790 ;
        RECT 46.690 214.630 46.970 214.910 ;
        RECT 47.210 214.630 47.490 214.910 ;
        RECT 46.690 211.110 46.970 211.390 ;
        RECT 47.210 211.110 47.490 211.390 ;
        RECT 46.690 210.230 46.970 210.510 ;
        RECT 47.210 210.230 47.490 210.510 ;
        RECT 40.570 207.150 40.850 207.430 ;
        RECT 41.090 207.150 41.370 207.430 ;
        RECT 44.530 207.150 44.810 207.430 ;
        RECT 45.050 207.150 45.330 207.430 ;
        RECT 40.570 205.390 40.850 205.670 ;
        RECT 41.090 205.390 41.370 205.670 ;
        RECT 44.530 205.390 44.810 205.670 ;
        RECT 45.050 205.390 45.330 205.670 ;
        RECT 40.570 204.510 40.850 204.790 ;
        RECT 41.090 204.510 41.370 204.790 ;
        RECT 44.530 204.510 44.810 204.790 ;
        RECT 45.050 204.510 45.330 204.790 ;
        RECT 38.490 204.070 38.770 204.350 ;
        RECT 39.010 204.070 39.290 204.350 ;
        RECT 40.570 203.630 40.850 203.910 ;
        RECT 41.090 203.630 41.370 203.910 ;
        RECT 44.530 203.630 44.810 203.910 ;
        RECT 45.050 203.630 45.330 203.910 ;
        RECT 40.570 202.750 40.850 203.030 ;
        RECT 41.090 202.750 41.370 203.030 ;
        RECT 44.530 202.750 44.810 203.030 ;
        RECT 45.050 202.750 45.330 203.030 ;
        RECT 28.130 201.870 28.410 202.150 ;
        RECT 28.650 201.870 28.930 202.150 ;
        RECT 32.090 201.870 32.370 202.150 ;
        RECT 32.610 201.870 32.890 202.150 ;
        RECT 53.330 220.350 53.610 220.630 ;
        RECT 53.850 220.350 54.130 220.630 ;
        RECT 57.210 220.350 57.490 220.630 ;
        RECT 57.730 220.350 58.010 220.630 ;
        RECT 53.330 219.470 53.610 219.750 ;
        RECT 53.850 219.470 54.130 219.750 ;
        RECT 57.290 219.470 57.570 219.750 ;
        RECT 57.810 219.470 58.090 219.750 ;
        RECT 51.170 217.270 51.450 217.550 ;
        RECT 51.690 217.270 51.970 217.550 ;
        RECT 51.170 215.510 51.450 215.790 ;
        RECT 51.690 215.510 51.970 215.790 ;
        RECT 51.170 214.630 51.450 214.910 ;
        RECT 51.690 214.630 51.970 214.910 ;
        RECT 51.170 211.110 51.450 211.390 ;
        RECT 51.690 211.110 51.970 211.390 ;
        RECT 51.170 210.230 51.450 210.510 ;
        RECT 51.690 210.230 51.970 210.510 ;
        RECT 53.330 216.830 53.610 217.110 ;
        RECT 53.850 216.830 54.130 217.110 ;
        RECT 59.450 218.150 59.730 218.430 ;
        RECT 59.970 218.150 60.250 218.430 ;
        RECT 57.290 216.830 57.570 217.110 ;
        RECT 57.810 216.830 58.090 217.110 ;
        RECT 53.330 214.190 53.610 214.470 ;
        RECT 53.850 214.190 54.130 214.470 ;
        RECT 57.290 214.190 57.570 214.470 ;
        RECT 57.810 214.190 58.090 214.470 ;
        RECT 53.330 213.310 53.610 213.590 ;
        RECT 53.850 213.310 54.130 213.590 ;
        RECT 53.330 212.430 53.610 212.710 ;
        RECT 53.850 212.430 54.130 212.710 ;
        RECT 57.290 212.430 57.570 212.710 ;
        RECT 57.810 212.430 58.090 212.710 ;
        RECT 57.290 211.550 57.570 211.830 ;
        RECT 57.810 211.550 58.090 211.830 ;
        RECT 53.330 209.790 53.610 210.070 ;
        RECT 53.850 209.790 54.130 210.070 ;
        RECT 59.450 212.870 59.730 213.150 ;
        RECT 59.970 212.870 60.250 213.150 ;
        RECT 57.290 209.790 57.570 210.070 ;
        RECT 57.810 209.790 58.090 210.070 ;
        RECT 53.330 207.150 53.610 207.430 ;
        RECT 53.850 207.150 54.130 207.430 ;
        RECT 57.290 207.150 57.570 207.430 ;
        RECT 57.810 207.150 58.090 207.430 ;
        RECT 59.450 208.470 59.730 208.750 ;
        RECT 59.970 208.470 60.250 208.750 ;
        RECT 59.370 207.590 59.650 207.870 ;
        RECT 59.890 207.590 60.170 207.870 ;
        RECT 53.330 205.390 53.610 205.670 ;
        RECT 53.850 205.390 54.130 205.670 ;
        RECT 57.290 205.390 57.570 205.670 ;
        RECT 57.810 205.390 58.090 205.670 ;
        RECT 53.330 204.510 53.610 204.790 ;
        RECT 53.850 204.510 54.130 204.790 ;
        RECT 57.290 204.510 57.570 204.790 ;
        RECT 57.810 204.510 58.090 204.790 ;
        RECT 59.370 204.070 59.650 204.350 ;
        RECT 59.890 204.070 60.170 204.350 ;
        RECT 53.330 203.630 53.610 203.910 ;
        RECT 53.850 203.630 54.130 203.910 ;
        RECT 57.290 203.630 57.570 203.910 ;
        RECT 57.810 203.630 58.090 203.910 ;
        RECT 53.330 202.750 53.610 203.030 ;
        RECT 53.850 202.750 54.130 203.030 ;
        RECT 57.290 202.750 57.570 203.030 ;
        RECT 57.810 202.750 58.090 203.030 ;
        RECT 40.570 201.870 40.850 202.150 ;
        RECT 41.090 201.870 41.370 202.150 ;
        RECT 44.530 201.870 44.810 202.150 ;
        RECT 45.050 201.870 45.330 202.150 ;
        RECT 65.850 220.350 66.130 220.630 ;
        RECT 66.370 220.350 66.650 220.630 ;
        RECT 69.730 220.350 70.010 220.630 ;
        RECT 70.250 220.350 70.530 220.630 ;
        RECT 65.770 219.470 66.050 219.750 ;
        RECT 66.290 219.470 66.570 219.750 ;
        RECT 69.730 219.470 70.010 219.750 ;
        RECT 70.250 219.470 70.530 219.750 ;
        RECT 63.610 218.150 63.890 218.430 ;
        RECT 64.130 218.150 64.410 218.430 ;
        RECT 65.770 216.830 66.050 217.110 ;
        RECT 66.290 216.830 66.570 217.110 ;
        RECT 69.730 216.830 70.010 217.110 ;
        RECT 70.250 216.830 70.530 217.110 ;
        RECT 63.610 212.870 63.890 213.150 ;
        RECT 64.130 212.870 64.410 213.150 ;
        RECT 65.770 214.190 66.050 214.470 ;
        RECT 66.290 214.190 66.570 214.470 ;
        RECT 69.730 214.190 70.010 214.470 ;
        RECT 70.250 214.190 70.530 214.470 ;
        RECT 69.730 213.310 70.010 213.590 ;
        RECT 70.250 213.310 70.530 213.590 ;
        RECT 65.770 212.430 66.050 212.710 ;
        RECT 66.290 212.430 66.570 212.710 ;
        RECT 69.730 212.430 70.010 212.710 ;
        RECT 70.250 212.430 70.530 212.710 ;
        RECT 65.770 211.550 66.050 211.830 ;
        RECT 66.290 211.550 66.570 211.830 ;
        RECT 63.610 208.470 63.890 208.750 ;
        RECT 64.130 208.470 64.410 208.750 ;
        RECT 63.690 207.590 63.970 207.870 ;
        RECT 64.210 207.590 64.490 207.870 ;
        RECT 65.770 209.790 66.050 210.070 ;
        RECT 66.290 209.790 66.570 210.070 ;
        RECT 69.730 209.790 70.010 210.070 ;
        RECT 70.250 209.790 70.530 210.070 ;
        RECT 71.890 217.270 72.170 217.550 ;
        RECT 72.410 217.270 72.690 217.550 ;
        RECT 71.890 215.510 72.170 215.790 ;
        RECT 72.410 215.510 72.690 215.790 ;
        RECT 71.890 214.630 72.170 214.910 ;
        RECT 72.410 214.630 72.690 214.910 ;
        RECT 71.890 211.110 72.170 211.390 ;
        RECT 72.410 211.110 72.690 211.390 ;
        RECT 71.890 210.230 72.170 210.510 ;
        RECT 72.410 210.230 72.690 210.510 ;
        RECT 65.770 207.150 66.050 207.430 ;
        RECT 66.290 207.150 66.570 207.430 ;
        RECT 69.730 207.150 70.010 207.430 ;
        RECT 70.250 207.150 70.530 207.430 ;
        RECT 65.770 205.390 66.050 205.670 ;
        RECT 66.290 205.390 66.570 205.670 ;
        RECT 69.730 205.390 70.010 205.670 ;
        RECT 70.250 205.390 70.530 205.670 ;
        RECT 65.770 204.510 66.050 204.790 ;
        RECT 66.290 204.510 66.570 204.790 ;
        RECT 69.730 204.510 70.010 204.790 ;
        RECT 70.250 204.510 70.530 204.790 ;
        RECT 63.690 204.070 63.970 204.350 ;
        RECT 64.210 204.070 64.490 204.350 ;
        RECT 65.770 203.630 66.050 203.910 ;
        RECT 66.290 203.630 66.570 203.910 ;
        RECT 69.730 203.630 70.010 203.910 ;
        RECT 70.250 203.630 70.530 203.910 ;
        RECT 65.770 202.750 66.050 203.030 ;
        RECT 66.290 202.750 66.570 203.030 ;
        RECT 69.730 202.750 70.010 203.030 ;
        RECT 70.250 202.750 70.530 203.030 ;
        RECT 53.330 201.870 53.610 202.150 ;
        RECT 53.850 201.870 54.130 202.150 ;
        RECT 57.290 201.870 57.570 202.150 ;
        RECT 57.810 201.870 58.090 202.150 ;
        RECT 78.530 220.350 78.810 220.630 ;
        RECT 79.050 220.350 79.330 220.630 ;
        RECT 82.410 220.350 82.690 220.630 ;
        RECT 82.930 220.350 83.210 220.630 ;
        RECT 78.530 219.470 78.810 219.750 ;
        RECT 79.050 219.470 79.330 219.750 ;
        RECT 82.490 219.470 82.770 219.750 ;
        RECT 83.010 219.470 83.290 219.750 ;
        RECT 76.370 217.270 76.650 217.550 ;
        RECT 76.890 217.270 77.170 217.550 ;
        RECT 76.370 215.510 76.650 215.790 ;
        RECT 76.890 215.510 77.170 215.790 ;
        RECT 76.370 214.630 76.650 214.910 ;
        RECT 76.890 214.630 77.170 214.910 ;
        RECT 76.370 211.110 76.650 211.390 ;
        RECT 76.890 211.110 77.170 211.390 ;
        RECT 76.370 210.230 76.650 210.510 ;
        RECT 76.890 210.230 77.170 210.510 ;
        RECT 78.530 216.830 78.810 217.110 ;
        RECT 79.050 216.830 79.330 217.110 ;
        RECT 84.650 218.150 84.930 218.430 ;
        RECT 85.170 218.150 85.450 218.430 ;
        RECT 82.490 216.830 82.770 217.110 ;
        RECT 83.010 216.830 83.290 217.110 ;
        RECT 78.530 214.190 78.810 214.470 ;
        RECT 79.050 214.190 79.330 214.470 ;
        RECT 82.490 214.190 82.770 214.470 ;
        RECT 83.010 214.190 83.290 214.470 ;
        RECT 78.530 213.310 78.810 213.590 ;
        RECT 79.050 213.310 79.330 213.590 ;
        RECT 78.530 212.430 78.810 212.710 ;
        RECT 79.050 212.430 79.330 212.710 ;
        RECT 82.490 212.430 82.770 212.710 ;
        RECT 83.010 212.430 83.290 212.710 ;
        RECT 82.490 211.550 82.770 211.830 ;
        RECT 83.010 211.550 83.290 211.830 ;
        RECT 78.530 209.790 78.810 210.070 ;
        RECT 79.050 209.790 79.330 210.070 ;
        RECT 84.650 212.870 84.930 213.150 ;
        RECT 85.170 212.870 85.450 213.150 ;
        RECT 82.490 209.790 82.770 210.070 ;
        RECT 83.010 209.790 83.290 210.070 ;
        RECT 78.530 207.150 78.810 207.430 ;
        RECT 79.050 207.150 79.330 207.430 ;
        RECT 82.490 207.150 82.770 207.430 ;
        RECT 83.010 207.150 83.290 207.430 ;
        RECT 84.650 208.470 84.930 208.750 ;
        RECT 85.170 208.470 85.450 208.750 ;
        RECT 84.570 207.590 84.850 207.870 ;
        RECT 85.090 207.590 85.370 207.870 ;
        RECT 78.530 205.390 78.810 205.670 ;
        RECT 79.050 205.390 79.330 205.670 ;
        RECT 82.490 205.390 82.770 205.670 ;
        RECT 83.010 205.390 83.290 205.670 ;
        RECT 78.530 204.510 78.810 204.790 ;
        RECT 79.050 204.510 79.330 204.790 ;
        RECT 82.490 204.510 82.770 204.790 ;
        RECT 83.010 204.510 83.290 204.790 ;
        RECT 84.570 204.070 84.850 204.350 ;
        RECT 85.090 204.070 85.370 204.350 ;
        RECT 78.530 203.630 78.810 203.910 ;
        RECT 79.050 203.630 79.330 203.910 ;
        RECT 82.490 203.630 82.770 203.910 ;
        RECT 83.010 203.630 83.290 203.910 ;
        RECT 78.530 202.750 78.810 203.030 ;
        RECT 79.050 202.750 79.330 203.030 ;
        RECT 82.490 202.750 82.770 203.030 ;
        RECT 83.010 202.750 83.290 203.030 ;
        RECT 65.770 201.870 66.050 202.150 ;
        RECT 66.290 201.870 66.570 202.150 ;
        RECT 69.730 201.870 70.010 202.150 ;
        RECT 70.250 201.870 70.530 202.150 ;
        RECT 91.050 220.350 91.330 220.630 ;
        RECT 91.570 220.350 91.850 220.630 ;
        RECT 94.930 220.350 95.210 220.630 ;
        RECT 95.450 220.350 95.730 220.630 ;
        RECT 90.970 219.470 91.250 219.750 ;
        RECT 91.490 219.470 91.770 219.750 ;
        RECT 94.930 219.470 95.210 219.750 ;
        RECT 95.450 219.470 95.730 219.750 ;
        RECT 88.810 218.150 89.090 218.430 ;
        RECT 89.330 218.150 89.610 218.430 ;
        RECT 90.970 216.830 91.250 217.110 ;
        RECT 91.490 216.830 91.770 217.110 ;
        RECT 94.930 216.830 95.210 217.110 ;
        RECT 95.450 216.830 95.730 217.110 ;
        RECT 88.810 212.870 89.090 213.150 ;
        RECT 89.330 212.870 89.610 213.150 ;
        RECT 90.970 214.190 91.250 214.470 ;
        RECT 91.490 214.190 91.770 214.470 ;
        RECT 94.930 214.190 95.210 214.470 ;
        RECT 95.450 214.190 95.730 214.470 ;
        RECT 94.930 213.310 95.210 213.590 ;
        RECT 95.450 213.310 95.730 213.590 ;
        RECT 90.970 212.430 91.250 212.710 ;
        RECT 91.490 212.430 91.770 212.710 ;
        RECT 94.930 212.430 95.210 212.710 ;
        RECT 95.450 212.430 95.730 212.710 ;
        RECT 90.970 211.550 91.250 211.830 ;
        RECT 91.490 211.550 91.770 211.830 ;
        RECT 88.810 208.470 89.090 208.750 ;
        RECT 89.330 208.470 89.610 208.750 ;
        RECT 88.890 207.590 89.170 207.870 ;
        RECT 89.410 207.590 89.690 207.870 ;
        RECT 90.970 209.790 91.250 210.070 ;
        RECT 91.490 209.790 91.770 210.070 ;
        RECT 94.930 209.790 95.210 210.070 ;
        RECT 95.450 209.790 95.730 210.070 ;
        RECT 97.090 217.270 97.370 217.550 ;
        RECT 97.610 217.270 97.890 217.550 ;
        RECT 97.090 215.510 97.370 215.790 ;
        RECT 97.610 215.510 97.890 215.790 ;
        RECT 97.090 214.630 97.370 214.910 ;
        RECT 97.610 214.630 97.890 214.910 ;
        RECT 97.090 211.110 97.370 211.390 ;
        RECT 97.610 211.110 97.890 211.390 ;
        RECT 97.090 210.230 97.370 210.510 ;
        RECT 97.610 210.230 97.890 210.510 ;
        RECT 90.970 207.150 91.250 207.430 ;
        RECT 91.490 207.150 91.770 207.430 ;
        RECT 94.930 207.150 95.210 207.430 ;
        RECT 95.450 207.150 95.730 207.430 ;
        RECT 90.970 205.390 91.250 205.670 ;
        RECT 91.490 205.390 91.770 205.670 ;
        RECT 94.930 205.390 95.210 205.670 ;
        RECT 95.450 205.390 95.730 205.670 ;
        RECT 90.970 204.510 91.250 204.790 ;
        RECT 91.490 204.510 91.770 204.790 ;
        RECT 94.930 204.510 95.210 204.790 ;
        RECT 95.450 204.510 95.730 204.790 ;
        RECT 88.890 204.070 89.170 204.350 ;
        RECT 89.410 204.070 89.690 204.350 ;
        RECT 90.970 203.630 91.250 203.910 ;
        RECT 91.490 203.630 91.770 203.910 ;
        RECT 94.930 203.630 95.210 203.910 ;
        RECT 95.450 203.630 95.730 203.910 ;
        RECT 90.970 202.750 91.250 203.030 ;
        RECT 91.490 202.750 91.770 203.030 ;
        RECT 94.930 202.750 95.210 203.030 ;
        RECT 95.450 202.750 95.730 203.030 ;
        RECT 78.530 201.870 78.810 202.150 ;
        RECT 79.050 201.870 79.330 202.150 ;
        RECT 82.490 201.870 82.770 202.150 ;
        RECT 83.010 201.870 83.290 202.150 ;
        RECT 103.730 220.350 104.010 220.630 ;
        RECT 104.250 220.350 104.530 220.630 ;
        RECT 107.610 220.350 107.890 220.630 ;
        RECT 108.130 220.350 108.410 220.630 ;
        RECT 103.730 219.470 104.010 219.750 ;
        RECT 104.250 219.470 104.530 219.750 ;
        RECT 107.690 219.470 107.970 219.750 ;
        RECT 108.210 219.470 108.490 219.750 ;
        RECT 101.570 217.270 101.850 217.550 ;
        RECT 102.090 217.270 102.370 217.550 ;
        RECT 101.570 215.510 101.850 215.790 ;
        RECT 102.090 215.510 102.370 215.790 ;
        RECT 101.570 214.630 101.850 214.910 ;
        RECT 102.090 214.630 102.370 214.910 ;
        RECT 101.570 211.110 101.850 211.390 ;
        RECT 102.090 211.110 102.370 211.390 ;
        RECT 101.570 210.230 101.850 210.510 ;
        RECT 102.090 210.230 102.370 210.510 ;
        RECT 103.730 216.830 104.010 217.110 ;
        RECT 104.250 216.830 104.530 217.110 ;
        RECT 109.850 218.150 110.130 218.430 ;
        RECT 110.370 218.150 110.650 218.430 ;
        RECT 107.690 216.830 107.970 217.110 ;
        RECT 108.210 216.830 108.490 217.110 ;
        RECT 103.730 214.190 104.010 214.470 ;
        RECT 104.250 214.190 104.530 214.470 ;
        RECT 107.690 214.190 107.970 214.470 ;
        RECT 108.210 214.190 108.490 214.470 ;
        RECT 103.730 213.310 104.010 213.590 ;
        RECT 104.250 213.310 104.530 213.590 ;
        RECT 103.730 212.430 104.010 212.710 ;
        RECT 104.250 212.430 104.530 212.710 ;
        RECT 107.690 212.430 107.970 212.710 ;
        RECT 108.210 212.430 108.490 212.710 ;
        RECT 107.690 211.550 107.970 211.830 ;
        RECT 108.210 211.550 108.490 211.830 ;
        RECT 103.730 209.790 104.010 210.070 ;
        RECT 104.250 209.790 104.530 210.070 ;
        RECT 109.850 212.870 110.130 213.150 ;
        RECT 110.370 212.870 110.650 213.150 ;
        RECT 107.690 209.790 107.970 210.070 ;
        RECT 108.210 209.790 108.490 210.070 ;
        RECT 103.730 207.150 104.010 207.430 ;
        RECT 104.250 207.150 104.530 207.430 ;
        RECT 107.690 207.150 107.970 207.430 ;
        RECT 108.210 207.150 108.490 207.430 ;
        RECT 109.850 208.470 110.130 208.750 ;
        RECT 110.370 208.470 110.650 208.750 ;
        RECT 109.770 207.590 110.050 207.870 ;
        RECT 110.290 207.590 110.570 207.870 ;
        RECT 103.730 205.390 104.010 205.670 ;
        RECT 104.250 205.390 104.530 205.670 ;
        RECT 107.690 205.390 107.970 205.670 ;
        RECT 108.210 205.390 108.490 205.670 ;
        RECT 103.730 204.510 104.010 204.790 ;
        RECT 104.250 204.510 104.530 204.790 ;
        RECT 107.690 204.510 107.970 204.790 ;
        RECT 108.210 204.510 108.490 204.790 ;
        RECT 109.770 204.070 110.050 204.350 ;
        RECT 110.290 204.070 110.570 204.350 ;
        RECT 103.730 203.630 104.010 203.910 ;
        RECT 104.250 203.630 104.530 203.910 ;
        RECT 107.690 203.630 107.970 203.910 ;
        RECT 108.210 203.630 108.490 203.910 ;
        RECT 103.730 202.750 104.010 203.030 ;
        RECT 104.250 202.750 104.530 203.030 ;
        RECT 107.690 202.750 107.970 203.030 ;
        RECT 108.210 202.750 108.490 203.030 ;
        RECT 90.970 201.870 91.250 202.150 ;
        RECT 91.490 201.870 91.770 202.150 ;
        RECT 94.930 201.870 95.210 202.150 ;
        RECT 95.450 201.870 95.730 202.150 ;
        RECT 116.250 221.230 116.530 221.510 ;
        RECT 116.770 221.230 117.050 221.510 ;
        RECT 116.170 220.350 116.450 220.630 ;
        RECT 116.690 220.350 116.970 220.630 ;
        RECT 120.130 220.350 120.410 220.630 ;
        RECT 120.650 220.350 120.930 220.630 ;
        RECT 116.170 219.470 116.450 219.750 ;
        RECT 116.690 219.470 116.970 219.750 ;
        RECT 116.170 218.590 116.450 218.870 ;
        RECT 116.690 218.590 116.970 218.870 ;
        RECT 120.130 218.590 120.410 218.870 ;
        RECT 120.650 218.590 120.930 218.870 ;
        RECT 120.130 217.710 120.410 217.990 ;
        RECT 120.650 217.710 120.930 217.990 ;
        RECT 114.010 217.270 114.290 217.550 ;
        RECT 114.530 217.270 114.810 217.550 ;
        RECT 114.170 216.390 114.450 216.670 ;
        RECT 114.690 216.390 114.970 216.670 ;
        RECT 116.170 215.950 116.450 216.230 ;
        RECT 116.690 215.950 116.970 216.230 ;
        RECT 120.130 215.950 120.410 216.230 ;
        RECT 120.650 215.950 120.930 216.230 ;
        RECT 116.170 215.070 116.450 215.350 ;
        RECT 116.690 215.070 116.970 215.350 ;
        RECT 116.170 214.190 116.450 214.470 ;
        RECT 116.690 214.190 116.970 214.470 ;
        RECT 120.130 214.190 120.410 214.470 ;
        RECT 120.650 214.190 120.930 214.470 ;
        RECT 116.170 213.310 116.450 213.590 ;
        RECT 116.690 213.310 116.970 213.590 ;
        RECT 114.010 211.110 114.290 211.390 ;
        RECT 114.530 211.110 114.810 211.390 ;
        RECT 116.170 212.430 116.450 212.710 ;
        RECT 116.690 212.430 116.970 212.710 ;
        RECT 120.130 212.430 120.410 212.710 ;
        RECT 120.650 212.430 120.930 212.710 ;
        RECT 116.170 211.550 116.450 211.830 ;
        RECT 116.690 211.550 116.970 211.830 ;
        RECT 114.170 210.230 114.450 210.510 ;
        RECT 114.690 210.230 114.970 210.510 ;
        RECT 116.170 209.790 116.450 210.070 ;
        RECT 116.690 209.790 116.970 210.070 ;
        RECT 120.130 209.790 120.410 210.070 ;
        RECT 120.650 209.790 120.930 210.070 ;
        RECT 116.330 208.910 116.610 209.190 ;
        RECT 116.850 208.910 117.130 209.190 ;
        RECT 114.010 207.590 114.290 207.870 ;
        RECT 114.530 207.590 114.810 207.870 ;
        RECT 116.170 208.030 116.450 208.310 ;
        RECT 116.690 208.030 116.970 208.310 ;
        RECT 120.130 208.030 120.410 208.310 ;
        RECT 120.650 208.030 120.930 208.310 ;
        RECT 116.170 206.270 116.450 206.550 ;
        RECT 116.690 206.270 116.970 206.550 ;
        RECT 114.010 205.830 114.290 206.110 ;
        RECT 114.530 205.830 114.810 206.110 ;
        RECT 116.170 205.390 116.450 205.670 ;
        RECT 116.690 205.390 116.970 205.670 ;
        RECT 120.130 205.390 120.410 205.670 ;
        RECT 120.650 205.390 120.930 205.670 ;
        RECT 116.170 204.510 116.450 204.790 ;
        RECT 116.690 204.510 116.970 204.790 ;
        RECT 114.170 204.070 114.450 204.350 ;
        RECT 114.690 204.070 114.970 204.350 ;
        RECT 116.170 203.630 116.450 203.910 ;
        RECT 116.690 203.630 116.970 203.910 ;
        RECT 120.130 203.630 120.410 203.910 ;
        RECT 120.650 203.630 120.930 203.910 ;
        RECT 116.170 202.750 116.450 203.030 ;
        RECT 116.690 202.750 116.970 203.030 ;
        RECT 120.130 202.750 120.410 203.030 ;
        RECT 120.650 202.750 120.930 203.030 ;
        RECT 103.730 201.870 104.010 202.150 ;
        RECT 104.250 201.870 104.530 202.150 ;
        RECT 107.690 201.870 107.970 202.150 ;
        RECT 108.210 201.870 108.490 202.150 ;
        RECT 116.170 201.870 116.450 202.150 ;
        RECT 116.690 201.870 116.970 202.150 ;
        RECT 120.130 201.870 120.410 202.150 ;
        RECT 120.650 201.870 120.930 202.150 ;
        RECT 133.290 219.430 133.630 219.770 ;
        RECT 13.290 200.540 13.570 200.820 ;
        RECT 13.810 200.540 14.090 200.820 ;
        RECT 34.170 200.540 34.450 200.820 ;
        RECT 34.690 200.540 34.970 200.820 ;
        RECT 38.490 200.540 38.770 200.820 ;
        RECT 39.010 200.540 39.290 200.820 ;
        RECT 59.370 200.540 59.650 200.820 ;
        RECT 59.890 200.540 60.170 200.820 ;
        RECT 63.690 200.540 63.970 200.820 ;
        RECT 64.210 200.540 64.490 200.820 ;
        RECT 84.570 200.540 84.850 200.820 ;
        RECT 85.090 200.540 85.370 200.820 ;
        RECT 88.890 200.540 89.170 200.820 ;
        RECT 89.410 200.540 89.690 200.820 ;
        RECT 109.770 200.540 110.050 200.820 ;
        RECT 110.290 200.540 110.570 200.820 ;
        RECT 111.860 200.560 112.140 200.840 ;
        RECT 132.110 200.510 132.450 200.850 ;
        RECT 15.370 199.650 15.650 199.930 ;
        RECT 15.890 199.650 16.170 199.930 ;
        RECT 32.090 199.650 32.370 199.930 ;
        RECT 32.610 199.650 32.890 199.930 ;
        RECT 40.570 199.650 40.850 199.930 ;
        RECT 41.090 199.650 41.370 199.930 ;
        RECT 57.290 199.650 57.570 199.930 ;
        RECT 57.810 199.650 58.090 199.930 ;
        RECT 65.770 199.650 66.050 199.930 ;
        RECT 66.290 199.650 66.570 199.930 ;
        RECT 82.490 199.650 82.770 199.930 ;
        RECT 83.010 199.650 83.290 199.930 ;
        RECT 90.970 199.650 91.250 199.930 ;
        RECT 91.490 199.650 91.770 199.930 ;
        RECT 107.690 199.650 107.970 199.930 ;
        RECT 108.210 199.650 108.490 199.930 ;
        RECT 116.170 199.650 116.450 199.930 ;
        RECT 116.690 199.650 116.970 199.930 ;
        RECT 15.370 199.130 15.650 199.410 ;
        RECT 15.890 199.130 16.170 199.410 ;
        RECT 32.090 199.130 32.370 199.410 ;
        RECT 32.610 199.130 32.890 199.410 ;
        RECT 40.570 199.130 40.850 199.410 ;
        RECT 41.090 199.130 41.370 199.410 ;
        RECT 57.290 199.130 57.570 199.410 ;
        RECT 57.810 199.130 58.090 199.410 ;
        RECT 65.770 199.130 66.050 199.410 ;
        RECT 66.290 199.130 66.570 199.410 ;
        RECT 82.490 199.130 82.770 199.410 ;
        RECT 83.010 199.130 83.290 199.410 ;
        RECT 90.970 199.130 91.250 199.410 ;
        RECT 91.490 199.130 91.770 199.410 ;
        RECT 107.690 199.130 107.970 199.410 ;
        RECT 108.210 199.130 108.490 199.410 ;
        RECT 116.170 199.130 116.450 199.410 ;
        RECT 116.690 199.130 116.970 199.410 ;
        RECT 19.330 198.210 19.610 198.490 ;
        RECT 19.850 198.210 20.130 198.490 ;
        RECT 22.110 198.210 22.390 198.490 ;
        RECT 22.630 198.210 22.910 198.490 ;
        RECT 25.150 198.210 25.430 198.490 ;
        RECT 25.670 198.210 25.950 198.490 ;
        RECT 28.130 198.210 28.410 198.490 ;
        RECT 28.650 198.210 28.930 198.490 ;
        RECT 44.530 198.210 44.810 198.490 ;
        RECT 45.050 198.210 45.330 198.490 ;
        RECT 47.310 198.210 47.590 198.490 ;
        RECT 47.830 198.210 48.110 198.490 ;
        RECT 50.350 198.210 50.630 198.490 ;
        RECT 50.870 198.210 51.150 198.490 ;
        RECT 53.330 198.210 53.610 198.490 ;
        RECT 53.850 198.210 54.130 198.490 ;
        RECT 69.730 198.210 70.010 198.490 ;
        RECT 70.250 198.210 70.530 198.490 ;
        RECT 72.510 198.210 72.790 198.490 ;
        RECT 73.030 198.210 73.310 198.490 ;
        RECT 75.550 198.210 75.830 198.490 ;
        RECT 76.070 198.210 76.350 198.490 ;
        RECT 78.530 198.210 78.810 198.490 ;
        RECT 79.050 198.210 79.330 198.490 ;
        RECT 94.930 198.210 95.210 198.490 ;
        RECT 95.450 198.210 95.730 198.490 ;
        RECT 97.710 198.210 97.990 198.490 ;
        RECT 98.230 198.210 98.510 198.490 ;
        RECT 100.750 198.210 101.030 198.490 ;
        RECT 101.270 198.210 101.550 198.490 ;
        RECT 103.730 198.210 104.010 198.490 ;
        RECT 104.250 198.210 104.530 198.490 ;
        RECT 120.130 198.210 120.410 198.490 ;
        RECT 120.650 198.210 120.930 198.490 ;
        RECT 19.330 197.690 19.610 197.970 ;
        RECT 19.850 197.690 20.130 197.970 ;
        RECT 22.110 197.690 22.390 197.970 ;
        RECT 22.630 197.690 22.910 197.970 ;
        RECT 25.150 197.690 25.430 197.970 ;
        RECT 25.670 197.690 25.950 197.970 ;
        RECT 28.130 197.690 28.410 197.970 ;
        RECT 28.650 197.690 28.930 197.970 ;
        RECT 44.530 197.690 44.810 197.970 ;
        RECT 45.050 197.690 45.330 197.970 ;
        RECT 47.310 197.690 47.590 197.970 ;
        RECT 47.830 197.690 48.110 197.970 ;
        RECT 50.350 197.690 50.630 197.970 ;
        RECT 50.870 197.690 51.150 197.970 ;
        RECT 53.330 197.690 53.610 197.970 ;
        RECT 53.850 197.690 54.130 197.970 ;
        RECT 69.730 197.690 70.010 197.970 ;
        RECT 70.250 197.690 70.530 197.970 ;
        RECT 72.510 197.690 72.790 197.970 ;
        RECT 73.030 197.690 73.310 197.970 ;
        RECT 75.550 197.690 75.830 197.970 ;
        RECT 76.070 197.690 76.350 197.970 ;
        RECT 78.530 197.690 78.810 197.970 ;
        RECT 79.050 197.690 79.330 197.970 ;
        RECT 94.930 197.690 95.210 197.970 ;
        RECT 95.450 197.690 95.730 197.970 ;
        RECT 97.710 197.690 97.990 197.970 ;
        RECT 98.230 197.690 98.510 197.970 ;
        RECT 100.750 197.690 101.030 197.970 ;
        RECT 101.270 197.690 101.550 197.970 ;
        RECT 103.730 197.690 104.010 197.970 ;
        RECT 104.250 197.690 104.530 197.970 ;
        RECT 120.130 197.690 120.410 197.970 ;
        RECT 120.650 197.690 120.930 197.970 ;
        RECT 2.660 183.470 2.940 183.750 ;
        RECT 2.660 182.950 2.940 183.230 ;
        RECT 19.230 194.610 19.510 194.890 ;
        RECT 19.750 194.610 20.030 194.890 ;
        RECT 28.030 194.610 28.310 194.890 ;
        RECT 28.550 194.610 28.830 194.890 ;
        RECT 44.430 194.610 44.710 194.890 ;
        RECT 44.950 194.610 45.230 194.890 ;
        RECT 53.230 194.610 53.510 194.890 ;
        RECT 53.750 194.610 54.030 194.890 ;
        RECT 69.630 194.610 69.910 194.890 ;
        RECT 70.150 194.610 70.430 194.890 ;
        RECT 78.430 194.610 78.710 194.890 ;
        RECT 78.950 194.610 79.230 194.890 ;
        RECT 94.830 194.610 95.110 194.890 ;
        RECT 95.350 194.610 95.630 194.890 ;
        RECT 103.630 194.610 103.910 194.890 ;
        RECT 104.150 194.610 104.430 194.890 ;
        RECT 120.030 194.610 120.310 194.890 ;
        RECT 120.550 194.610 120.830 194.890 ;
        RECT 19.230 194.090 19.510 194.370 ;
        RECT 19.750 194.090 20.030 194.370 ;
        RECT 28.030 194.090 28.310 194.370 ;
        RECT 28.550 194.090 28.830 194.370 ;
        RECT 44.430 194.090 44.710 194.370 ;
        RECT 44.950 194.090 45.230 194.370 ;
        RECT 53.230 194.090 53.510 194.370 ;
        RECT 53.750 194.090 54.030 194.370 ;
        RECT 69.630 194.090 69.910 194.370 ;
        RECT 70.150 194.090 70.430 194.370 ;
        RECT 78.430 194.090 78.710 194.370 ;
        RECT 78.950 194.090 79.230 194.370 ;
        RECT 94.830 194.090 95.110 194.370 ;
        RECT 95.350 194.090 95.630 194.370 ;
        RECT 103.630 194.090 103.910 194.370 ;
        RECT 104.150 194.090 104.430 194.370 ;
        RECT 120.030 194.090 120.310 194.370 ;
        RECT 120.550 194.090 120.830 194.370 ;
        RECT 15.270 191.010 15.550 191.290 ;
        RECT 15.790 191.010 16.070 191.290 ;
        RECT 31.990 191.010 32.270 191.290 ;
        RECT 32.510 191.010 32.790 191.290 ;
        RECT 40.470 191.010 40.750 191.290 ;
        RECT 40.990 191.010 41.270 191.290 ;
        RECT 57.190 191.010 57.470 191.290 ;
        RECT 57.710 191.010 57.990 191.290 ;
        RECT 65.670 191.010 65.950 191.290 ;
        RECT 66.190 191.010 66.470 191.290 ;
        RECT 82.390 191.010 82.670 191.290 ;
        RECT 82.910 191.010 83.190 191.290 ;
        RECT 90.870 191.010 91.150 191.290 ;
        RECT 91.390 191.010 91.670 191.290 ;
        RECT 107.590 191.010 107.870 191.290 ;
        RECT 108.110 191.010 108.390 191.290 ;
        RECT 116.070 191.010 116.350 191.290 ;
        RECT 116.590 191.010 116.870 191.290 ;
        RECT 15.270 190.490 15.550 190.770 ;
        RECT 15.790 190.490 16.070 190.770 ;
        RECT 31.990 190.490 32.270 190.770 ;
        RECT 32.510 190.490 32.790 190.770 ;
        RECT 40.470 190.490 40.750 190.770 ;
        RECT 40.990 190.490 41.270 190.770 ;
        RECT 57.190 190.490 57.470 190.770 ;
        RECT 57.710 190.490 57.990 190.770 ;
        RECT 65.670 190.490 65.950 190.770 ;
        RECT 66.190 190.490 66.470 190.770 ;
        RECT 82.390 190.490 82.670 190.770 ;
        RECT 82.910 190.490 83.190 190.770 ;
        RECT 90.870 190.490 91.150 190.770 ;
        RECT 91.390 190.490 91.670 190.770 ;
        RECT 107.590 190.490 107.870 190.770 ;
        RECT 108.110 190.490 108.390 190.770 ;
        RECT 116.070 190.490 116.350 190.770 ;
        RECT 116.590 190.490 116.870 190.770 ;
        RECT 15.270 187.170 15.550 187.450 ;
        RECT 15.790 187.170 16.070 187.450 ;
        RECT 19.230 187.170 19.510 187.450 ;
        RECT 19.750 187.170 20.030 187.450 ;
        RECT 28.030 187.170 28.310 187.450 ;
        RECT 28.550 187.170 28.830 187.450 ;
        RECT 31.990 187.170 32.270 187.450 ;
        RECT 32.510 187.170 32.790 187.450 ;
        RECT 15.270 186.290 15.550 186.570 ;
        RECT 15.790 186.290 16.070 186.570 ;
        RECT 19.230 186.290 19.510 186.570 ;
        RECT 19.750 186.290 20.030 186.570 ;
        RECT 19.230 185.580 19.510 185.860 ;
        RECT 19.750 185.580 20.030 185.860 ;
        RECT 13.110 183.210 13.390 183.490 ;
        RECT 13.630 183.210 13.910 183.490 ;
        RECT 15.270 184.530 15.550 184.810 ;
        RECT 15.790 184.530 16.070 184.810 ;
        RECT 19.230 184.530 19.510 184.810 ;
        RECT 19.750 184.530 20.030 184.810 ;
        RECT 15.270 183.650 15.550 183.930 ;
        RECT 15.790 183.650 16.070 183.930 ;
        RECT 15.270 181.890 15.550 182.170 ;
        RECT 15.790 181.890 16.070 182.170 ;
        RECT 19.230 181.890 19.510 182.170 ;
        RECT 19.750 181.890 20.030 182.170 ;
        RECT 15.270 180.130 15.550 180.410 ;
        RECT 15.790 180.130 16.070 180.410 ;
        RECT 19.230 180.130 19.510 180.410 ;
        RECT 19.750 180.130 20.030 180.410 ;
        RECT 19.230 179.250 19.510 179.530 ;
        RECT 19.750 179.250 20.030 179.530 ;
        RECT 13.110 178.810 13.390 179.090 ;
        RECT 13.630 178.810 13.910 179.090 ;
        RECT 15.270 177.490 15.550 177.770 ;
        RECT 15.790 177.490 16.070 177.770 ;
        RECT 19.230 177.490 19.510 177.770 ;
        RECT 19.750 177.490 20.030 177.770 ;
        RECT 15.270 176.610 15.550 176.890 ;
        RECT 15.790 176.610 16.070 176.890 ;
        RECT 15.270 175.730 15.550 176.010 ;
        RECT 15.790 175.730 16.070 176.010 ;
        RECT 19.230 175.730 19.510 176.010 ;
        RECT 19.750 175.730 20.030 176.010 ;
        RECT 21.390 174.410 21.670 174.690 ;
        RECT 21.910 174.410 22.190 174.690 ;
        RECT 15.270 173.970 15.550 174.250 ;
        RECT 15.790 173.970 16.070 174.250 ;
        RECT 19.230 173.970 19.510 174.250 ;
        RECT 19.750 173.970 20.030 174.250 ;
        RECT 15.270 173.090 15.550 173.370 ;
        RECT 15.790 173.090 16.070 173.370 ;
        RECT 15.270 171.330 15.550 171.610 ;
        RECT 15.790 171.330 16.070 171.610 ;
        RECT 13.110 170.890 13.390 171.170 ;
        RECT 13.630 170.890 13.910 171.170 ;
        RECT 21.390 171.770 21.670 172.050 ;
        RECT 21.910 171.770 22.190 172.050 ;
        RECT 19.230 171.330 19.510 171.610 ;
        RECT 19.750 171.330 20.030 171.610 ;
        RECT 15.270 169.570 15.550 169.850 ;
        RECT 15.790 169.570 16.070 169.850 ;
        RECT 15.270 168.690 15.550 168.970 ;
        RECT 15.790 168.690 16.070 168.970 ;
        RECT 19.230 168.690 19.510 168.970 ;
        RECT 19.750 168.690 20.030 168.970 ;
        RECT 15.270 166.930 15.550 167.210 ;
        RECT 15.790 166.930 16.070 167.210 ;
        RECT 19.230 166.930 19.510 167.210 ;
        RECT 19.750 166.930 20.030 167.210 ;
        RECT 18.190 166.310 18.470 166.590 ;
        RECT 18.190 165.790 18.470 166.070 ;
        RECT 15.270 165.170 15.550 165.450 ;
        RECT 15.790 165.170 16.070 165.450 ;
        RECT 19.230 165.170 19.510 165.450 ;
        RECT 19.750 165.170 20.030 165.450 ;
        RECT 15.270 164.290 15.550 164.570 ;
        RECT 15.790 164.290 16.070 164.570 ;
        RECT 19.230 164.290 19.510 164.570 ;
        RECT 19.750 164.290 20.030 164.570 ;
        RECT 15.270 162.530 15.550 162.810 ;
        RECT 15.790 162.530 16.070 162.810 ;
        RECT 19.230 162.530 19.510 162.810 ;
        RECT 19.750 162.530 20.030 162.810 ;
        RECT 17.405 161.910 17.685 162.190 ;
        RECT 13.110 161.210 13.390 161.490 ;
        RECT 13.630 161.210 13.910 161.490 ;
        RECT 17.405 161.390 17.685 161.670 ;
        RECT 15.270 160.770 15.550 161.050 ;
        RECT 15.790 160.770 16.070 161.050 ;
        RECT 19.230 160.770 19.510 161.050 ;
        RECT 19.750 160.770 20.030 161.050 ;
        RECT 15.270 159.890 15.550 160.170 ;
        RECT 15.790 159.890 16.070 160.170 ;
        RECT 19.230 159.890 19.510 160.170 ;
        RECT 19.750 159.890 20.030 160.170 ;
        RECT 15.270 158.130 15.550 158.410 ;
        RECT 15.790 158.130 16.070 158.410 ;
        RECT 19.230 158.130 19.510 158.410 ;
        RECT 19.750 158.130 20.030 158.410 ;
        RECT 16.690 157.510 16.970 157.790 ;
        RECT 13.270 156.810 13.550 157.090 ;
        RECT 13.790 156.810 14.070 157.090 ;
        RECT 16.690 156.990 16.970 157.270 ;
        RECT 19.230 157.250 19.510 157.530 ;
        RECT 19.750 157.250 20.030 157.530 ;
        RECT 15.270 156.370 15.550 156.650 ;
        RECT 15.790 156.370 16.070 156.650 ;
        RECT 19.230 156.370 19.510 156.650 ;
        RECT 19.750 156.370 20.030 156.650 ;
        RECT 15.270 155.490 15.550 155.770 ;
        RECT 15.790 155.490 16.070 155.770 ;
        RECT 19.230 155.490 19.510 155.770 ;
        RECT 19.750 155.490 20.030 155.770 ;
        RECT 15.270 153.730 15.550 154.010 ;
        RECT 15.790 153.730 16.070 154.010 ;
        RECT 19.230 153.730 19.510 154.010 ;
        RECT 19.750 153.730 20.030 154.010 ;
        RECT 15.270 151.970 15.550 152.250 ;
        RECT 15.790 151.970 16.070 152.250 ;
        RECT 19.230 151.970 19.510 152.250 ;
        RECT 19.750 151.970 20.030 152.250 ;
        RECT 13.110 150.650 13.390 150.930 ;
        RECT 13.630 150.650 13.910 150.930 ;
        RECT 21.390 150.650 21.670 150.930 ;
        RECT 21.910 150.650 22.190 150.930 ;
        RECT 13.110 148.890 13.390 149.170 ;
        RECT 13.630 148.890 13.910 149.170 ;
        RECT 13.110 147.130 13.390 147.410 ;
        RECT 13.630 147.130 13.910 147.410 ;
        RECT 15.270 148.450 15.550 148.730 ;
        RECT 15.790 148.450 16.070 148.730 ;
        RECT 19.230 148.450 19.510 148.730 ;
        RECT 19.750 148.450 20.030 148.730 ;
        RECT 15.270 147.570 15.550 147.850 ;
        RECT 15.790 147.570 16.070 147.850 ;
        RECT 13.270 145.370 13.550 145.650 ;
        RECT 13.790 145.370 14.070 145.650 ;
        RECT 15.270 144.930 15.550 145.210 ;
        RECT 15.790 144.930 16.070 145.210 ;
        RECT 19.230 144.930 19.510 145.210 ;
        RECT 19.750 144.930 20.030 145.210 ;
        RECT 15.270 143.170 15.550 143.450 ;
        RECT 15.790 143.170 16.070 143.450 ;
        RECT 19.230 143.170 19.510 143.450 ;
        RECT 19.750 143.170 20.030 143.450 ;
        RECT 19.230 142.290 19.510 142.570 ;
        RECT 19.750 142.290 20.030 142.570 ;
        RECT 15.270 141.410 15.550 141.690 ;
        RECT 15.790 141.410 16.070 141.690 ;
        RECT 15.270 140.530 15.550 140.810 ;
        RECT 15.790 140.530 16.070 140.810 ;
        RECT 13.270 140.090 13.550 140.370 ;
        RECT 13.790 140.090 14.070 140.370 ;
        RECT 15.270 137.890 15.550 138.170 ;
        RECT 15.790 137.890 16.070 138.170 ;
        RECT 19.230 137.890 19.510 138.170 ;
        RECT 19.750 137.890 20.030 138.170 ;
        RECT 19.230 137.010 19.510 137.290 ;
        RECT 19.750 137.010 20.030 137.290 ;
        RECT 13.110 136.570 13.390 136.850 ;
        RECT 13.630 136.570 13.910 136.850 ;
        RECT 15.270 135.250 15.550 135.530 ;
        RECT 15.790 135.250 16.070 135.530 ;
        RECT 19.230 135.250 19.510 135.530 ;
        RECT 19.750 135.250 20.030 135.530 ;
        RECT 40.470 187.170 40.750 187.450 ;
        RECT 40.990 187.170 41.270 187.450 ;
        RECT 44.430 187.170 44.710 187.450 ;
        RECT 44.950 187.170 45.230 187.450 ;
        RECT 28.030 186.290 28.310 186.570 ;
        RECT 28.550 186.290 28.830 186.570 ;
        RECT 31.990 186.290 32.270 186.570 ;
        RECT 32.510 186.290 32.790 186.570 ;
        RECT 27.870 185.410 28.150 185.690 ;
        RECT 28.390 185.410 28.670 185.690 ;
        RECT 28.030 184.530 28.310 184.810 ;
        RECT 28.550 184.530 28.830 184.810 ;
        RECT 31.990 184.530 32.270 184.810 ;
        RECT 32.510 184.530 32.790 184.810 ;
        RECT 31.990 183.650 32.270 183.930 ;
        RECT 32.510 183.650 32.790 183.930 ;
        RECT 33.990 183.210 34.270 183.490 ;
        RECT 34.510 183.210 34.790 183.490 ;
        RECT 28.030 181.890 28.310 182.170 ;
        RECT 28.550 181.890 28.830 182.170 ;
        RECT 31.990 181.890 32.270 182.170 ;
        RECT 32.510 181.890 32.790 182.170 ;
        RECT 28.030 180.130 28.310 180.410 ;
        RECT 28.550 180.130 28.830 180.410 ;
        RECT 31.990 180.130 32.270 180.410 ;
        RECT 32.510 180.130 32.790 180.410 ;
        RECT 28.030 179.250 28.310 179.530 ;
        RECT 28.550 179.250 28.830 179.530 ;
        RECT 34.150 178.810 34.430 179.090 ;
        RECT 34.670 178.810 34.950 179.090 ;
        RECT 28.030 177.490 28.310 177.770 ;
        RECT 28.550 177.490 28.830 177.770 ;
        RECT 31.990 177.490 32.270 177.770 ;
        RECT 32.510 177.490 32.790 177.770 ;
        RECT 31.830 176.610 32.110 176.890 ;
        RECT 32.350 176.610 32.630 176.890 ;
        RECT 28.030 175.730 28.310 176.010 ;
        RECT 28.550 175.730 28.830 176.010 ;
        RECT 31.990 175.730 32.270 176.010 ;
        RECT 32.510 175.730 32.790 176.010 ;
        RECT 25.870 174.410 26.150 174.690 ;
        RECT 26.390 174.410 26.670 174.690 ;
        RECT 28.030 173.970 28.310 174.250 ;
        RECT 28.550 173.970 28.830 174.250 ;
        RECT 31.990 173.970 32.270 174.250 ;
        RECT 32.510 173.970 32.790 174.250 ;
        RECT 31.990 173.090 32.270 173.370 ;
        RECT 32.510 173.090 32.790 173.370 ;
        RECT 25.870 171.770 26.150 172.050 ;
        RECT 26.390 171.770 26.670 172.050 ;
        RECT 28.030 171.330 28.310 171.610 ;
        RECT 28.550 171.330 28.830 171.610 ;
        RECT 31.990 171.330 32.270 171.610 ;
        RECT 32.510 171.330 32.790 171.610 ;
        RECT 33.990 170.890 34.270 171.170 ;
        RECT 34.510 170.890 34.790 171.170 ;
        RECT 31.990 169.570 32.270 169.850 ;
        RECT 32.510 169.570 32.790 169.850 ;
        RECT 28.030 168.690 28.310 168.970 ;
        RECT 28.550 168.690 28.830 168.970 ;
        RECT 31.990 168.690 32.270 168.970 ;
        RECT 32.510 168.690 32.790 168.970 ;
        RECT 28.030 166.930 28.310 167.210 ;
        RECT 28.550 166.930 28.830 167.210 ;
        RECT 29.590 166.310 29.870 166.590 ;
        RECT 31.990 166.930 32.270 167.210 ;
        RECT 32.510 166.930 32.790 167.210 ;
        RECT 29.590 165.790 29.870 166.070 ;
        RECT 28.030 165.170 28.310 165.450 ;
        RECT 28.550 165.170 28.830 165.450 ;
        RECT 31.990 165.170 32.270 165.450 ;
        RECT 32.510 165.170 32.790 165.450 ;
        RECT 28.030 164.290 28.310 164.570 ;
        RECT 28.550 164.290 28.830 164.570 ;
        RECT 31.990 164.290 32.270 164.570 ;
        RECT 32.510 164.290 32.790 164.570 ;
        RECT 28.030 162.530 28.310 162.810 ;
        RECT 28.550 162.530 28.830 162.810 ;
        RECT 30.375 161.910 30.655 162.190 ;
        RECT 31.990 162.530 32.270 162.810 ;
        RECT 32.510 162.530 32.790 162.810 ;
        RECT 30.375 161.390 30.655 161.670 ;
        RECT 34.150 161.210 34.430 161.490 ;
        RECT 34.670 161.210 34.950 161.490 ;
        RECT 28.030 160.770 28.310 161.050 ;
        RECT 28.550 160.770 28.830 161.050 ;
        RECT 31.990 160.770 32.270 161.050 ;
        RECT 32.510 160.770 32.790 161.050 ;
        RECT 28.030 159.890 28.310 160.170 ;
        RECT 28.550 159.890 28.830 160.170 ;
        RECT 31.990 159.890 32.270 160.170 ;
        RECT 32.510 159.890 32.790 160.170 ;
        RECT 28.030 158.130 28.310 158.410 ;
        RECT 28.550 158.130 28.830 158.410 ;
        RECT 31.990 158.130 32.270 158.410 ;
        RECT 32.510 158.130 32.790 158.410 ;
        RECT 28.030 157.250 28.310 157.530 ;
        RECT 28.550 157.250 28.830 157.530 ;
        RECT 31.090 157.510 31.370 157.790 ;
        RECT 31.090 156.990 31.370 157.270 ;
        RECT 33.990 156.810 34.270 157.090 ;
        RECT 34.510 156.810 34.790 157.090 ;
        RECT 28.030 156.370 28.310 156.650 ;
        RECT 28.550 156.370 28.830 156.650 ;
        RECT 31.990 156.370 32.270 156.650 ;
        RECT 32.510 156.370 32.790 156.650 ;
        RECT 28.030 155.490 28.310 155.770 ;
        RECT 28.550 155.490 28.830 155.770 ;
        RECT 31.990 155.490 32.270 155.770 ;
        RECT 32.510 155.490 32.790 155.770 ;
        RECT 28.030 153.730 28.310 154.010 ;
        RECT 28.550 153.730 28.830 154.010 ;
        RECT 31.990 153.730 32.270 154.010 ;
        RECT 32.510 153.730 32.790 154.010 ;
        RECT 28.030 151.970 28.310 152.250 ;
        RECT 28.550 151.970 28.830 152.250 ;
        RECT 31.990 151.970 32.270 152.250 ;
        RECT 32.510 151.970 32.790 152.250 ;
        RECT 25.710 150.650 25.990 150.930 ;
        RECT 26.230 150.650 26.510 150.930 ;
        RECT 34.150 150.650 34.430 150.930 ;
        RECT 34.670 150.650 34.950 150.930 ;
        RECT 28.030 148.450 28.310 148.730 ;
        RECT 28.550 148.450 28.830 148.730 ;
        RECT 31.990 148.450 32.270 148.730 ;
        RECT 32.510 148.450 32.790 148.730 ;
        RECT 31.990 147.570 32.270 147.850 ;
        RECT 32.510 147.570 32.790 147.850 ;
        RECT 33.990 148.890 34.270 149.170 ;
        RECT 34.510 148.890 34.790 149.170 ;
        RECT 34.150 147.130 34.430 147.410 ;
        RECT 34.670 147.130 34.950 147.410 ;
        RECT 28.030 144.930 28.310 145.210 ;
        RECT 28.550 144.930 28.830 145.210 ;
        RECT 31.990 144.930 32.270 145.210 ;
        RECT 32.510 144.930 32.790 145.210 ;
        RECT 33.990 145.370 34.270 145.650 ;
        RECT 34.510 145.370 34.790 145.650 ;
        RECT 28.030 143.170 28.310 143.450 ;
        RECT 28.550 143.170 28.830 143.450 ;
        RECT 31.990 143.170 32.270 143.450 ;
        RECT 32.510 143.170 32.790 143.450 ;
        RECT 28.030 142.290 28.310 142.570 ;
        RECT 28.550 142.290 28.830 142.570 ;
        RECT 31.990 141.410 32.270 141.690 ;
        RECT 32.510 141.410 32.790 141.690 ;
        RECT 31.990 140.530 32.270 140.810 ;
        RECT 32.510 140.530 32.790 140.810 ;
        RECT 33.990 140.090 34.270 140.370 ;
        RECT 34.510 140.090 34.790 140.370 ;
        RECT 28.030 137.890 28.310 138.170 ;
        RECT 28.550 137.890 28.830 138.170 ;
        RECT 31.990 137.890 32.270 138.170 ;
        RECT 32.510 137.890 32.790 138.170 ;
        RECT 28.030 137.010 28.310 137.290 ;
        RECT 28.550 137.010 28.830 137.290 ;
        RECT 34.150 136.570 34.430 136.850 ;
        RECT 34.670 136.570 34.950 136.850 ;
        RECT 28.030 135.250 28.310 135.530 ;
        RECT 28.550 135.250 28.830 135.530 ;
        RECT 31.990 135.250 32.270 135.530 ;
        RECT 32.510 135.250 32.790 135.530 ;
        RECT 15.270 134.370 15.550 134.650 ;
        RECT 15.790 134.370 16.070 134.650 ;
        RECT 19.230 134.370 19.510 134.650 ;
        RECT 19.750 134.370 20.030 134.650 ;
        RECT 53.230 187.170 53.510 187.450 ;
        RECT 53.750 187.170 54.030 187.450 ;
        RECT 57.190 187.170 57.470 187.450 ;
        RECT 57.710 187.170 57.990 187.450 ;
        RECT 40.470 186.290 40.750 186.570 ;
        RECT 40.990 186.290 41.270 186.570 ;
        RECT 44.430 186.290 44.710 186.570 ;
        RECT 44.950 186.290 45.230 186.570 ;
        RECT 44.430 185.580 44.710 185.860 ;
        RECT 44.950 185.580 45.230 185.860 ;
        RECT 38.310 183.210 38.590 183.490 ;
        RECT 38.830 183.210 39.110 183.490 ;
        RECT 40.470 184.530 40.750 184.810 ;
        RECT 40.990 184.530 41.270 184.810 ;
        RECT 44.430 184.530 44.710 184.810 ;
        RECT 44.950 184.530 45.230 184.810 ;
        RECT 40.470 183.650 40.750 183.930 ;
        RECT 40.990 183.650 41.270 183.930 ;
        RECT 40.470 181.890 40.750 182.170 ;
        RECT 40.990 181.890 41.270 182.170 ;
        RECT 44.430 181.890 44.710 182.170 ;
        RECT 44.950 181.890 45.230 182.170 ;
        RECT 40.470 180.130 40.750 180.410 ;
        RECT 40.990 180.130 41.270 180.410 ;
        RECT 44.430 180.130 44.710 180.410 ;
        RECT 44.950 180.130 45.230 180.410 ;
        RECT 44.430 179.250 44.710 179.530 ;
        RECT 44.950 179.250 45.230 179.530 ;
        RECT 38.310 178.810 38.590 179.090 ;
        RECT 38.830 178.810 39.110 179.090 ;
        RECT 40.470 177.490 40.750 177.770 ;
        RECT 40.990 177.490 41.270 177.770 ;
        RECT 44.430 177.490 44.710 177.770 ;
        RECT 44.950 177.490 45.230 177.770 ;
        RECT 40.470 176.610 40.750 176.890 ;
        RECT 40.990 176.610 41.270 176.890 ;
        RECT 40.470 175.730 40.750 176.010 ;
        RECT 40.990 175.730 41.270 176.010 ;
        RECT 44.430 175.730 44.710 176.010 ;
        RECT 44.950 175.730 45.230 176.010 ;
        RECT 46.590 174.410 46.870 174.690 ;
        RECT 47.110 174.410 47.390 174.690 ;
        RECT 40.470 173.970 40.750 174.250 ;
        RECT 40.990 173.970 41.270 174.250 ;
        RECT 44.430 173.970 44.710 174.250 ;
        RECT 44.950 173.970 45.230 174.250 ;
        RECT 40.470 173.090 40.750 173.370 ;
        RECT 40.990 173.090 41.270 173.370 ;
        RECT 40.470 171.330 40.750 171.610 ;
        RECT 40.990 171.330 41.270 171.610 ;
        RECT 38.310 170.890 38.590 171.170 ;
        RECT 38.830 170.890 39.110 171.170 ;
        RECT 46.590 171.770 46.870 172.050 ;
        RECT 47.110 171.770 47.390 172.050 ;
        RECT 44.430 171.330 44.710 171.610 ;
        RECT 44.950 171.330 45.230 171.610 ;
        RECT 40.470 169.570 40.750 169.850 ;
        RECT 40.990 169.570 41.270 169.850 ;
        RECT 40.470 168.690 40.750 168.970 ;
        RECT 40.990 168.690 41.270 168.970 ;
        RECT 44.430 168.690 44.710 168.970 ;
        RECT 44.950 168.690 45.230 168.970 ;
        RECT 40.470 166.930 40.750 167.210 ;
        RECT 40.990 166.930 41.270 167.210 ;
        RECT 44.430 166.930 44.710 167.210 ;
        RECT 44.950 166.930 45.230 167.210 ;
        RECT 43.390 166.310 43.670 166.590 ;
        RECT 43.390 165.790 43.670 166.070 ;
        RECT 40.470 165.170 40.750 165.450 ;
        RECT 40.990 165.170 41.270 165.450 ;
        RECT 44.430 165.170 44.710 165.450 ;
        RECT 44.950 165.170 45.230 165.450 ;
        RECT 40.470 164.290 40.750 164.570 ;
        RECT 40.990 164.290 41.270 164.570 ;
        RECT 44.430 164.290 44.710 164.570 ;
        RECT 44.950 164.290 45.230 164.570 ;
        RECT 40.470 162.530 40.750 162.810 ;
        RECT 40.990 162.530 41.270 162.810 ;
        RECT 44.430 162.530 44.710 162.810 ;
        RECT 44.950 162.530 45.230 162.810 ;
        RECT 42.605 161.910 42.885 162.190 ;
        RECT 38.310 161.210 38.590 161.490 ;
        RECT 38.830 161.210 39.110 161.490 ;
        RECT 42.605 161.390 42.885 161.670 ;
        RECT 40.470 160.770 40.750 161.050 ;
        RECT 40.990 160.770 41.270 161.050 ;
        RECT 44.430 160.770 44.710 161.050 ;
        RECT 44.950 160.770 45.230 161.050 ;
        RECT 40.470 159.890 40.750 160.170 ;
        RECT 40.990 159.890 41.270 160.170 ;
        RECT 44.430 159.890 44.710 160.170 ;
        RECT 44.950 159.890 45.230 160.170 ;
        RECT 40.470 158.130 40.750 158.410 ;
        RECT 40.990 158.130 41.270 158.410 ;
        RECT 44.430 158.130 44.710 158.410 ;
        RECT 44.950 158.130 45.230 158.410 ;
        RECT 41.890 157.510 42.170 157.790 ;
        RECT 38.470 156.810 38.750 157.090 ;
        RECT 38.990 156.810 39.270 157.090 ;
        RECT 41.890 156.990 42.170 157.270 ;
        RECT 44.430 157.250 44.710 157.530 ;
        RECT 44.950 157.250 45.230 157.530 ;
        RECT 40.470 156.370 40.750 156.650 ;
        RECT 40.990 156.370 41.270 156.650 ;
        RECT 44.430 156.370 44.710 156.650 ;
        RECT 44.950 156.370 45.230 156.650 ;
        RECT 40.470 155.490 40.750 155.770 ;
        RECT 40.990 155.490 41.270 155.770 ;
        RECT 44.430 155.490 44.710 155.770 ;
        RECT 44.950 155.490 45.230 155.770 ;
        RECT 40.470 153.730 40.750 154.010 ;
        RECT 40.990 153.730 41.270 154.010 ;
        RECT 44.430 153.730 44.710 154.010 ;
        RECT 44.950 153.730 45.230 154.010 ;
        RECT 40.470 151.970 40.750 152.250 ;
        RECT 40.990 151.970 41.270 152.250 ;
        RECT 44.430 151.970 44.710 152.250 ;
        RECT 44.950 151.970 45.230 152.250 ;
        RECT 38.310 150.650 38.590 150.930 ;
        RECT 38.830 150.650 39.110 150.930 ;
        RECT 46.590 150.650 46.870 150.930 ;
        RECT 47.110 150.650 47.390 150.930 ;
        RECT 38.310 148.890 38.590 149.170 ;
        RECT 38.830 148.890 39.110 149.170 ;
        RECT 38.310 147.130 38.590 147.410 ;
        RECT 38.830 147.130 39.110 147.410 ;
        RECT 40.470 148.450 40.750 148.730 ;
        RECT 40.990 148.450 41.270 148.730 ;
        RECT 44.430 148.450 44.710 148.730 ;
        RECT 44.950 148.450 45.230 148.730 ;
        RECT 40.470 147.570 40.750 147.850 ;
        RECT 40.990 147.570 41.270 147.850 ;
        RECT 38.470 145.370 38.750 145.650 ;
        RECT 38.990 145.370 39.270 145.650 ;
        RECT 40.470 144.930 40.750 145.210 ;
        RECT 40.990 144.930 41.270 145.210 ;
        RECT 44.430 144.930 44.710 145.210 ;
        RECT 44.950 144.930 45.230 145.210 ;
        RECT 40.470 143.170 40.750 143.450 ;
        RECT 40.990 143.170 41.270 143.450 ;
        RECT 44.430 143.170 44.710 143.450 ;
        RECT 44.950 143.170 45.230 143.450 ;
        RECT 44.430 142.290 44.710 142.570 ;
        RECT 44.950 142.290 45.230 142.570 ;
        RECT 40.470 141.410 40.750 141.690 ;
        RECT 40.990 141.410 41.270 141.690 ;
        RECT 40.470 140.530 40.750 140.810 ;
        RECT 40.990 140.530 41.270 140.810 ;
        RECT 38.470 140.090 38.750 140.370 ;
        RECT 38.990 140.090 39.270 140.370 ;
        RECT 40.470 137.890 40.750 138.170 ;
        RECT 40.990 137.890 41.270 138.170 ;
        RECT 44.430 137.890 44.710 138.170 ;
        RECT 44.950 137.890 45.230 138.170 ;
        RECT 44.430 137.010 44.710 137.290 ;
        RECT 44.950 137.010 45.230 137.290 ;
        RECT 38.310 136.570 38.590 136.850 ;
        RECT 38.830 136.570 39.110 136.850 ;
        RECT 40.470 135.250 40.750 135.530 ;
        RECT 40.990 135.250 41.270 135.530 ;
        RECT 44.430 135.250 44.710 135.530 ;
        RECT 44.950 135.250 45.230 135.530 ;
        RECT 28.030 134.370 28.310 134.650 ;
        RECT 28.550 134.370 28.830 134.650 ;
        RECT 31.990 134.370 32.270 134.650 ;
        RECT 32.510 134.370 32.790 134.650 ;
        RECT 65.670 187.170 65.950 187.450 ;
        RECT 66.190 187.170 66.470 187.450 ;
        RECT 69.630 187.170 69.910 187.450 ;
        RECT 70.150 187.170 70.430 187.450 ;
        RECT 53.230 186.290 53.510 186.570 ;
        RECT 53.750 186.290 54.030 186.570 ;
        RECT 57.190 186.290 57.470 186.570 ;
        RECT 57.710 186.290 57.990 186.570 ;
        RECT 53.070 185.410 53.350 185.690 ;
        RECT 53.590 185.410 53.870 185.690 ;
        RECT 53.230 184.530 53.510 184.810 ;
        RECT 53.750 184.530 54.030 184.810 ;
        RECT 57.190 184.530 57.470 184.810 ;
        RECT 57.710 184.530 57.990 184.810 ;
        RECT 57.190 183.650 57.470 183.930 ;
        RECT 57.710 183.650 57.990 183.930 ;
        RECT 59.190 183.210 59.470 183.490 ;
        RECT 59.710 183.210 59.990 183.490 ;
        RECT 53.230 181.890 53.510 182.170 ;
        RECT 53.750 181.890 54.030 182.170 ;
        RECT 57.190 181.890 57.470 182.170 ;
        RECT 57.710 181.890 57.990 182.170 ;
        RECT 53.230 180.130 53.510 180.410 ;
        RECT 53.750 180.130 54.030 180.410 ;
        RECT 57.190 180.130 57.470 180.410 ;
        RECT 57.710 180.130 57.990 180.410 ;
        RECT 53.230 179.250 53.510 179.530 ;
        RECT 53.750 179.250 54.030 179.530 ;
        RECT 59.350 178.810 59.630 179.090 ;
        RECT 59.870 178.810 60.150 179.090 ;
        RECT 53.230 177.490 53.510 177.770 ;
        RECT 53.750 177.490 54.030 177.770 ;
        RECT 57.190 177.490 57.470 177.770 ;
        RECT 57.710 177.490 57.990 177.770 ;
        RECT 57.030 176.610 57.310 176.890 ;
        RECT 57.550 176.610 57.830 176.890 ;
        RECT 53.230 175.730 53.510 176.010 ;
        RECT 53.750 175.730 54.030 176.010 ;
        RECT 57.190 175.730 57.470 176.010 ;
        RECT 57.710 175.730 57.990 176.010 ;
        RECT 51.070 174.410 51.350 174.690 ;
        RECT 51.590 174.410 51.870 174.690 ;
        RECT 53.230 173.970 53.510 174.250 ;
        RECT 53.750 173.970 54.030 174.250 ;
        RECT 57.190 173.970 57.470 174.250 ;
        RECT 57.710 173.970 57.990 174.250 ;
        RECT 57.190 173.090 57.470 173.370 ;
        RECT 57.710 173.090 57.990 173.370 ;
        RECT 51.070 171.770 51.350 172.050 ;
        RECT 51.590 171.770 51.870 172.050 ;
        RECT 53.230 171.330 53.510 171.610 ;
        RECT 53.750 171.330 54.030 171.610 ;
        RECT 57.190 171.330 57.470 171.610 ;
        RECT 57.710 171.330 57.990 171.610 ;
        RECT 59.190 170.890 59.470 171.170 ;
        RECT 59.710 170.890 59.990 171.170 ;
        RECT 57.190 169.570 57.470 169.850 ;
        RECT 57.710 169.570 57.990 169.850 ;
        RECT 53.230 168.690 53.510 168.970 ;
        RECT 53.750 168.690 54.030 168.970 ;
        RECT 57.190 168.690 57.470 168.970 ;
        RECT 57.710 168.690 57.990 168.970 ;
        RECT 53.230 166.930 53.510 167.210 ;
        RECT 53.750 166.930 54.030 167.210 ;
        RECT 54.790 166.310 55.070 166.590 ;
        RECT 57.190 166.930 57.470 167.210 ;
        RECT 57.710 166.930 57.990 167.210 ;
        RECT 54.790 165.790 55.070 166.070 ;
        RECT 53.230 165.170 53.510 165.450 ;
        RECT 53.750 165.170 54.030 165.450 ;
        RECT 57.190 165.170 57.470 165.450 ;
        RECT 57.710 165.170 57.990 165.450 ;
        RECT 53.230 164.290 53.510 164.570 ;
        RECT 53.750 164.290 54.030 164.570 ;
        RECT 57.190 164.290 57.470 164.570 ;
        RECT 57.710 164.290 57.990 164.570 ;
        RECT 53.230 162.530 53.510 162.810 ;
        RECT 53.750 162.530 54.030 162.810 ;
        RECT 55.575 161.910 55.855 162.190 ;
        RECT 57.190 162.530 57.470 162.810 ;
        RECT 57.710 162.530 57.990 162.810 ;
        RECT 55.575 161.390 55.855 161.670 ;
        RECT 59.350 161.210 59.630 161.490 ;
        RECT 59.870 161.210 60.150 161.490 ;
        RECT 53.230 160.770 53.510 161.050 ;
        RECT 53.750 160.770 54.030 161.050 ;
        RECT 57.190 160.770 57.470 161.050 ;
        RECT 57.710 160.770 57.990 161.050 ;
        RECT 53.230 159.890 53.510 160.170 ;
        RECT 53.750 159.890 54.030 160.170 ;
        RECT 57.190 159.890 57.470 160.170 ;
        RECT 57.710 159.890 57.990 160.170 ;
        RECT 53.230 158.130 53.510 158.410 ;
        RECT 53.750 158.130 54.030 158.410 ;
        RECT 57.190 158.130 57.470 158.410 ;
        RECT 57.710 158.130 57.990 158.410 ;
        RECT 53.230 157.250 53.510 157.530 ;
        RECT 53.750 157.250 54.030 157.530 ;
        RECT 56.290 157.510 56.570 157.790 ;
        RECT 56.290 156.990 56.570 157.270 ;
        RECT 59.190 156.810 59.470 157.090 ;
        RECT 59.710 156.810 59.990 157.090 ;
        RECT 53.230 156.370 53.510 156.650 ;
        RECT 53.750 156.370 54.030 156.650 ;
        RECT 57.190 156.370 57.470 156.650 ;
        RECT 57.710 156.370 57.990 156.650 ;
        RECT 53.230 155.490 53.510 155.770 ;
        RECT 53.750 155.490 54.030 155.770 ;
        RECT 57.190 155.490 57.470 155.770 ;
        RECT 57.710 155.490 57.990 155.770 ;
        RECT 53.230 153.730 53.510 154.010 ;
        RECT 53.750 153.730 54.030 154.010 ;
        RECT 57.190 153.730 57.470 154.010 ;
        RECT 57.710 153.730 57.990 154.010 ;
        RECT 53.230 151.970 53.510 152.250 ;
        RECT 53.750 151.970 54.030 152.250 ;
        RECT 57.190 151.970 57.470 152.250 ;
        RECT 57.710 151.970 57.990 152.250 ;
        RECT 50.910 150.650 51.190 150.930 ;
        RECT 51.430 150.650 51.710 150.930 ;
        RECT 59.350 150.650 59.630 150.930 ;
        RECT 59.870 150.650 60.150 150.930 ;
        RECT 53.230 148.450 53.510 148.730 ;
        RECT 53.750 148.450 54.030 148.730 ;
        RECT 57.190 148.450 57.470 148.730 ;
        RECT 57.710 148.450 57.990 148.730 ;
        RECT 57.190 147.570 57.470 147.850 ;
        RECT 57.710 147.570 57.990 147.850 ;
        RECT 59.190 148.890 59.470 149.170 ;
        RECT 59.710 148.890 59.990 149.170 ;
        RECT 59.350 147.130 59.630 147.410 ;
        RECT 59.870 147.130 60.150 147.410 ;
        RECT 53.230 144.930 53.510 145.210 ;
        RECT 53.750 144.930 54.030 145.210 ;
        RECT 57.190 144.930 57.470 145.210 ;
        RECT 57.710 144.930 57.990 145.210 ;
        RECT 59.190 145.370 59.470 145.650 ;
        RECT 59.710 145.370 59.990 145.650 ;
        RECT 53.230 143.170 53.510 143.450 ;
        RECT 53.750 143.170 54.030 143.450 ;
        RECT 57.190 143.170 57.470 143.450 ;
        RECT 57.710 143.170 57.990 143.450 ;
        RECT 53.230 142.290 53.510 142.570 ;
        RECT 53.750 142.290 54.030 142.570 ;
        RECT 57.190 141.410 57.470 141.690 ;
        RECT 57.710 141.410 57.990 141.690 ;
        RECT 57.190 140.530 57.470 140.810 ;
        RECT 57.710 140.530 57.990 140.810 ;
        RECT 59.190 140.090 59.470 140.370 ;
        RECT 59.710 140.090 59.990 140.370 ;
        RECT 53.230 137.890 53.510 138.170 ;
        RECT 53.750 137.890 54.030 138.170 ;
        RECT 57.190 137.890 57.470 138.170 ;
        RECT 57.710 137.890 57.990 138.170 ;
        RECT 53.230 137.010 53.510 137.290 ;
        RECT 53.750 137.010 54.030 137.290 ;
        RECT 59.350 136.570 59.630 136.850 ;
        RECT 59.870 136.570 60.150 136.850 ;
        RECT 53.230 135.250 53.510 135.530 ;
        RECT 53.750 135.250 54.030 135.530 ;
        RECT 57.190 135.250 57.470 135.530 ;
        RECT 57.710 135.250 57.990 135.530 ;
        RECT 40.470 134.370 40.750 134.650 ;
        RECT 40.990 134.370 41.270 134.650 ;
        RECT 44.430 134.370 44.710 134.650 ;
        RECT 44.950 134.370 45.230 134.650 ;
        RECT 78.430 187.170 78.710 187.450 ;
        RECT 78.950 187.170 79.230 187.450 ;
        RECT 82.390 187.170 82.670 187.450 ;
        RECT 82.910 187.170 83.190 187.450 ;
        RECT 65.670 186.290 65.950 186.570 ;
        RECT 66.190 186.290 66.470 186.570 ;
        RECT 69.630 186.290 69.910 186.570 ;
        RECT 70.150 186.290 70.430 186.570 ;
        RECT 69.630 185.580 69.910 185.860 ;
        RECT 70.150 185.580 70.430 185.860 ;
        RECT 63.510 183.210 63.790 183.490 ;
        RECT 64.030 183.210 64.310 183.490 ;
        RECT 65.670 184.530 65.950 184.810 ;
        RECT 66.190 184.530 66.470 184.810 ;
        RECT 69.630 184.530 69.910 184.810 ;
        RECT 70.150 184.530 70.430 184.810 ;
        RECT 65.670 183.650 65.950 183.930 ;
        RECT 66.190 183.650 66.470 183.930 ;
        RECT 65.670 181.890 65.950 182.170 ;
        RECT 66.190 181.890 66.470 182.170 ;
        RECT 69.630 181.890 69.910 182.170 ;
        RECT 70.150 181.890 70.430 182.170 ;
        RECT 65.670 180.130 65.950 180.410 ;
        RECT 66.190 180.130 66.470 180.410 ;
        RECT 69.630 180.130 69.910 180.410 ;
        RECT 70.150 180.130 70.430 180.410 ;
        RECT 69.630 179.250 69.910 179.530 ;
        RECT 70.150 179.250 70.430 179.530 ;
        RECT 63.510 178.810 63.790 179.090 ;
        RECT 64.030 178.810 64.310 179.090 ;
        RECT 65.670 177.490 65.950 177.770 ;
        RECT 66.190 177.490 66.470 177.770 ;
        RECT 69.630 177.490 69.910 177.770 ;
        RECT 70.150 177.490 70.430 177.770 ;
        RECT 65.670 176.610 65.950 176.890 ;
        RECT 66.190 176.610 66.470 176.890 ;
        RECT 65.670 175.730 65.950 176.010 ;
        RECT 66.190 175.730 66.470 176.010 ;
        RECT 69.630 175.730 69.910 176.010 ;
        RECT 70.150 175.730 70.430 176.010 ;
        RECT 71.790 174.410 72.070 174.690 ;
        RECT 72.310 174.410 72.590 174.690 ;
        RECT 65.670 173.970 65.950 174.250 ;
        RECT 66.190 173.970 66.470 174.250 ;
        RECT 69.630 173.970 69.910 174.250 ;
        RECT 70.150 173.970 70.430 174.250 ;
        RECT 65.670 173.090 65.950 173.370 ;
        RECT 66.190 173.090 66.470 173.370 ;
        RECT 65.670 171.330 65.950 171.610 ;
        RECT 66.190 171.330 66.470 171.610 ;
        RECT 63.510 170.890 63.790 171.170 ;
        RECT 64.030 170.890 64.310 171.170 ;
        RECT 71.790 171.770 72.070 172.050 ;
        RECT 72.310 171.770 72.590 172.050 ;
        RECT 69.630 171.330 69.910 171.610 ;
        RECT 70.150 171.330 70.430 171.610 ;
        RECT 65.670 169.570 65.950 169.850 ;
        RECT 66.190 169.570 66.470 169.850 ;
        RECT 65.670 168.690 65.950 168.970 ;
        RECT 66.190 168.690 66.470 168.970 ;
        RECT 69.630 168.690 69.910 168.970 ;
        RECT 70.150 168.690 70.430 168.970 ;
        RECT 65.670 166.930 65.950 167.210 ;
        RECT 66.190 166.930 66.470 167.210 ;
        RECT 69.630 166.930 69.910 167.210 ;
        RECT 70.150 166.930 70.430 167.210 ;
        RECT 68.590 166.310 68.870 166.590 ;
        RECT 68.590 165.790 68.870 166.070 ;
        RECT 65.670 165.170 65.950 165.450 ;
        RECT 66.190 165.170 66.470 165.450 ;
        RECT 69.630 165.170 69.910 165.450 ;
        RECT 70.150 165.170 70.430 165.450 ;
        RECT 65.670 164.290 65.950 164.570 ;
        RECT 66.190 164.290 66.470 164.570 ;
        RECT 69.630 164.290 69.910 164.570 ;
        RECT 70.150 164.290 70.430 164.570 ;
        RECT 65.670 162.530 65.950 162.810 ;
        RECT 66.190 162.530 66.470 162.810 ;
        RECT 69.630 162.530 69.910 162.810 ;
        RECT 70.150 162.530 70.430 162.810 ;
        RECT 67.805 161.910 68.085 162.190 ;
        RECT 63.510 161.210 63.790 161.490 ;
        RECT 64.030 161.210 64.310 161.490 ;
        RECT 67.805 161.390 68.085 161.670 ;
        RECT 65.670 160.770 65.950 161.050 ;
        RECT 66.190 160.770 66.470 161.050 ;
        RECT 69.630 160.770 69.910 161.050 ;
        RECT 70.150 160.770 70.430 161.050 ;
        RECT 65.670 159.890 65.950 160.170 ;
        RECT 66.190 159.890 66.470 160.170 ;
        RECT 69.630 159.890 69.910 160.170 ;
        RECT 70.150 159.890 70.430 160.170 ;
        RECT 65.670 158.130 65.950 158.410 ;
        RECT 66.190 158.130 66.470 158.410 ;
        RECT 69.630 158.130 69.910 158.410 ;
        RECT 70.150 158.130 70.430 158.410 ;
        RECT 67.090 157.510 67.370 157.790 ;
        RECT 63.670 156.810 63.950 157.090 ;
        RECT 64.190 156.810 64.470 157.090 ;
        RECT 67.090 156.990 67.370 157.270 ;
        RECT 69.630 157.250 69.910 157.530 ;
        RECT 70.150 157.250 70.430 157.530 ;
        RECT 65.670 156.370 65.950 156.650 ;
        RECT 66.190 156.370 66.470 156.650 ;
        RECT 69.630 156.370 69.910 156.650 ;
        RECT 70.150 156.370 70.430 156.650 ;
        RECT 65.670 155.490 65.950 155.770 ;
        RECT 66.190 155.490 66.470 155.770 ;
        RECT 69.630 155.490 69.910 155.770 ;
        RECT 70.150 155.490 70.430 155.770 ;
        RECT 65.670 153.730 65.950 154.010 ;
        RECT 66.190 153.730 66.470 154.010 ;
        RECT 69.630 153.730 69.910 154.010 ;
        RECT 70.150 153.730 70.430 154.010 ;
        RECT 65.670 151.970 65.950 152.250 ;
        RECT 66.190 151.970 66.470 152.250 ;
        RECT 69.630 151.970 69.910 152.250 ;
        RECT 70.150 151.970 70.430 152.250 ;
        RECT 63.510 150.650 63.790 150.930 ;
        RECT 64.030 150.650 64.310 150.930 ;
        RECT 71.790 150.650 72.070 150.930 ;
        RECT 72.310 150.650 72.590 150.930 ;
        RECT 63.510 148.890 63.790 149.170 ;
        RECT 64.030 148.890 64.310 149.170 ;
        RECT 63.510 147.130 63.790 147.410 ;
        RECT 64.030 147.130 64.310 147.410 ;
        RECT 65.670 148.450 65.950 148.730 ;
        RECT 66.190 148.450 66.470 148.730 ;
        RECT 69.630 148.450 69.910 148.730 ;
        RECT 70.150 148.450 70.430 148.730 ;
        RECT 65.670 147.570 65.950 147.850 ;
        RECT 66.190 147.570 66.470 147.850 ;
        RECT 63.670 145.370 63.950 145.650 ;
        RECT 64.190 145.370 64.470 145.650 ;
        RECT 65.670 144.930 65.950 145.210 ;
        RECT 66.190 144.930 66.470 145.210 ;
        RECT 69.630 144.930 69.910 145.210 ;
        RECT 70.150 144.930 70.430 145.210 ;
        RECT 65.670 143.170 65.950 143.450 ;
        RECT 66.190 143.170 66.470 143.450 ;
        RECT 69.630 143.170 69.910 143.450 ;
        RECT 70.150 143.170 70.430 143.450 ;
        RECT 69.630 142.290 69.910 142.570 ;
        RECT 70.150 142.290 70.430 142.570 ;
        RECT 65.670 141.410 65.950 141.690 ;
        RECT 66.190 141.410 66.470 141.690 ;
        RECT 65.670 140.530 65.950 140.810 ;
        RECT 66.190 140.530 66.470 140.810 ;
        RECT 63.670 140.090 63.950 140.370 ;
        RECT 64.190 140.090 64.470 140.370 ;
        RECT 65.670 137.890 65.950 138.170 ;
        RECT 66.190 137.890 66.470 138.170 ;
        RECT 69.630 137.890 69.910 138.170 ;
        RECT 70.150 137.890 70.430 138.170 ;
        RECT 69.630 137.010 69.910 137.290 ;
        RECT 70.150 137.010 70.430 137.290 ;
        RECT 63.510 136.570 63.790 136.850 ;
        RECT 64.030 136.570 64.310 136.850 ;
        RECT 65.670 135.250 65.950 135.530 ;
        RECT 66.190 135.250 66.470 135.530 ;
        RECT 69.630 135.250 69.910 135.530 ;
        RECT 70.150 135.250 70.430 135.530 ;
        RECT 53.230 134.370 53.510 134.650 ;
        RECT 53.750 134.370 54.030 134.650 ;
        RECT 57.190 134.370 57.470 134.650 ;
        RECT 57.710 134.370 57.990 134.650 ;
        RECT 90.870 187.170 91.150 187.450 ;
        RECT 91.390 187.170 91.670 187.450 ;
        RECT 94.830 187.170 95.110 187.450 ;
        RECT 95.350 187.170 95.630 187.450 ;
        RECT 78.430 186.290 78.710 186.570 ;
        RECT 78.950 186.290 79.230 186.570 ;
        RECT 82.390 186.290 82.670 186.570 ;
        RECT 82.910 186.290 83.190 186.570 ;
        RECT 78.270 185.410 78.550 185.690 ;
        RECT 78.790 185.410 79.070 185.690 ;
        RECT 78.430 184.530 78.710 184.810 ;
        RECT 78.950 184.530 79.230 184.810 ;
        RECT 82.390 184.530 82.670 184.810 ;
        RECT 82.910 184.530 83.190 184.810 ;
        RECT 82.390 183.650 82.670 183.930 ;
        RECT 82.910 183.650 83.190 183.930 ;
        RECT 84.390 183.210 84.670 183.490 ;
        RECT 84.910 183.210 85.190 183.490 ;
        RECT 78.430 181.890 78.710 182.170 ;
        RECT 78.950 181.890 79.230 182.170 ;
        RECT 82.390 181.890 82.670 182.170 ;
        RECT 82.910 181.890 83.190 182.170 ;
        RECT 78.430 180.130 78.710 180.410 ;
        RECT 78.950 180.130 79.230 180.410 ;
        RECT 82.390 180.130 82.670 180.410 ;
        RECT 82.910 180.130 83.190 180.410 ;
        RECT 78.430 179.250 78.710 179.530 ;
        RECT 78.950 179.250 79.230 179.530 ;
        RECT 84.550 178.810 84.830 179.090 ;
        RECT 85.070 178.810 85.350 179.090 ;
        RECT 78.430 177.490 78.710 177.770 ;
        RECT 78.950 177.490 79.230 177.770 ;
        RECT 82.390 177.490 82.670 177.770 ;
        RECT 82.910 177.490 83.190 177.770 ;
        RECT 82.230 176.610 82.510 176.890 ;
        RECT 82.750 176.610 83.030 176.890 ;
        RECT 78.430 175.730 78.710 176.010 ;
        RECT 78.950 175.730 79.230 176.010 ;
        RECT 82.390 175.730 82.670 176.010 ;
        RECT 82.910 175.730 83.190 176.010 ;
        RECT 76.270 174.410 76.550 174.690 ;
        RECT 76.790 174.410 77.070 174.690 ;
        RECT 78.430 173.970 78.710 174.250 ;
        RECT 78.950 173.970 79.230 174.250 ;
        RECT 82.390 173.970 82.670 174.250 ;
        RECT 82.910 173.970 83.190 174.250 ;
        RECT 82.390 173.090 82.670 173.370 ;
        RECT 82.910 173.090 83.190 173.370 ;
        RECT 76.270 171.770 76.550 172.050 ;
        RECT 76.790 171.770 77.070 172.050 ;
        RECT 78.430 171.330 78.710 171.610 ;
        RECT 78.950 171.330 79.230 171.610 ;
        RECT 82.390 171.330 82.670 171.610 ;
        RECT 82.910 171.330 83.190 171.610 ;
        RECT 84.390 170.890 84.670 171.170 ;
        RECT 84.910 170.890 85.190 171.170 ;
        RECT 82.390 169.570 82.670 169.850 ;
        RECT 82.910 169.570 83.190 169.850 ;
        RECT 78.430 168.690 78.710 168.970 ;
        RECT 78.950 168.690 79.230 168.970 ;
        RECT 82.390 168.690 82.670 168.970 ;
        RECT 82.910 168.690 83.190 168.970 ;
        RECT 78.430 166.930 78.710 167.210 ;
        RECT 78.950 166.930 79.230 167.210 ;
        RECT 79.990 166.310 80.270 166.590 ;
        RECT 82.390 166.930 82.670 167.210 ;
        RECT 82.910 166.930 83.190 167.210 ;
        RECT 79.990 165.790 80.270 166.070 ;
        RECT 78.430 165.170 78.710 165.450 ;
        RECT 78.950 165.170 79.230 165.450 ;
        RECT 82.390 165.170 82.670 165.450 ;
        RECT 82.910 165.170 83.190 165.450 ;
        RECT 78.430 164.290 78.710 164.570 ;
        RECT 78.950 164.290 79.230 164.570 ;
        RECT 82.390 164.290 82.670 164.570 ;
        RECT 82.910 164.290 83.190 164.570 ;
        RECT 78.430 162.530 78.710 162.810 ;
        RECT 78.950 162.530 79.230 162.810 ;
        RECT 80.775 161.910 81.055 162.190 ;
        RECT 82.390 162.530 82.670 162.810 ;
        RECT 82.910 162.530 83.190 162.810 ;
        RECT 80.775 161.390 81.055 161.670 ;
        RECT 84.550 161.210 84.830 161.490 ;
        RECT 85.070 161.210 85.350 161.490 ;
        RECT 78.430 160.770 78.710 161.050 ;
        RECT 78.950 160.770 79.230 161.050 ;
        RECT 82.390 160.770 82.670 161.050 ;
        RECT 82.910 160.770 83.190 161.050 ;
        RECT 78.430 159.890 78.710 160.170 ;
        RECT 78.950 159.890 79.230 160.170 ;
        RECT 82.390 159.890 82.670 160.170 ;
        RECT 82.910 159.890 83.190 160.170 ;
        RECT 78.430 158.130 78.710 158.410 ;
        RECT 78.950 158.130 79.230 158.410 ;
        RECT 82.390 158.130 82.670 158.410 ;
        RECT 82.910 158.130 83.190 158.410 ;
        RECT 78.430 157.250 78.710 157.530 ;
        RECT 78.950 157.250 79.230 157.530 ;
        RECT 81.490 157.510 81.770 157.790 ;
        RECT 81.490 156.990 81.770 157.270 ;
        RECT 84.390 156.810 84.670 157.090 ;
        RECT 84.910 156.810 85.190 157.090 ;
        RECT 78.430 156.370 78.710 156.650 ;
        RECT 78.950 156.370 79.230 156.650 ;
        RECT 82.390 156.370 82.670 156.650 ;
        RECT 82.910 156.370 83.190 156.650 ;
        RECT 78.430 155.490 78.710 155.770 ;
        RECT 78.950 155.490 79.230 155.770 ;
        RECT 82.390 155.490 82.670 155.770 ;
        RECT 82.910 155.490 83.190 155.770 ;
        RECT 78.430 153.730 78.710 154.010 ;
        RECT 78.950 153.730 79.230 154.010 ;
        RECT 82.390 153.730 82.670 154.010 ;
        RECT 82.910 153.730 83.190 154.010 ;
        RECT 78.430 151.970 78.710 152.250 ;
        RECT 78.950 151.970 79.230 152.250 ;
        RECT 82.390 151.970 82.670 152.250 ;
        RECT 82.910 151.970 83.190 152.250 ;
        RECT 76.110 150.650 76.390 150.930 ;
        RECT 76.630 150.650 76.910 150.930 ;
        RECT 84.550 150.650 84.830 150.930 ;
        RECT 85.070 150.650 85.350 150.930 ;
        RECT 78.430 148.450 78.710 148.730 ;
        RECT 78.950 148.450 79.230 148.730 ;
        RECT 82.390 148.450 82.670 148.730 ;
        RECT 82.910 148.450 83.190 148.730 ;
        RECT 82.390 147.570 82.670 147.850 ;
        RECT 82.910 147.570 83.190 147.850 ;
        RECT 84.390 148.890 84.670 149.170 ;
        RECT 84.910 148.890 85.190 149.170 ;
        RECT 84.550 147.130 84.830 147.410 ;
        RECT 85.070 147.130 85.350 147.410 ;
        RECT 78.430 144.930 78.710 145.210 ;
        RECT 78.950 144.930 79.230 145.210 ;
        RECT 82.390 144.930 82.670 145.210 ;
        RECT 82.910 144.930 83.190 145.210 ;
        RECT 84.390 145.370 84.670 145.650 ;
        RECT 84.910 145.370 85.190 145.650 ;
        RECT 78.430 143.170 78.710 143.450 ;
        RECT 78.950 143.170 79.230 143.450 ;
        RECT 82.390 143.170 82.670 143.450 ;
        RECT 82.910 143.170 83.190 143.450 ;
        RECT 78.430 142.290 78.710 142.570 ;
        RECT 78.950 142.290 79.230 142.570 ;
        RECT 82.390 141.410 82.670 141.690 ;
        RECT 82.910 141.410 83.190 141.690 ;
        RECT 82.390 140.530 82.670 140.810 ;
        RECT 82.910 140.530 83.190 140.810 ;
        RECT 84.390 140.090 84.670 140.370 ;
        RECT 84.910 140.090 85.190 140.370 ;
        RECT 78.430 137.890 78.710 138.170 ;
        RECT 78.950 137.890 79.230 138.170 ;
        RECT 82.390 137.890 82.670 138.170 ;
        RECT 82.910 137.890 83.190 138.170 ;
        RECT 78.430 137.010 78.710 137.290 ;
        RECT 78.950 137.010 79.230 137.290 ;
        RECT 84.550 136.570 84.830 136.850 ;
        RECT 85.070 136.570 85.350 136.850 ;
        RECT 78.430 135.250 78.710 135.530 ;
        RECT 78.950 135.250 79.230 135.530 ;
        RECT 82.390 135.250 82.670 135.530 ;
        RECT 82.910 135.250 83.190 135.530 ;
        RECT 65.670 134.370 65.950 134.650 ;
        RECT 66.190 134.370 66.470 134.650 ;
        RECT 69.630 134.370 69.910 134.650 ;
        RECT 70.150 134.370 70.430 134.650 ;
        RECT 103.630 187.170 103.910 187.450 ;
        RECT 104.150 187.170 104.430 187.450 ;
        RECT 107.590 187.170 107.870 187.450 ;
        RECT 108.110 187.170 108.390 187.450 ;
        RECT 90.870 186.290 91.150 186.570 ;
        RECT 91.390 186.290 91.670 186.570 ;
        RECT 94.830 186.290 95.110 186.570 ;
        RECT 95.350 186.290 95.630 186.570 ;
        RECT 94.830 185.580 95.110 185.860 ;
        RECT 95.350 185.580 95.630 185.860 ;
        RECT 88.710 183.210 88.990 183.490 ;
        RECT 89.230 183.210 89.510 183.490 ;
        RECT 90.870 184.530 91.150 184.810 ;
        RECT 91.390 184.530 91.670 184.810 ;
        RECT 94.830 184.530 95.110 184.810 ;
        RECT 95.350 184.530 95.630 184.810 ;
        RECT 90.870 183.650 91.150 183.930 ;
        RECT 91.390 183.650 91.670 183.930 ;
        RECT 90.870 181.890 91.150 182.170 ;
        RECT 91.390 181.890 91.670 182.170 ;
        RECT 94.830 181.890 95.110 182.170 ;
        RECT 95.350 181.890 95.630 182.170 ;
        RECT 90.870 180.130 91.150 180.410 ;
        RECT 91.390 180.130 91.670 180.410 ;
        RECT 94.830 180.130 95.110 180.410 ;
        RECT 95.350 180.130 95.630 180.410 ;
        RECT 94.830 179.250 95.110 179.530 ;
        RECT 95.350 179.250 95.630 179.530 ;
        RECT 88.710 178.810 88.990 179.090 ;
        RECT 89.230 178.810 89.510 179.090 ;
        RECT 90.870 177.490 91.150 177.770 ;
        RECT 91.390 177.490 91.670 177.770 ;
        RECT 94.830 177.490 95.110 177.770 ;
        RECT 95.350 177.490 95.630 177.770 ;
        RECT 90.870 176.610 91.150 176.890 ;
        RECT 91.390 176.610 91.670 176.890 ;
        RECT 90.870 175.730 91.150 176.010 ;
        RECT 91.390 175.730 91.670 176.010 ;
        RECT 94.830 175.730 95.110 176.010 ;
        RECT 95.350 175.730 95.630 176.010 ;
        RECT 96.990 174.410 97.270 174.690 ;
        RECT 97.510 174.410 97.790 174.690 ;
        RECT 90.870 173.970 91.150 174.250 ;
        RECT 91.390 173.970 91.670 174.250 ;
        RECT 94.830 173.970 95.110 174.250 ;
        RECT 95.350 173.970 95.630 174.250 ;
        RECT 90.870 173.090 91.150 173.370 ;
        RECT 91.390 173.090 91.670 173.370 ;
        RECT 90.870 171.330 91.150 171.610 ;
        RECT 91.390 171.330 91.670 171.610 ;
        RECT 88.710 170.890 88.990 171.170 ;
        RECT 89.230 170.890 89.510 171.170 ;
        RECT 96.990 171.770 97.270 172.050 ;
        RECT 97.510 171.770 97.790 172.050 ;
        RECT 94.830 171.330 95.110 171.610 ;
        RECT 95.350 171.330 95.630 171.610 ;
        RECT 90.870 169.570 91.150 169.850 ;
        RECT 91.390 169.570 91.670 169.850 ;
        RECT 90.870 168.690 91.150 168.970 ;
        RECT 91.390 168.690 91.670 168.970 ;
        RECT 94.830 168.690 95.110 168.970 ;
        RECT 95.350 168.690 95.630 168.970 ;
        RECT 90.870 166.930 91.150 167.210 ;
        RECT 91.390 166.930 91.670 167.210 ;
        RECT 94.830 166.930 95.110 167.210 ;
        RECT 95.350 166.930 95.630 167.210 ;
        RECT 93.790 166.310 94.070 166.590 ;
        RECT 93.790 165.790 94.070 166.070 ;
        RECT 90.870 165.170 91.150 165.450 ;
        RECT 91.390 165.170 91.670 165.450 ;
        RECT 94.830 165.170 95.110 165.450 ;
        RECT 95.350 165.170 95.630 165.450 ;
        RECT 90.870 164.290 91.150 164.570 ;
        RECT 91.390 164.290 91.670 164.570 ;
        RECT 94.830 164.290 95.110 164.570 ;
        RECT 95.350 164.290 95.630 164.570 ;
        RECT 90.870 162.530 91.150 162.810 ;
        RECT 91.390 162.530 91.670 162.810 ;
        RECT 94.830 162.530 95.110 162.810 ;
        RECT 95.350 162.530 95.630 162.810 ;
        RECT 93.005 161.910 93.285 162.190 ;
        RECT 88.710 161.210 88.990 161.490 ;
        RECT 89.230 161.210 89.510 161.490 ;
        RECT 93.005 161.390 93.285 161.670 ;
        RECT 90.870 160.770 91.150 161.050 ;
        RECT 91.390 160.770 91.670 161.050 ;
        RECT 94.830 160.770 95.110 161.050 ;
        RECT 95.350 160.770 95.630 161.050 ;
        RECT 90.870 159.890 91.150 160.170 ;
        RECT 91.390 159.890 91.670 160.170 ;
        RECT 94.830 159.890 95.110 160.170 ;
        RECT 95.350 159.890 95.630 160.170 ;
        RECT 90.870 158.130 91.150 158.410 ;
        RECT 91.390 158.130 91.670 158.410 ;
        RECT 94.830 158.130 95.110 158.410 ;
        RECT 95.350 158.130 95.630 158.410 ;
        RECT 92.290 157.510 92.570 157.790 ;
        RECT 88.870 156.810 89.150 157.090 ;
        RECT 89.390 156.810 89.670 157.090 ;
        RECT 92.290 156.990 92.570 157.270 ;
        RECT 94.830 157.250 95.110 157.530 ;
        RECT 95.350 157.250 95.630 157.530 ;
        RECT 90.870 156.370 91.150 156.650 ;
        RECT 91.390 156.370 91.670 156.650 ;
        RECT 94.830 156.370 95.110 156.650 ;
        RECT 95.350 156.370 95.630 156.650 ;
        RECT 90.870 155.490 91.150 155.770 ;
        RECT 91.390 155.490 91.670 155.770 ;
        RECT 94.830 155.490 95.110 155.770 ;
        RECT 95.350 155.490 95.630 155.770 ;
        RECT 90.870 153.730 91.150 154.010 ;
        RECT 91.390 153.730 91.670 154.010 ;
        RECT 94.830 153.730 95.110 154.010 ;
        RECT 95.350 153.730 95.630 154.010 ;
        RECT 90.870 151.970 91.150 152.250 ;
        RECT 91.390 151.970 91.670 152.250 ;
        RECT 94.830 151.970 95.110 152.250 ;
        RECT 95.350 151.970 95.630 152.250 ;
        RECT 88.710 150.650 88.990 150.930 ;
        RECT 89.230 150.650 89.510 150.930 ;
        RECT 96.990 150.650 97.270 150.930 ;
        RECT 97.510 150.650 97.790 150.930 ;
        RECT 88.710 148.890 88.990 149.170 ;
        RECT 89.230 148.890 89.510 149.170 ;
        RECT 88.710 147.130 88.990 147.410 ;
        RECT 89.230 147.130 89.510 147.410 ;
        RECT 90.870 148.450 91.150 148.730 ;
        RECT 91.390 148.450 91.670 148.730 ;
        RECT 94.830 148.450 95.110 148.730 ;
        RECT 95.350 148.450 95.630 148.730 ;
        RECT 90.870 147.570 91.150 147.850 ;
        RECT 91.390 147.570 91.670 147.850 ;
        RECT 88.870 145.370 89.150 145.650 ;
        RECT 89.390 145.370 89.670 145.650 ;
        RECT 90.870 144.930 91.150 145.210 ;
        RECT 91.390 144.930 91.670 145.210 ;
        RECT 94.830 144.930 95.110 145.210 ;
        RECT 95.350 144.930 95.630 145.210 ;
        RECT 90.870 143.170 91.150 143.450 ;
        RECT 91.390 143.170 91.670 143.450 ;
        RECT 94.830 143.170 95.110 143.450 ;
        RECT 95.350 143.170 95.630 143.450 ;
        RECT 94.830 142.290 95.110 142.570 ;
        RECT 95.350 142.290 95.630 142.570 ;
        RECT 90.870 141.410 91.150 141.690 ;
        RECT 91.390 141.410 91.670 141.690 ;
        RECT 90.870 140.530 91.150 140.810 ;
        RECT 91.390 140.530 91.670 140.810 ;
        RECT 88.870 140.090 89.150 140.370 ;
        RECT 89.390 140.090 89.670 140.370 ;
        RECT 90.870 137.890 91.150 138.170 ;
        RECT 91.390 137.890 91.670 138.170 ;
        RECT 94.830 137.890 95.110 138.170 ;
        RECT 95.350 137.890 95.630 138.170 ;
        RECT 94.830 137.010 95.110 137.290 ;
        RECT 95.350 137.010 95.630 137.290 ;
        RECT 88.710 136.570 88.990 136.850 ;
        RECT 89.230 136.570 89.510 136.850 ;
        RECT 90.870 135.250 91.150 135.530 ;
        RECT 91.390 135.250 91.670 135.530 ;
        RECT 94.830 135.250 95.110 135.530 ;
        RECT 95.350 135.250 95.630 135.530 ;
        RECT 78.430 134.370 78.710 134.650 ;
        RECT 78.950 134.370 79.230 134.650 ;
        RECT 82.390 134.370 82.670 134.650 ;
        RECT 82.910 134.370 83.190 134.650 ;
        RECT 103.630 186.290 103.910 186.570 ;
        RECT 104.150 186.290 104.430 186.570 ;
        RECT 107.590 186.290 107.870 186.570 ;
        RECT 108.110 186.290 108.390 186.570 ;
        RECT 103.470 185.410 103.750 185.690 ;
        RECT 103.990 185.410 104.270 185.690 ;
        RECT 103.630 184.530 103.910 184.810 ;
        RECT 104.150 184.530 104.430 184.810 ;
        RECT 107.590 184.530 107.870 184.810 ;
        RECT 108.110 184.530 108.390 184.810 ;
        RECT 107.590 183.650 107.870 183.930 ;
        RECT 108.110 183.650 108.390 183.930 ;
        RECT 109.590 183.210 109.870 183.490 ;
        RECT 110.110 183.210 110.390 183.490 ;
        RECT 116.070 182.770 116.350 183.050 ;
        RECT 116.590 182.770 116.870 183.050 ;
        RECT 120.030 182.770 120.310 183.050 ;
        RECT 120.550 182.770 120.830 183.050 ;
        RECT 103.630 181.890 103.910 182.170 ;
        RECT 104.150 181.890 104.430 182.170 ;
        RECT 107.590 181.890 107.870 182.170 ;
        RECT 108.110 181.890 108.390 182.170 ;
        RECT 103.630 180.130 103.910 180.410 ;
        RECT 104.150 180.130 104.430 180.410 ;
        RECT 107.590 180.130 107.870 180.410 ;
        RECT 108.110 180.130 108.390 180.410 ;
        RECT 103.630 179.250 103.910 179.530 ;
        RECT 104.150 179.250 104.430 179.530 ;
        RECT 109.750 178.810 110.030 179.090 ;
        RECT 110.270 178.810 110.550 179.090 ;
        RECT 103.630 177.490 103.910 177.770 ;
        RECT 104.150 177.490 104.430 177.770 ;
        RECT 107.590 177.490 107.870 177.770 ;
        RECT 108.110 177.490 108.390 177.770 ;
        RECT 107.430 176.610 107.710 176.890 ;
        RECT 107.950 176.610 108.230 176.890 ;
        RECT 103.630 175.730 103.910 176.010 ;
        RECT 104.150 175.730 104.430 176.010 ;
        RECT 107.590 175.730 107.870 176.010 ;
        RECT 108.110 175.730 108.390 176.010 ;
        RECT 101.470 174.410 101.750 174.690 ;
        RECT 101.990 174.410 102.270 174.690 ;
        RECT 103.630 173.970 103.910 174.250 ;
        RECT 104.150 173.970 104.430 174.250 ;
        RECT 107.590 173.970 107.870 174.250 ;
        RECT 108.110 173.970 108.390 174.250 ;
        RECT 107.590 173.090 107.870 173.370 ;
        RECT 108.110 173.090 108.390 173.370 ;
        RECT 101.470 171.770 101.750 172.050 ;
        RECT 101.990 171.770 102.270 172.050 ;
        RECT 103.630 171.330 103.910 171.610 ;
        RECT 104.150 171.330 104.430 171.610 ;
        RECT 109.590 172.650 109.870 172.930 ;
        RECT 110.110 172.650 110.390 172.930 ;
        RECT 107.590 171.330 107.870 171.610 ;
        RECT 108.110 171.330 108.390 171.610 ;
        RECT 109.590 170.890 109.870 171.170 ;
        RECT 110.110 170.890 110.390 171.170 ;
        RECT 107.590 169.570 107.870 169.850 ;
        RECT 108.110 169.570 108.390 169.850 ;
        RECT 103.630 168.690 103.910 168.970 ;
        RECT 104.150 168.690 104.430 168.970 ;
        RECT 107.590 168.690 107.870 168.970 ;
        RECT 108.110 168.690 108.390 168.970 ;
        RECT 103.630 166.930 103.910 167.210 ;
        RECT 104.150 166.930 104.430 167.210 ;
        RECT 105.190 166.310 105.470 166.590 ;
        RECT 107.590 166.930 107.870 167.210 ;
        RECT 108.110 166.930 108.390 167.210 ;
        RECT 105.190 165.790 105.470 166.070 ;
        RECT 103.630 165.170 103.910 165.450 ;
        RECT 104.150 165.170 104.430 165.450 ;
        RECT 107.590 165.170 107.870 165.450 ;
        RECT 108.110 165.170 108.390 165.450 ;
        RECT 103.630 164.290 103.910 164.570 ;
        RECT 104.150 164.290 104.430 164.570 ;
        RECT 107.590 164.290 107.870 164.570 ;
        RECT 108.110 164.290 108.390 164.570 ;
        RECT 103.630 162.530 103.910 162.810 ;
        RECT 104.150 162.530 104.430 162.810 ;
        RECT 105.975 161.910 106.255 162.190 ;
        RECT 107.590 162.530 107.870 162.810 ;
        RECT 108.110 162.530 108.390 162.810 ;
        RECT 105.975 161.390 106.255 161.670 ;
        RECT 109.750 161.210 110.030 161.490 ;
        RECT 110.270 161.210 110.550 161.490 ;
        RECT 103.630 160.770 103.910 161.050 ;
        RECT 104.150 160.770 104.430 161.050 ;
        RECT 107.590 160.770 107.870 161.050 ;
        RECT 108.110 160.770 108.390 161.050 ;
        RECT 103.630 159.890 103.910 160.170 ;
        RECT 104.150 159.890 104.430 160.170 ;
        RECT 107.590 159.890 107.870 160.170 ;
        RECT 108.110 159.890 108.390 160.170 ;
        RECT 103.630 158.130 103.910 158.410 ;
        RECT 104.150 158.130 104.430 158.410 ;
        RECT 107.590 158.130 107.870 158.410 ;
        RECT 108.110 158.130 108.390 158.410 ;
        RECT 103.630 157.250 103.910 157.530 ;
        RECT 104.150 157.250 104.430 157.530 ;
        RECT 106.690 157.510 106.970 157.790 ;
        RECT 106.690 156.990 106.970 157.270 ;
        RECT 109.590 156.810 109.870 157.090 ;
        RECT 110.110 156.810 110.390 157.090 ;
        RECT 103.630 156.370 103.910 156.650 ;
        RECT 104.150 156.370 104.430 156.650 ;
        RECT 107.590 156.370 107.870 156.650 ;
        RECT 108.110 156.370 108.390 156.650 ;
        RECT 103.630 155.490 103.910 155.770 ;
        RECT 104.150 155.490 104.430 155.770 ;
        RECT 107.590 155.490 107.870 155.770 ;
        RECT 108.110 155.490 108.390 155.770 ;
        RECT 103.630 153.730 103.910 154.010 ;
        RECT 104.150 153.730 104.430 154.010 ;
        RECT 107.590 153.730 107.870 154.010 ;
        RECT 108.110 153.730 108.390 154.010 ;
        RECT 103.630 151.970 103.910 152.250 ;
        RECT 104.150 151.970 104.430 152.250 ;
        RECT 107.590 151.970 107.870 152.250 ;
        RECT 108.110 151.970 108.390 152.250 ;
        RECT 101.310 150.650 101.590 150.930 ;
        RECT 101.830 150.650 102.110 150.930 ;
        RECT 109.750 150.650 110.030 150.930 ;
        RECT 110.270 150.650 110.550 150.930 ;
        RECT 103.630 148.450 103.910 148.730 ;
        RECT 104.150 148.450 104.430 148.730 ;
        RECT 107.590 148.450 107.870 148.730 ;
        RECT 108.110 148.450 108.390 148.730 ;
        RECT 107.590 147.570 107.870 147.850 ;
        RECT 108.110 147.570 108.390 147.850 ;
        RECT 109.590 148.890 109.870 149.170 ;
        RECT 110.110 148.890 110.390 149.170 ;
        RECT 109.750 147.130 110.030 147.410 ;
        RECT 110.270 147.130 110.550 147.410 ;
        RECT 103.630 144.930 103.910 145.210 ;
        RECT 104.150 144.930 104.430 145.210 ;
        RECT 107.590 144.930 107.870 145.210 ;
        RECT 108.110 144.930 108.390 145.210 ;
        RECT 109.590 145.370 109.870 145.650 ;
        RECT 110.110 145.370 110.390 145.650 ;
        RECT 103.630 143.170 103.910 143.450 ;
        RECT 104.150 143.170 104.430 143.450 ;
        RECT 107.590 143.170 107.870 143.450 ;
        RECT 108.110 143.170 108.390 143.450 ;
        RECT 103.630 142.290 103.910 142.570 ;
        RECT 104.150 142.290 104.430 142.570 ;
        RECT 107.590 141.410 107.870 141.690 ;
        RECT 108.110 141.410 108.390 141.690 ;
        RECT 107.590 140.530 107.870 140.810 ;
        RECT 108.110 140.530 108.390 140.810 ;
        RECT 109.590 140.090 109.870 140.370 ;
        RECT 110.110 140.090 110.390 140.370 ;
        RECT 103.630 137.890 103.910 138.170 ;
        RECT 104.150 137.890 104.430 138.170 ;
        RECT 107.590 137.890 107.870 138.170 ;
        RECT 108.110 137.890 108.390 138.170 ;
        RECT 103.630 137.010 103.910 137.290 ;
        RECT 104.150 137.010 104.430 137.290 ;
        RECT 109.750 136.570 110.030 136.850 ;
        RECT 110.270 136.570 110.550 136.850 ;
        RECT 103.630 135.250 103.910 135.530 ;
        RECT 104.150 135.250 104.430 135.530 ;
        RECT 107.590 135.250 107.870 135.530 ;
        RECT 108.110 135.250 108.390 135.530 ;
        RECT 90.870 134.370 91.150 134.650 ;
        RECT 91.390 134.370 91.670 134.650 ;
        RECT 94.830 134.370 95.110 134.650 ;
        RECT 95.350 134.370 95.630 134.650 ;
        RECT 116.070 181.890 116.350 182.170 ;
        RECT 116.590 181.890 116.870 182.170 ;
        RECT 120.030 181.890 120.310 182.170 ;
        RECT 120.550 181.890 120.830 182.170 ;
        RECT 113.910 180.740 114.190 181.020 ;
        RECT 114.430 180.740 114.710 181.020 ;
        RECT 116.070 180.130 116.350 180.410 ;
        RECT 116.590 180.130 116.870 180.410 ;
        RECT 120.030 180.130 120.310 180.410 ;
        RECT 120.550 180.130 120.830 180.410 ;
        RECT 116.070 179.250 116.350 179.530 ;
        RECT 116.590 179.250 116.870 179.530 ;
        RECT 113.910 178.810 114.190 179.090 ;
        RECT 114.430 178.810 114.710 179.090 ;
        RECT 116.070 177.490 116.350 177.770 ;
        RECT 116.590 177.490 116.870 177.770 ;
        RECT 120.030 177.490 120.310 177.770 ;
        RECT 120.550 177.490 120.830 177.770 ;
        RECT 116.070 176.610 116.350 176.890 ;
        RECT 116.590 176.610 116.870 176.890 ;
        RECT 120.030 176.610 120.310 176.890 ;
        RECT 120.550 176.610 120.830 176.890 ;
        RECT 122.190 177.930 122.470 178.210 ;
        RECT 122.710 177.930 122.990 178.210 ;
        RECT 116.070 174.850 116.350 175.130 ;
        RECT 116.590 174.850 116.870 175.130 ;
        RECT 120.030 174.850 120.310 175.130 ;
        RECT 120.550 174.850 120.830 175.130 ;
        RECT 113.910 173.530 114.190 173.810 ;
        RECT 114.430 173.530 114.710 173.810 ;
        RECT 116.070 173.090 116.350 173.370 ;
        RECT 116.590 173.090 116.870 173.370 ;
        RECT 120.030 173.090 120.310 173.370 ;
        RECT 120.550 173.090 120.830 173.370 ;
        RECT 114.070 167.370 114.350 167.650 ;
        RECT 114.590 167.370 114.870 167.650 ;
        RECT 120.030 166.930 120.310 167.210 ;
        RECT 120.550 166.930 120.830 167.210 ;
        RECT 113.910 166.490 114.190 166.770 ;
        RECT 114.430 166.490 114.710 166.770 ;
        RECT 116.070 166.050 116.350 166.330 ;
        RECT 116.590 166.050 116.870 166.330 ;
        RECT 120.030 165.170 120.310 165.450 ;
        RECT 120.550 165.170 120.830 165.450 ;
        RECT 114.070 163.850 114.350 164.130 ;
        RECT 114.590 163.850 114.870 164.130 ;
        RECT 120.030 163.410 120.310 163.690 ;
        RECT 120.550 163.410 120.830 163.690 ;
        RECT 120.030 162.530 120.310 162.810 ;
        RECT 120.550 162.530 120.830 162.810 ;
        RECT 120.030 161.650 120.310 161.930 ;
        RECT 120.550 161.650 120.830 161.930 ;
        RECT 120.030 159.890 120.310 160.170 ;
        RECT 120.550 159.890 120.830 160.170 ;
        RECT 116.070 159.010 116.350 159.290 ;
        RECT 116.590 159.010 116.870 159.290 ;
        RECT 116.070 158.130 116.350 158.410 ;
        RECT 116.590 158.130 116.870 158.410 ;
        RECT 120.030 158.130 120.310 158.410 ;
        RECT 120.550 158.130 120.830 158.410 ;
        RECT 116.070 156.370 116.350 156.650 ;
        RECT 116.590 156.370 116.870 156.650 ;
        RECT 120.030 156.370 120.310 156.650 ;
        RECT 120.550 156.370 120.830 156.650 ;
        RECT 120.030 155.490 120.310 155.770 ;
        RECT 120.550 155.490 120.830 155.770 ;
        RECT 122.190 161.210 122.470 161.490 ;
        RECT 122.710 161.210 122.990 161.490 ;
        RECT 116.070 154.610 116.350 154.890 ;
        RECT 116.590 154.610 116.870 154.890 ;
        RECT 120.030 154.610 120.310 154.890 ;
        RECT 120.550 154.610 120.830 154.890 ;
        RECT 116.070 153.730 116.350 154.010 ;
        RECT 116.590 153.730 116.870 154.010 ;
        RECT 120.030 153.730 120.310 154.010 ;
        RECT 120.550 153.730 120.830 154.010 ;
        RECT 116.070 151.970 116.350 152.250 ;
        RECT 116.590 151.970 116.870 152.250 ;
        RECT 116.230 151.260 116.510 151.540 ;
        RECT 116.750 151.260 117.030 151.540 ;
        RECT 120.030 151.970 120.310 152.250 ;
        RECT 120.550 151.970 120.830 152.250 ;
        RECT 116.070 150.210 116.350 150.490 ;
        RECT 116.590 150.210 116.870 150.490 ;
        RECT 120.030 150.210 120.310 150.490 ;
        RECT 120.550 150.210 120.830 150.490 ;
        RECT 120.030 149.330 120.310 149.610 ;
        RECT 120.550 149.330 120.830 149.610 ;
        RECT 122.190 150.650 122.470 150.930 ;
        RECT 122.710 150.650 122.990 150.930 ;
        RECT 122.190 148.010 122.470 148.290 ;
        RECT 122.710 148.010 122.990 148.290 ;
        RECT 120.030 147.570 120.310 147.850 ;
        RECT 120.550 147.570 120.830 147.850 ;
        RECT 114.070 144.490 114.350 144.770 ;
        RECT 114.590 144.490 114.870 144.770 ;
        RECT 120.030 145.810 120.310 146.090 ;
        RECT 120.550 145.810 120.830 146.090 ;
        RECT 122.190 145.370 122.470 145.650 ;
        RECT 122.710 145.370 122.990 145.650 ;
        RECT 120.030 144.050 120.310 144.330 ;
        RECT 120.550 144.050 120.830 144.330 ;
        RECT 116.070 143.170 116.350 143.450 ;
        RECT 116.590 143.170 116.870 143.450 ;
        RECT 114.070 140.970 114.350 141.250 ;
        RECT 114.590 140.970 114.870 141.250 ;
        RECT 120.030 137.010 120.310 137.290 ;
        RECT 120.550 137.010 120.830 137.290 ;
        RECT 113.910 136.570 114.190 136.850 ;
        RECT 114.430 136.570 114.710 136.850 ;
        RECT 116.070 136.130 116.350 136.410 ;
        RECT 116.590 136.130 116.870 136.410 ;
        RECT 116.070 135.250 116.350 135.530 ;
        RECT 116.590 135.250 116.870 135.530 ;
        RECT 120.030 135.250 120.310 135.530 ;
        RECT 120.550 135.250 120.830 135.530 ;
        RECT 103.630 134.370 103.910 134.650 ;
        RECT 104.150 134.370 104.430 134.650 ;
        RECT 107.590 134.370 107.870 134.650 ;
        RECT 108.110 134.370 108.390 134.650 ;
        RECT 116.070 134.370 116.350 134.650 ;
        RECT 116.590 134.370 116.870 134.650 ;
        RECT 120.030 134.370 120.310 134.650 ;
        RECT 120.550 134.370 120.830 134.650 ;
        RECT 22.830 105.510 23.110 105.790 ;
        RECT 22.830 104.990 23.110 105.270 ;
        RECT 56.180 105.250 56.460 105.530 ;
        RECT 56.700 105.250 56.980 105.530 ;
        RECT 79.280 105.250 79.560 105.530 ;
        RECT 79.800 105.250 80.080 105.530 ;
        RECT 113.150 105.510 113.430 105.790 ;
        RECT 113.150 104.990 113.430 105.270 ;
        RECT 21.510 102.490 21.790 102.770 ;
        RECT 25.470 102.490 25.750 102.770 ;
        RECT 42.630 102.490 42.910 102.770 ;
        RECT 46.590 102.490 46.870 102.770 ;
        RECT 21.510 101.970 21.790 102.250 ;
        RECT 25.470 101.970 25.750 102.250 ;
        RECT 42.630 101.970 42.910 102.250 ;
        RECT 46.590 101.970 46.870 102.250 ;
        RECT 56.180 102.230 56.460 102.510 ;
        RECT 56.700 102.230 56.980 102.510 ;
        RECT 79.280 102.230 79.560 102.510 ;
        RECT 79.800 102.230 80.080 102.510 ;
        RECT 89.390 102.490 89.670 102.770 ;
        RECT 93.350 102.490 93.630 102.770 ;
        RECT 110.510 102.490 110.790 102.770 ;
        RECT 114.470 102.490 114.750 102.770 ;
        RECT 89.390 101.970 89.670 102.250 ;
        RECT 93.350 101.970 93.630 102.250 ;
        RECT 110.510 101.970 110.790 102.250 ;
        RECT 114.470 101.970 114.750 102.250 ;
        RECT 18.870 99.470 19.150 99.750 ;
        RECT 20.190 99.470 20.470 99.750 ;
        RECT 26.790 99.470 27.070 99.750 ;
        RECT 28.110 99.470 28.390 99.750 ;
        RECT 39.990 99.470 40.270 99.750 ;
        RECT 41.310 99.470 41.590 99.750 ;
        RECT 47.910 99.470 48.190 99.750 ;
        RECT 49.230 99.470 49.510 99.750 ;
        RECT 18.870 98.950 19.150 99.230 ;
        RECT 20.190 98.950 20.470 99.230 ;
        RECT 26.790 98.950 27.070 99.230 ;
        RECT 28.110 98.950 28.390 99.230 ;
        RECT 39.990 98.950 40.270 99.230 ;
        RECT 41.310 98.950 41.590 99.230 ;
        RECT 47.910 98.950 48.190 99.230 ;
        RECT 49.230 98.950 49.510 99.230 ;
        RECT 56.180 99.210 56.460 99.490 ;
        RECT 56.700 99.210 56.980 99.490 ;
        RECT 79.280 99.210 79.560 99.490 ;
        RECT 79.800 99.210 80.080 99.490 ;
        RECT 86.750 99.470 87.030 99.750 ;
        RECT 88.070 99.470 88.350 99.750 ;
        RECT 94.670 99.470 94.950 99.750 ;
        RECT 95.990 99.470 96.270 99.750 ;
        RECT 107.870 99.470 108.150 99.750 ;
        RECT 109.190 99.470 109.470 99.750 ;
        RECT 115.790 99.470 116.070 99.750 ;
        RECT 117.110 99.470 117.390 99.750 ;
        RECT 86.750 98.950 87.030 99.230 ;
        RECT 88.070 98.950 88.350 99.230 ;
        RECT 94.670 98.950 94.950 99.230 ;
        RECT 95.990 98.950 96.270 99.230 ;
        RECT 107.870 98.950 108.150 99.230 ;
        RECT 109.190 98.950 109.470 99.230 ;
        RECT 115.790 98.950 116.070 99.230 ;
        RECT 117.110 98.950 117.390 99.230 ;
        RECT 24.150 96.450 24.430 96.730 ;
        RECT 43.950 96.450 44.230 96.730 ;
        RECT 24.150 95.930 24.430 96.210 ;
        RECT 43.950 95.930 44.230 96.210 ;
        RECT 56.180 96.190 56.460 96.470 ;
        RECT 56.700 96.190 56.980 96.470 ;
        RECT 79.280 96.190 79.560 96.470 ;
        RECT 79.800 96.190 80.080 96.470 ;
        RECT 92.030 96.450 92.310 96.730 ;
        RECT 111.830 96.450 112.110 96.730 ;
        RECT 92.030 95.930 92.310 96.210 ;
        RECT 111.830 95.930 112.110 96.210 ;
        RECT 13.590 93.430 13.870 93.710 ;
        RECT 14.910 93.430 15.190 93.710 ;
        RECT 16.230 93.430 16.510 93.710 ;
        RECT 17.550 93.430 17.830 93.710 ;
        RECT 29.430 93.430 29.710 93.710 ;
        RECT 30.750 93.430 31.030 93.710 ;
        RECT 32.070 93.430 32.350 93.710 ;
        RECT 33.390 93.430 33.670 93.710 ;
        RECT 34.710 93.430 34.990 93.710 ;
        RECT 36.030 93.430 36.310 93.710 ;
        RECT 37.350 93.430 37.630 93.710 ;
        RECT 38.670 93.430 38.950 93.710 ;
        RECT 50.550 93.430 50.830 93.710 ;
        RECT 51.870 93.430 52.150 93.710 ;
        RECT 53.190 93.430 53.470 93.710 ;
        RECT 54.510 93.430 54.790 93.710 ;
        RECT 13.590 92.910 13.870 93.190 ;
        RECT 14.910 92.910 15.190 93.190 ;
        RECT 16.230 92.910 16.510 93.190 ;
        RECT 17.550 92.910 17.830 93.190 ;
        RECT 29.430 92.910 29.710 93.190 ;
        RECT 30.750 92.910 31.030 93.190 ;
        RECT 32.070 92.910 32.350 93.190 ;
        RECT 33.390 92.910 33.670 93.190 ;
        RECT 34.710 92.910 34.990 93.190 ;
        RECT 36.030 92.910 36.310 93.190 ;
        RECT 37.350 92.910 37.630 93.190 ;
        RECT 38.670 92.910 38.950 93.190 ;
        RECT 50.550 92.910 50.830 93.190 ;
        RECT 51.870 92.910 52.150 93.190 ;
        RECT 53.190 92.910 53.470 93.190 ;
        RECT 54.510 92.910 54.790 93.190 ;
        RECT 56.180 93.170 56.460 93.450 ;
        RECT 56.700 93.170 56.980 93.450 ;
        RECT 79.280 93.170 79.560 93.450 ;
        RECT 79.800 93.170 80.080 93.450 ;
        RECT 81.470 93.430 81.750 93.710 ;
        RECT 82.790 93.430 83.070 93.710 ;
        RECT 84.110 93.430 84.390 93.710 ;
        RECT 85.430 93.430 85.710 93.710 ;
        RECT 97.310 93.430 97.590 93.710 ;
        RECT 98.630 93.430 98.910 93.710 ;
        RECT 99.950 93.430 100.230 93.710 ;
        RECT 101.270 93.430 101.550 93.710 ;
        RECT 102.590 93.430 102.870 93.710 ;
        RECT 103.910 93.430 104.190 93.710 ;
        RECT 105.230 93.430 105.510 93.710 ;
        RECT 106.550 93.430 106.830 93.710 ;
        RECT 118.430 93.430 118.710 93.710 ;
        RECT 119.750 93.430 120.030 93.710 ;
        RECT 121.070 93.430 121.350 93.710 ;
        RECT 122.390 93.430 122.670 93.710 ;
        RECT 81.470 92.910 81.750 93.190 ;
        RECT 82.790 92.910 83.070 93.190 ;
        RECT 84.110 92.910 84.390 93.190 ;
        RECT 85.430 92.910 85.710 93.190 ;
        RECT 97.310 92.910 97.590 93.190 ;
        RECT 98.630 92.910 98.910 93.190 ;
        RECT 99.950 92.910 100.230 93.190 ;
        RECT 101.270 92.910 101.550 93.190 ;
        RECT 102.590 92.910 102.870 93.190 ;
        RECT 103.910 92.910 104.190 93.190 ;
        RECT 105.230 92.910 105.510 93.190 ;
        RECT 106.550 92.910 106.830 93.190 ;
        RECT 118.430 92.910 118.710 93.190 ;
        RECT 119.750 92.910 120.030 93.190 ;
        RECT 121.070 92.910 121.350 93.190 ;
        RECT 122.390 92.910 122.670 93.190 ;
        RECT 7.350 90.090 7.630 90.370 ;
        RECT 7.870 90.090 8.150 90.370 ;
        RECT 45.270 90.410 45.550 90.690 ;
        RECT 7.350 89.570 7.630 89.850 ;
        RECT 7.870 89.570 8.150 89.850 ;
        RECT 45.270 89.890 45.550 90.170 ;
        RECT 56.180 90.150 56.460 90.430 ;
        RECT 56.700 90.150 56.980 90.430 ;
        RECT 79.280 90.150 79.560 90.430 ;
        RECT 79.800 90.150 80.080 90.430 ;
        RECT 90.710 90.410 90.990 90.690 ;
        RECT 90.710 89.890 90.990 90.170 ;
        RECT 128.660 89.750 128.940 90.030 ;
        RECT 128.660 89.230 128.940 89.510 ;
        RECT 22.830 88.510 23.110 88.790 ;
        RECT 22.830 87.990 23.110 88.270 ;
        RECT 56.180 88.250 56.460 88.530 ;
        RECT 56.700 88.250 56.980 88.530 ;
        RECT 79.280 88.250 79.560 88.530 ;
        RECT 79.800 88.250 80.080 88.530 ;
        RECT 113.150 88.510 113.430 88.790 ;
        RECT 113.150 87.990 113.430 88.270 ;
        RECT 21.510 85.490 21.790 85.770 ;
        RECT 25.470 85.490 25.750 85.770 ;
        RECT 42.630 85.490 42.910 85.770 ;
        RECT 46.590 85.490 46.870 85.770 ;
        RECT 21.510 84.970 21.790 85.250 ;
        RECT 25.470 84.970 25.750 85.250 ;
        RECT 42.630 84.970 42.910 85.250 ;
        RECT 46.590 84.970 46.870 85.250 ;
        RECT 56.180 85.230 56.460 85.510 ;
        RECT 56.700 85.230 56.980 85.510 ;
        RECT 79.280 85.230 79.560 85.510 ;
        RECT 79.800 85.230 80.080 85.510 ;
        RECT 89.390 85.490 89.670 85.770 ;
        RECT 93.350 85.490 93.630 85.770 ;
        RECT 110.510 85.490 110.790 85.770 ;
        RECT 114.470 85.490 114.750 85.770 ;
        RECT 89.390 84.970 89.670 85.250 ;
        RECT 93.350 84.970 93.630 85.250 ;
        RECT 110.510 84.970 110.790 85.250 ;
        RECT 114.470 84.970 114.750 85.250 ;
        RECT 18.870 82.470 19.150 82.750 ;
        RECT 20.190 82.470 20.470 82.750 ;
        RECT 26.790 82.470 27.070 82.750 ;
        RECT 28.110 82.470 28.390 82.750 ;
        RECT 39.990 82.470 40.270 82.750 ;
        RECT 41.310 82.470 41.590 82.750 ;
        RECT 47.910 82.470 48.190 82.750 ;
        RECT 49.230 82.470 49.510 82.750 ;
        RECT 18.870 81.950 19.150 82.230 ;
        RECT 20.190 81.950 20.470 82.230 ;
        RECT 26.790 81.950 27.070 82.230 ;
        RECT 28.110 81.950 28.390 82.230 ;
        RECT 39.990 81.950 40.270 82.230 ;
        RECT 41.310 81.950 41.590 82.230 ;
        RECT 47.910 81.950 48.190 82.230 ;
        RECT 49.230 81.950 49.510 82.230 ;
        RECT 56.180 82.210 56.460 82.490 ;
        RECT 56.700 82.210 56.980 82.490 ;
        RECT 79.280 82.210 79.560 82.490 ;
        RECT 79.800 82.210 80.080 82.490 ;
        RECT 86.750 82.470 87.030 82.750 ;
        RECT 88.070 82.470 88.350 82.750 ;
        RECT 94.670 82.470 94.950 82.750 ;
        RECT 95.990 82.470 96.270 82.750 ;
        RECT 107.870 82.470 108.150 82.750 ;
        RECT 109.190 82.470 109.470 82.750 ;
        RECT 115.790 82.470 116.070 82.750 ;
        RECT 117.110 82.470 117.390 82.750 ;
        RECT 86.750 81.950 87.030 82.230 ;
        RECT 88.070 81.950 88.350 82.230 ;
        RECT 94.670 81.950 94.950 82.230 ;
        RECT 95.990 81.950 96.270 82.230 ;
        RECT 107.870 81.950 108.150 82.230 ;
        RECT 109.190 81.950 109.470 82.230 ;
        RECT 115.790 81.950 116.070 82.230 ;
        RECT 117.110 81.950 117.390 82.230 ;
        RECT 24.150 79.450 24.430 79.730 ;
        RECT 43.950 79.450 44.230 79.730 ;
        RECT 24.150 78.930 24.430 79.210 ;
        RECT 43.950 78.930 44.230 79.210 ;
        RECT 56.180 79.190 56.460 79.470 ;
        RECT 56.700 79.190 56.980 79.470 ;
        RECT 79.280 79.190 79.560 79.470 ;
        RECT 79.800 79.190 80.080 79.470 ;
        RECT 92.030 79.450 92.310 79.730 ;
        RECT 111.830 79.450 112.110 79.730 ;
        RECT 92.030 78.930 92.310 79.210 ;
        RECT 111.830 78.930 112.110 79.210 ;
        RECT 13.590 76.430 13.870 76.710 ;
        RECT 14.910 76.430 15.190 76.710 ;
        RECT 16.230 76.430 16.510 76.710 ;
        RECT 17.550 76.430 17.830 76.710 ;
        RECT 29.430 76.430 29.710 76.710 ;
        RECT 30.750 76.430 31.030 76.710 ;
        RECT 32.070 76.430 32.350 76.710 ;
        RECT 33.390 76.430 33.670 76.710 ;
        RECT 34.710 76.430 34.990 76.710 ;
        RECT 36.030 76.430 36.310 76.710 ;
        RECT 37.350 76.430 37.630 76.710 ;
        RECT 38.670 76.430 38.950 76.710 ;
        RECT 50.550 76.430 50.830 76.710 ;
        RECT 51.870 76.430 52.150 76.710 ;
        RECT 53.190 76.430 53.470 76.710 ;
        RECT 54.510 76.430 54.790 76.710 ;
        RECT 13.590 75.910 13.870 76.190 ;
        RECT 14.910 75.910 15.190 76.190 ;
        RECT 16.230 75.910 16.510 76.190 ;
        RECT 17.550 75.910 17.830 76.190 ;
        RECT 29.430 75.910 29.710 76.190 ;
        RECT 30.750 75.910 31.030 76.190 ;
        RECT 32.070 75.910 32.350 76.190 ;
        RECT 33.390 75.910 33.670 76.190 ;
        RECT 34.710 75.910 34.990 76.190 ;
        RECT 36.030 75.910 36.310 76.190 ;
        RECT 37.350 75.910 37.630 76.190 ;
        RECT 38.670 75.910 38.950 76.190 ;
        RECT 50.550 75.910 50.830 76.190 ;
        RECT 51.870 75.910 52.150 76.190 ;
        RECT 53.190 75.910 53.470 76.190 ;
        RECT 54.510 75.910 54.790 76.190 ;
        RECT 56.180 76.170 56.460 76.450 ;
        RECT 56.700 76.170 56.980 76.450 ;
        RECT 79.280 76.170 79.560 76.450 ;
        RECT 79.800 76.170 80.080 76.450 ;
        RECT 81.470 76.430 81.750 76.710 ;
        RECT 82.790 76.430 83.070 76.710 ;
        RECT 84.110 76.430 84.390 76.710 ;
        RECT 85.430 76.430 85.710 76.710 ;
        RECT 97.310 76.430 97.590 76.710 ;
        RECT 98.630 76.430 98.910 76.710 ;
        RECT 99.950 76.430 100.230 76.710 ;
        RECT 101.270 76.430 101.550 76.710 ;
        RECT 102.590 76.430 102.870 76.710 ;
        RECT 103.910 76.430 104.190 76.710 ;
        RECT 105.230 76.430 105.510 76.710 ;
        RECT 106.550 76.430 106.830 76.710 ;
        RECT 118.430 76.430 118.710 76.710 ;
        RECT 119.750 76.430 120.030 76.710 ;
        RECT 121.070 76.430 121.350 76.710 ;
        RECT 122.390 76.430 122.670 76.710 ;
        RECT 81.470 75.910 81.750 76.190 ;
        RECT 82.790 75.910 83.070 76.190 ;
        RECT 84.110 75.910 84.390 76.190 ;
        RECT 85.430 75.910 85.710 76.190 ;
        RECT 97.310 75.910 97.590 76.190 ;
        RECT 98.630 75.910 98.910 76.190 ;
        RECT 99.950 75.910 100.230 76.190 ;
        RECT 101.270 75.910 101.550 76.190 ;
        RECT 102.590 75.910 102.870 76.190 ;
        RECT 103.910 75.910 104.190 76.190 ;
        RECT 105.230 75.910 105.510 76.190 ;
        RECT 106.550 75.910 106.830 76.190 ;
        RECT 118.430 75.910 118.710 76.190 ;
        RECT 119.750 75.910 120.030 76.190 ;
        RECT 121.070 75.910 121.350 76.190 ;
        RECT 122.390 75.910 122.670 76.190 ;
        RECT 7.350 73.090 7.630 73.370 ;
        RECT 7.870 73.090 8.150 73.370 ;
        RECT 45.270 73.410 45.550 73.690 ;
        RECT 7.350 72.570 7.630 72.850 ;
        RECT 7.870 72.570 8.150 72.850 ;
        RECT 45.270 72.890 45.550 73.170 ;
        RECT 56.180 73.150 56.460 73.430 ;
        RECT 56.700 73.150 56.980 73.430 ;
        RECT 79.280 73.150 79.560 73.430 ;
        RECT 79.800 73.150 80.080 73.430 ;
        RECT 90.710 73.410 90.990 73.690 ;
        RECT 90.710 72.890 90.990 73.170 ;
        RECT 128.660 72.750 128.940 73.030 ;
        RECT 128.660 72.230 128.940 72.510 ;
        RECT 22.830 71.510 23.110 71.790 ;
        RECT 22.830 70.990 23.110 71.270 ;
        RECT 56.180 71.250 56.460 71.530 ;
        RECT 56.700 71.250 56.980 71.530 ;
        RECT 79.280 71.250 79.560 71.530 ;
        RECT 79.800 71.250 80.080 71.530 ;
        RECT 113.150 71.510 113.430 71.790 ;
        RECT 113.150 70.990 113.430 71.270 ;
        RECT 21.510 68.490 21.790 68.770 ;
        RECT 25.470 68.490 25.750 68.770 ;
        RECT 42.630 68.490 42.910 68.770 ;
        RECT 46.590 68.490 46.870 68.770 ;
        RECT 21.510 67.970 21.790 68.250 ;
        RECT 25.470 67.970 25.750 68.250 ;
        RECT 42.630 67.970 42.910 68.250 ;
        RECT 46.590 67.970 46.870 68.250 ;
        RECT 56.180 68.230 56.460 68.510 ;
        RECT 56.700 68.230 56.980 68.510 ;
        RECT 79.280 68.230 79.560 68.510 ;
        RECT 79.800 68.230 80.080 68.510 ;
        RECT 89.390 68.490 89.670 68.770 ;
        RECT 93.350 68.490 93.630 68.770 ;
        RECT 110.510 68.490 110.790 68.770 ;
        RECT 114.470 68.490 114.750 68.770 ;
        RECT 89.390 67.970 89.670 68.250 ;
        RECT 93.350 67.970 93.630 68.250 ;
        RECT 110.510 67.970 110.790 68.250 ;
        RECT 114.470 67.970 114.750 68.250 ;
        RECT 18.870 65.470 19.150 65.750 ;
        RECT 20.190 65.470 20.470 65.750 ;
        RECT 26.790 65.470 27.070 65.750 ;
        RECT 28.110 65.470 28.390 65.750 ;
        RECT 39.990 65.470 40.270 65.750 ;
        RECT 41.310 65.470 41.590 65.750 ;
        RECT 47.910 65.470 48.190 65.750 ;
        RECT 49.230 65.470 49.510 65.750 ;
        RECT 18.870 64.950 19.150 65.230 ;
        RECT 20.190 64.950 20.470 65.230 ;
        RECT 26.790 64.950 27.070 65.230 ;
        RECT 28.110 64.950 28.390 65.230 ;
        RECT 39.990 64.950 40.270 65.230 ;
        RECT 41.310 64.950 41.590 65.230 ;
        RECT 47.910 64.950 48.190 65.230 ;
        RECT 49.230 64.950 49.510 65.230 ;
        RECT 56.180 65.210 56.460 65.490 ;
        RECT 56.700 65.210 56.980 65.490 ;
        RECT 79.280 65.210 79.560 65.490 ;
        RECT 79.800 65.210 80.080 65.490 ;
        RECT 86.750 65.470 87.030 65.750 ;
        RECT 88.070 65.470 88.350 65.750 ;
        RECT 94.670 65.470 94.950 65.750 ;
        RECT 95.990 65.470 96.270 65.750 ;
        RECT 107.870 65.470 108.150 65.750 ;
        RECT 109.190 65.470 109.470 65.750 ;
        RECT 115.790 65.470 116.070 65.750 ;
        RECT 117.110 65.470 117.390 65.750 ;
        RECT 86.750 64.950 87.030 65.230 ;
        RECT 88.070 64.950 88.350 65.230 ;
        RECT 94.670 64.950 94.950 65.230 ;
        RECT 95.990 64.950 96.270 65.230 ;
        RECT 107.870 64.950 108.150 65.230 ;
        RECT 109.190 64.950 109.470 65.230 ;
        RECT 115.790 64.950 116.070 65.230 ;
        RECT 117.110 64.950 117.390 65.230 ;
        RECT 24.150 62.450 24.430 62.730 ;
        RECT 43.950 62.450 44.230 62.730 ;
        RECT 24.150 61.930 24.430 62.210 ;
        RECT 43.950 61.930 44.230 62.210 ;
        RECT 56.180 62.190 56.460 62.470 ;
        RECT 56.700 62.190 56.980 62.470 ;
        RECT 79.280 62.190 79.560 62.470 ;
        RECT 79.800 62.190 80.080 62.470 ;
        RECT 92.030 62.450 92.310 62.730 ;
        RECT 111.830 62.450 112.110 62.730 ;
        RECT 92.030 61.930 92.310 62.210 ;
        RECT 111.830 61.930 112.110 62.210 ;
        RECT 13.590 59.430 13.870 59.710 ;
        RECT 14.910 59.430 15.190 59.710 ;
        RECT 16.230 59.430 16.510 59.710 ;
        RECT 17.550 59.430 17.830 59.710 ;
        RECT 29.430 59.430 29.710 59.710 ;
        RECT 30.750 59.430 31.030 59.710 ;
        RECT 32.070 59.430 32.350 59.710 ;
        RECT 33.390 59.430 33.670 59.710 ;
        RECT 34.710 59.430 34.990 59.710 ;
        RECT 36.030 59.430 36.310 59.710 ;
        RECT 37.350 59.430 37.630 59.710 ;
        RECT 38.670 59.430 38.950 59.710 ;
        RECT 50.550 59.430 50.830 59.710 ;
        RECT 51.870 59.430 52.150 59.710 ;
        RECT 53.190 59.430 53.470 59.710 ;
        RECT 54.510 59.430 54.790 59.710 ;
        RECT 13.590 58.910 13.870 59.190 ;
        RECT 14.910 58.910 15.190 59.190 ;
        RECT 16.230 58.910 16.510 59.190 ;
        RECT 17.550 58.910 17.830 59.190 ;
        RECT 29.430 58.910 29.710 59.190 ;
        RECT 30.750 58.910 31.030 59.190 ;
        RECT 32.070 58.910 32.350 59.190 ;
        RECT 33.390 58.910 33.670 59.190 ;
        RECT 34.710 58.910 34.990 59.190 ;
        RECT 36.030 58.910 36.310 59.190 ;
        RECT 37.350 58.910 37.630 59.190 ;
        RECT 38.670 58.910 38.950 59.190 ;
        RECT 50.550 58.910 50.830 59.190 ;
        RECT 51.870 58.910 52.150 59.190 ;
        RECT 53.190 58.910 53.470 59.190 ;
        RECT 54.510 58.910 54.790 59.190 ;
        RECT 56.180 59.170 56.460 59.450 ;
        RECT 56.700 59.170 56.980 59.450 ;
        RECT 79.280 59.170 79.560 59.450 ;
        RECT 79.800 59.170 80.080 59.450 ;
        RECT 81.470 59.430 81.750 59.710 ;
        RECT 82.790 59.430 83.070 59.710 ;
        RECT 84.110 59.430 84.390 59.710 ;
        RECT 85.430 59.430 85.710 59.710 ;
        RECT 97.310 59.430 97.590 59.710 ;
        RECT 98.630 59.430 98.910 59.710 ;
        RECT 99.950 59.430 100.230 59.710 ;
        RECT 101.270 59.430 101.550 59.710 ;
        RECT 102.590 59.430 102.870 59.710 ;
        RECT 103.910 59.430 104.190 59.710 ;
        RECT 105.230 59.430 105.510 59.710 ;
        RECT 106.550 59.430 106.830 59.710 ;
        RECT 118.430 59.430 118.710 59.710 ;
        RECT 119.750 59.430 120.030 59.710 ;
        RECT 121.070 59.430 121.350 59.710 ;
        RECT 122.390 59.430 122.670 59.710 ;
        RECT 81.470 58.910 81.750 59.190 ;
        RECT 82.790 58.910 83.070 59.190 ;
        RECT 84.110 58.910 84.390 59.190 ;
        RECT 85.430 58.910 85.710 59.190 ;
        RECT 97.310 58.910 97.590 59.190 ;
        RECT 98.630 58.910 98.910 59.190 ;
        RECT 99.950 58.910 100.230 59.190 ;
        RECT 101.270 58.910 101.550 59.190 ;
        RECT 102.590 58.910 102.870 59.190 ;
        RECT 103.910 58.910 104.190 59.190 ;
        RECT 105.230 58.910 105.510 59.190 ;
        RECT 106.550 58.910 106.830 59.190 ;
        RECT 118.430 58.910 118.710 59.190 ;
        RECT 119.750 58.910 120.030 59.190 ;
        RECT 121.070 58.910 121.350 59.190 ;
        RECT 122.390 58.910 122.670 59.190 ;
        RECT 7.350 56.090 7.630 56.370 ;
        RECT 7.870 56.090 8.150 56.370 ;
        RECT 45.270 56.410 45.550 56.690 ;
        RECT 7.350 55.570 7.630 55.850 ;
        RECT 7.870 55.570 8.150 55.850 ;
        RECT 45.270 55.890 45.550 56.170 ;
        RECT 56.730 56.410 57.010 56.690 ;
        RECT 56.730 55.890 57.010 56.170 ;
        RECT 79.250 56.410 79.530 56.690 ;
        RECT 79.250 55.890 79.530 56.170 ;
        RECT 90.710 56.410 90.990 56.690 ;
        RECT 90.710 55.890 90.990 56.170 ;
        RECT 128.660 55.750 128.940 56.030 ;
        RECT 128.660 55.230 128.940 55.510 ;
        RECT 22.830 54.510 23.110 54.790 ;
        RECT 22.830 53.990 23.110 54.270 ;
        RECT 56.180 54.250 56.460 54.530 ;
        RECT 56.700 54.250 56.980 54.530 ;
        RECT 79.280 54.250 79.560 54.530 ;
        RECT 79.800 54.250 80.080 54.530 ;
        RECT 113.150 54.510 113.430 54.790 ;
        RECT 113.150 53.990 113.430 54.270 ;
        RECT 21.510 51.490 21.790 51.770 ;
        RECT 25.470 51.490 25.750 51.770 ;
        RECT 42.630 51.490 42.910 51.770 ;
        RECT 46.590 51.490 46.870 51.770 ;
        RECT 21.510 50.970 21.790 51.250 ;
        RECT 25.470 50.970 25.750 51.250 ;
        RECT 42.630 50.970 42.910 51.250 ;
        RECT 46.590 50.970 46.870 51.250 ;
        RECT 56.180 51.230 56.460 51.510 ;
        RECT 56.700 51.230 56.980 51.510 ;
        RECT 79.280 51.230 79.560 51.510 ;
        RECT 79.800 51.230 80.080 51.510 ;
        RECT 89.390 51.490 89.670 51.770 ;
        RECT 93.350 51.490 93.630 51.770 ;
        RECT 110.510 51.490 110.790 51.770 ;
        RECT 114.470 51.490 114.750 51.770 ;
        RECT 89.390 50.970 89.670 51.250 ;
        RECT 93.350 50.970 93.630 51.250 ;
        RECT 110.510 50.970 110.790 51.250 ;
        RECT 114.470 50.970 114.750 51.250 ;
        RECT 18.870 48.470 19.150 48.750 ;
        RECT 20.190 48.470 20.470 48.750 ;
        RECT 26.790 48.470 27.070 48.750 ;
        RECT 28.110 48.470 28.390 48.750 ;
        RECT 39.990 48.470 40.270 48.750 ;
        RECT 41.310 48.470 41.590 48.750 ;
        RECT 47.910 48.470 48.190 48.750 ;
        RECT 49.230 48.470 49.510 48.750 ;
        RECT 18.870 47.950 19.150 48.230 ;
        RECT 20.190 47.950 20.470 48.230 ;
        RECT 26.790 47.950 27.070 48.230 ;
        RECT 28.110 47.950 28.390 48.230 ;
        RECT 39.990 47.950 40.270 48.230 ;
        RECT 41.310 47.950 41.590 48.230 ;
        RECT 47.910 47.950 48.190 48.230 ;
        RECT 49.230 47.950 49.510 48.230 ;
        RECT 56.180 48.210 56.460 48.490 ;
        RECT 56.700 48.210 56.980 48.490 ;
        RECT 79.280 48.210 79.560 48.490 ;
        RECT 79.800 48.210 80.080 48.490 ;
        RECT 86.750 48.470 87.030 48.750 ;
        RECT 88.070 48.470 88.350 48.750 ;
        RECT 94.670 48.470 94.950 48.750 ;
        RECT 95.990 48.470 96.270 48.750 ;
        RECT 107.870 48.470 108.150 48.750 ;
        RECT 109.190 48.470 109.470 48.750 ;
        RECT 115.790 48.470 116.070 48.750 ;
        RECT 117.110 48.470 117.390 48.750 ;
        RECT 86.750 47.950 87.030 48.230 ;
        RECT 88.070 47.950 88.350 48.230 ;
        RECT 94.670 47.950 94.950 48.230 ;
        RECT 95.990 47.950 96.270 48.230 ;
        RECT 107.870 47.950 108.150 48.230 ;
        RECT 109.190 47.950 109.470 48.230 ;
        RECT 115.790 47.950 116.070 48.230 ;
        RECT 117.110 47.950 117.390 48.230 ;
        RECT 24.150 45.450 24.430 45.730 ;
        RECT 43.950 45.450 44.230 45.730 ;
        RECT 24.150 44.930 24.430 45.210 ;
        RECT 43.950 44.930 44.230 45.210 ;
        RECT 56.180 45.190 56.460 45.470 ;
        RECT 56.700 45.190 56.980 45.470 ;
        RECT 79.280 45.190 79.560 45.470 ;
        RECT 79.800 45.190 80.080 45.470 ;
        RECT 92.030 45.450 92.310 45.730 ;
        RECT 111.830 45.450 112.110 45.730 ;
        RECT 92.030 44.930 92.310 45.210 ;
        RECT 111.830 44.930 112.110 45.210 ;
        RECT 13.590 42.430 13.870 42.710 ;
        RECT 14.910 42.430 15.190 42.710 ;
        RECT 16.230 42.430 16.510 42.710 ;
        RECT 17.550 42.430 17.830 42.710 ;
        RECT 29.430 42.430 29.710 42.710 ;
        RECT 30.750 42.430 31.030 42.710 ;
        RECT 32.070 42.430 32.350 42.710 ;
        RECT 33.390 42.430 33.670 42.710 ;
        RECT 34.710 42.430 34.990 42.710 ;
        RECT 36.030 42.430 36.310 42.710 ;
        RECT 37.350 42.430 37.630 42.710 ;
        RECT 38.670 42.430 38.950 42.710 ;
        RECT 50.550 42.430 50.830 42.710 ;
        RECT 51.870 42.430 52.150 42.710 ;
        RECT 53.190 42.430 53.470 42.710 ;
        RECT 54.510 42.430 54.790 42.710 ;
        RECT 13.590 41.910 13.870 42.190 ;
        RECT 14.910 41.910 15.190 42.190 ;
        RECT 16.230 41.910 16.510 42.190 ;
        RECT 17.550 41.910 17.830 42.190 ;
        RECT 29.430 41.910 29.710 42.190 ;
        RECT 30.750 41.910 31.030 42.190 ;
        RECT 32.070 41.910 32.350 42.190 ;
        RECT 33.390 41.910 33.670 42.190 ;
        RECT 34.710 41.910 34.990 42.190 ;
        RECT 36.030 41.910 36.310 42.190 ;
        RECT 37.350 41.910 37.630 42.190 ;
        RECT 38.670 41.910 38.950 42.190 ;
        RECT 50.550 41.910 50.830 42.190 ;
        RECT 51.870 41.910 52.150 42.190 ;
        RECT 53.190 41.910 53.470 42.190 ;
        RECT 54.510 41.910 54.790 42.190 ;
        RECT 56.180 42.170 56.460 42.450 ;
        RECT 56.700 42.170 56.980 42.450 ;
        RECT 79.280 42.170 79.560 42.450 ;
        RECT 79.800 42.170 80.080 42.450 ;
        RECT 81.470 42.430 81.750 42.710 ;
        RECT 82.790 42.430 83.070 42.710 ;
        RECT 84.110 42.430 84.390 42.710 ;
        RECT 85.430 42.430 85.710 42.710 ;
        RECT 97.310 42.430 97.590 42.710 ;
        RECT 98.630 42.430 98.910 42.710 ;
        RECT 99.950 42.430 100.230 42.710 ;
        RECT 101.270 42.430 101.550 42.710 ;
        RECT 102.590 42.430 102.870 42.710 ;
        RECT 103.910 42.430 104.190 42.710 ;
        RECT 105.230 42.430 105.510 42.710 ;
        RECT 106.550 42.430 106.830 42.710 ;
        RECT 118.430 42.430 118.710 42.710 ;
        RECT 119.750 42.430 120.030 42.710 ;
        RECT 121.070 42.430 121.350 42.710 ;
        RECT 122.390 42.430 122.670 42.710 ;
        RECT 81.470 41.910 81.750 42.190 ;
        RECT 82.790 41.910 83.070 42.190 ;
        RECT 84.110 41.910 84.390 42.190 ;
        RECT 85.430 41.910 85.710 42.190 ;
        RECT 97.310 41.910 97.590 42.190 ;
        RECT 98.630 41.910 98.910 42.190 ;
        RECT 99.950 41.910 100.230 42.190 ;
        RECT 101.270 41.910 101.550 42.190 ;
        RECT 102.590 41.910 102.870 42.190 ;
        RECT 103.910 41.910 104.190 42.190 ;
        RECT 105.230 41.910 105.510 42.190 ;
        RECT 106.550 41.910 106.830 42.190 ;
        RECT 118.430 41.910 118.710 42.190 ;
        RECT 119.750 41.910 120.030 42.190 ;
        RECT 121.070 41.910 121.350 42.190 ;
        RECT 122.390 41.910 122.670 42.190 ;
        RECT 7.350 39.090 7.630 39.370 ;
        RECT 7.870 39.090 8.150 39.370 ;
        RECT 45.270 39.410 45.550 39.690 ;
        RECT 7.350 38.570 7.630 38.850 ;
        RECT 7.870 38.570 8.150 38.850 ;
        RECT 45.270 38.890 45.550 39.170 ;
        RECT 56.180 39.150 56.460 39.430 ;
        RECT 56.700 39.150 56.980 39.430 ;
        RECT 79.280 39.150 79.560 39.430 ;
        RECT 79.800 39.150 80.080 39.430 ;
        RECT 90.710 39.410 90.990 39.690 ;
        RECT 90.710 38.890 90.990 39.170 ;
        RECT 128.660 38.750 128.940 39.030 ;
        RECT 128.660 38.230 128.940 38.510 ;
        RECT 44.550 36.280 45.630 36.600 ;
        RECT 11.790 35.480 12.870 35.800 ;
        RECT 44.550 34.680 45.630 35.000 ;
        RECT 11.790 33.880 12.870 34.200 ;
        RECT 44.550 33.080 45.630 33.400 ;
        RECT 90.630 36.280 91.710 36.600 ;
        RECT 123.390 35.480 124.470 35.800 ;
        RECT 90.630 34.680 91.710 35.000 ;
        RECT 123.390 33.880 124.470 34.200 ;
        RECT 90.630 33.080 91.710 33.400 ;
        RECT 11.790 32.280 12.870 32.600 ;
        RECT 123.390 32.280 124.470 32.600 ;
        RECT 44.550 31.480 45.630 31.800 ;
        RECT 11.790 30.680 12.870 31.000 ;
        RECT 44.550 29.880 45.630 30.200 ;
        RECT 90.630 31.480 91.710 31.800 ;
        RECT 123.390 30.680 124.470 31.000 ;
        RECT 11.790 29.080 12.870 29.400 ;
        RECT 44.550 28.280 45.630 28.600 ;
        RECT 52.330 29.380 52.610 29.660 ;
        RECT 52.850 29.380 53.130 29.660 ;
        RECT 56.290 29.380 56.570 29.660 ;
        RECT 56.810 29.380 57.090 29.660 ;
        RECT 11.790 27.480 12.870 27.800 ;
        RECT 44.550 26.680 45.630 27.000 ;
        RECT 11.790 25.880 12.870 26.200 ;
        RECT 44.550 25.080 45.630 25.400 ;
        RECT 11.790 24.280 12.870 24.600 ;
        RECT 44.550 23.480 45.630 23.800 ;
        RECT 79.170 29.380 79.450 29.660 ;
        RECT 79.690 29.380 79.970 29.660 ;
        RECT 83.130 29.380 83.410 29.660 ;
        RECT 83.650 29.380 83.930 29.660 ;
        RECT 52.330 28.500 52.610 28.780 ;
        RECT 52.850 28.500 53.130 28.780 ;
        RECT 56.290 28.500 56.570 28.780 ;
        RECT 56.810 28.500 57.090 28.780 ;
        RECT 56.290 27.620 56.570 27.900 ;
        RECT 56.810 27.620 57.090 27.900 ;
        RECT 52.330 26.740 52.610 27.020 ;
        RECT 52.850 26.740 53.130 27.020 ;
        RECT 56.290 26.740 56.570 27.020 ;
        RECT 56.810 26.740 57.090 27.020 ;
        RECT 52.330 25.860 52.610 26.140 ;
        RECT 52.850 25.860 53.130 26.140 ;
        RECT 56.290 25.860 56.570 26.140 ;
        RECT 56.810 25.860 57.090 26.140 ;
        RECT 11.790 22.680 12.870 23.000 ;
        RECT 44.550 21.880 45.630 22.200 ;
        RECT 11.790 21.080 12.870 21.400 ;
        RECT 44.550 20.280 45.630 20.600 ;
        RECT 11.790 19.480 12.870 19.800 ;
        RECT 44.550 18.680 45.630 19.000 ;
        RECT 11.790 17.880 12.870 18.200 ;
        RECT 44.550 17.080 45.630 17.400 ;
        RECT 11.790 16.280 12.870 16.600 ;
        RECT 44.550 15.480 45.630 15.800 ;
        RECT 11.790 14.680 12.870 15.000 ;
        RECT 44.550 13.880 45.630 14.200 ;
        RECT 52.330 24.980 52.610 25.260 ;
        RECT 52.850 24.980 53.130 25.260 ;
        RECT 56.290 24.980 56.570 25.260 ;
        RECT 56.810 24.980 57.090 25.260 ;
        RECT 52.330 24.270 52.610 24.550 ;
        RECT 52.850 24.270 53.130 24.550 ;
        RECT 52.330 23.220 52.610 23.500 ;
        RECT 52.850 23.220 53.130 23.500 ;
        RECT 56.290 23.220 56.570 23.500 ;
        RECT 56.810 23.220 57.090 23.500 ;
        RECT 52.330 22.340 52.610 22.620 ;
        RECT 52.850 22.340 53.130 22.620 ;
        RECT 56.130 22.340 56.410 22.620 ;
        RECT 56.650 22.340 56.930 22.620 ;
        RECT 52.330 21.460 52.610 21.740 ;
        RECT 52.850 21.460 53.130 21.740 ;
        RECT 58.450 21.900 58.730 22.180 ;
        RECT 58.970 21.900 59.250 22.180 ;
        RECT 58.450 21.020 58.730 21.300 ;
        RECT 58.970 21.020 59.250 21.300 ;
        RECT 56.290 20.580 56.570 20.860 ;
        RECT 56.810 20.580 57.090 20.860 ;
        RECT 56.290 19.700 56.570 19.980 ;
        RECT 56.810 19.700 57.090 19.980 ;
        RECT 52.330 18.820 52.610 19.100 ;
        RECT 52.850 18.820 53.130 19.100 ;
        RECT 50.170 18.380 50.450 18.660 ;
        RECT 50.690 18.380 50.970 18.660 ;
        RECT 52.330 17.940 52.610 18.220 ;
        RECT 52.850 17.940 53.130 18.220 ;
        RECT 56.290 17.940 56.570 18.220 ;
        RECT 56.810 17.940 57.090 18.220 ;
        RECT 50.170 17.500 50.450 17.780 ;
        RECT 50.690 17.500 50.970 17.780 ;
        RECT 52.330 16.180 52.610 16.460 ;
        RECT 52.850 16.180 53.130 16.460 ;
        RECT 56.290 16.350 56.570 16.630 ;
        RECT 56.810 16.350 57.090 16.630 ;
        RECT 58.370 15.740 58.650 16.020 ;
        RECT 58.890 15.740 59.170 16.020 ;
        RECT 52.330 15.300 52.610 15.580 ;
        RECT 52.850 15.300 53.130 15.580 ;
        RECT 56.290 15.300 56.570 15.580 ;
        RECT 56.810 15.300 57.090 15.580 ;
        RECT 52.330 14.420 52.610 14.700 ;
        RECT 52.850 14.420 53.130 14.700 ;
        RECT 56.290 14.420 56.570 14.700 ;
        RECT 56.810 14.420 57.090 14.700 ;
        RECT 11.790 13.080 12.870 13.400 ;
        RECT 63.330 25.860 63.610 26.140 ;
        RECT 63.850 25.860 64.130 26.140 ;
        RECT 65.650 26.300 65.930 26.580 ;
        RECT 66.170 26.300 66.450 26.580 ;
        RECT 69.810 26.300 70.090 26.580 ;
        RECT 70.330 26.300 70.610 26.580 ;
        RECT 52.330 13.540 52.610 13.820 ;
        RECT 52.850 13.540 53.130 13.820 ;
        RECT 56.290 13.540 56.570 13.820 ;
        RECT 56.810 13.540 57.090 13.820 ;
        RECT 63.330 18.820 63.610 19.100 ;
        RECT 63.850 18.820 64.130 19.100 ;
        RECT 63.490 17.940 63.770 18.220 ;
        RECT 64.010 17.940 64.290 18.220 ;
        RECT 65.490 17.500 65.770 17.780 ;
        RECT 66.010 17.500 66.290 17.780 ;
        RECT 63.330 14.420 63.610 14.700 ;
        RECT 63.850 14.420 64.130 14.700 ;
        RECT 71.970 25.860 72.250 26.140 ;
        RECT 72.490 25.860 72.770 26.140 ;
        RECT 79.170 28.500 79.450 28.780 ;
        RECT 79.690 28.500 79.970 28.780 ;
        RECT 83.130 28.500 83.410 28.780 ;
        RECT 83.650 28.500 83.930 28.780 ;
        RECT 79.170 27.620 79.450 27.900 ;
        RECT 79.690 27.620 79.970 27.900 ;
        RECT 79.170 26.740 79.450 27.020 ;
        RECT 79.690 26.740 79.970 27.020 ;
        RECT 83.130 26.740 83.410 27.020 ;
        RECT 83.650 26.740 83.930 27.020 ;
        RECT 79.170 25.860 79.450 26.140 ;
        RECT 79.690 25.860 79.970 26.140 ;
        RECT 83.130 25.860 83.410 26.140 ;
        RECT 83.650 25.860 83.930 26.140 ;
        RECT 71.970 18.820 72.250 19.100 ;
        RECT 72.490 18.820 72.770 19.100 ;
        RECT 71.970 17.940 72.250 18.220 ;
        RECT 72.490 17.940 72.770 18.220 ;
        RECT 69.970 17.500 70.250 17.780 ;
        RECT 70.490 17.500 70.770 17.780 ;
        RECT 72.130 14.420 72.410 14.700 ;
        RECT 72.650 14.420 72.930 14.700 ;
        RECT 90.630 29.880 91.710 30.200 ;
        RECT 123.390 29.080 124.470 29.400 ;
        RECT 90.630 28.280 91.710 28.600 ;
        RECT 123.390 27.480 124.470 27.800 ;
        RECT 79.170 24.980 79.450 25.260 ;
        RECT 79.690 24.980 79.970 25.260 ;
        RECT 83.130 24.980 83.410 25.260 ;
        RECT 83.650 24.980 83.930 25.260 ;
        RECT 83.130 24.270 83.410 24.550 ;
        RECT 83.650 24.270 83.930 24.550 ;
        RECT 79.170 23.220 79.450 23.500 ;
        RECT 79.690 23.220 79.970 23.500 ;
        RECT 83.130 23.220 83.410 23.500 ;
        RECT 83.650 23.220 83.930 23.500 ;
        RECT 79.330 22.340 79.610 22.620 ;
        RECT 79.850 22.340 80.130 22.620 ;
        RECT 83.130 22.340 83.410 22.620 ;
        RECT 83.650 22.340 83.930 22.620 ;
        RECT 77.010 21.900 77.290 22.180 ;
        RECT 77.530 21.900 77.810 22.180 ;
        RECT 77.010 21.020 77.290 21.300 ;
        RECT 77.530 21.020 77.810 21.300 ;
        RECT 83.130 21.460 83.410 21.740 ;
        RECT 83.650 21.460 83.930 21.740 ;
        RECT 79.170 20.580 79.450 20.860 ;
        RECT 79.690 20.580 79.970 20.860 ;
        RECT 79.170 19.700 79.450 19.980 ;
        RECT 79.690 19.700 79.970 19.980 ;
        RECT 83.130 18.820 83.410 19.100 ;
        RECT 83.650 18.820 83.930 19.100 ;
        RECT 85.290 18.380 85.570 18.660 ;
        RECT 85.810 18.380 86.090 18.660 ;
        RECT 79.170 17.940 79.450 18.220 ;
        RECT 79.690 17.940 79.970 18.220 ;
        RECT 83.130 17.940 83.410 18.220 ;
        RECT 83.650 17.940 83.930 18.220 ;
        RECT 85.290 17.500 85.570 17.780 ;
        RECT 85.810 17.500 86.090 17.780 ;
        RECT 79.170 16.350 79.450 16.630 ;
        RECT 79.690 16.350 79.970 16.630 ;
        RECT 83.130 16.180 83.410 16.460 ;
        RECT 83.650 16.180 83.930 16.460 ;
        RECT 77.090 15.740 77.370 16.020 ;
        RECT 77.610 15.740 77.890 16.020 ;
        RECT 79.170 15.300 79.450 15.580 ;
        RECT 79.690 15.300 79.970 15.580 ;
        RECT 83.130 15.300 83.410 15.580 ;
        RECT 83.650 15.300 83.930 15.580 ;
        RECT 79.170 14.420 79.450 14.700 ;
        RECT 79.690 14.420 79.970 14.700 ;
        RECT 83.130 14.420 83.410 14.700 ;
        RECT 83.650 14.420 83.930 14.700 ;
        RECT 90.630 26.680 91.710 27.000 ;
        RECT 123.390 25.880 124.470 26.200 ;
        RECT 90.630 25.080 91.710 25.400 ;
        RECT 123.390 24.280 124.470 24.600 ;
        RECT 90.630 23.480 91.710 23.800 ;
        RECT 123.390 22.680 124.470 23.000 ;
        RECT 90.630 21.880 91.710 22.200 ;
        RECT 123.390 21.080 124.470 21.400 ;
        RECT 90.630 20.280 91.710 20.600 ;
        RECT 123.390 19.480 124.470 19.800 ;
        RECT 90.630 18.680 91.710 19.000 ;
        RECT 123.390 17.880 124.470 18.200 ;
        RECT 79.170 13.540 79.450 13.820 ;
        RECT 79.690 13.540 79.970 13.820 ;
        RECT 83.130 13.540 83.410 13.820 ;
        RECT 83.650 13.540 83.930 13.820 ;
        RECT 90.630 17.080 91.710 17.400 ;
        RECT 123.390 16.280 124.470 16.600 ;
        RECT 90.630 15.480 91.710 15.800 ;
        RECT 123.390 14.680 124.470 15.000 ;
        RECT 90.630 13.880 91.710 14.200 ;
        RECT 123.390 13.080 124.470 13.400 ;
        RECT 56.290 10.220 56.570 10.500 ;
        RECT 56.810 10.220 57.090 10.500 ;
        RECT 79.170 10.220 79.450 10.500 ;
        RECT 79.690 10.220 79.970 10.500 ;
        RECT 56.290 9.700 56.570 9.980 ;
        RECT 56.810 9.700 57.090 9.980 ;
        RECT 79.170 9.700 79.450 9.980 ;
        RECT 79.690 9.700 79.970 9.980 ;
        RECT 52.330 6.620 52.610 6.900 ;
        RECT 52.850 6.620 53.130 6.900 ;
        RECT 83.130 6.620 83.410 6.900 ;
        RECT 83.650 6.620 83.930 6.900 ;
        RECT 52.330 6.100 52.610 6.380 ;
        RECT 52.850 6.100 53.130 6.380 ;
        RECT 83.130 6.100 83.410 6.380 ;
        RECT 83.650 6.100 83.930 6.380 ;
        RECT 135.240 208.115 135.480 208.355 ;
        RECT 146.550 208.085 146.850 208.385 ;
        RECT 140.095 206.345 140.375 206.625 ;
        RECT 140.615 206.345 140.895 206.625 ;
        RECT 144.055 206.345 144.335 206.625 ;
        RECT 144.575 206.345 144.855 206.625 ;
        RECT 140.095 205.465 140.375 205.745 ;
        RECT 140.615 205.465 140.895 205.745 ;
        RECT 144.055 205.465 144.335 205.745 ;
        RECT 144.575 205.465 144.855 205.745 ;
        RECT 144.215 204.585 145.015 204.865 ;
        RECT 140.095 203.705 140.375 203.985 ;
        RECT 140.615 203.705 140.895 203.985 ;
        RECT 144.055 203.705 144.335 203.985 ;
        RECT 144.575 203.705 144.855 203.985 ;
        RECT 140.255 202.825 141.055 203.105 ;
        RECT 138.095 200.625 138.895 200.905 ;
        RECT 140.095 201.945 140.375 202.225 ;
        RECT 140.615 201.945 140.895 202.225 ;
        RECT 144.055 201.945 144.335 202.225 ;
        RECT 144.575 201.945 144.855 202.225 ;
        RECT 140.095 201.065 140.375 201.345 ;
        RECT 140.615 201.065 140.895 201.345 ;
        RECT 144.055 201.065 144.335 201.345 ;
        RECT 144.575 201.065 144.855 201.345 ;
        RECT 58.370 5.010 58.650 5.290 ;
        RECT 58.890 5.010 59.170 5.290 ;
        RECT 77.090 5.010 77.370 5.290 ;
        RECT 77.610 5.010 77.890 5.290 ;
        RECT 58.890 3.950 59.170 4.230 ;
        RECT 59.410 3.950 59.690 4.230 ;
        RECT 76.570 3.950 76.850 4.230 ;
        RECT 77.090 3.950 77.370 4.230 ;
      LAYER met1 ;
        RECT 59.665 224.020 60.450 224.320 ;
        RECT 36.790 223.570 37.090 223.600 ;
        RECT 61.210 223.570 61.510 224.490 ;
        RECT 136.410 223.960 136.770 224.380 ;
        RECT 36.790 223.270 61.510 223.570 ;
        RECT 111.980 223.320 112.280 223.350 ;
        RECT 36.790 223.240 37.090 223.270 ;
        RECT 111.980 223.020 112.970 223.320 ;
        RECT 111.980 222.990 112.280 223.020 ;
        RECT 135.180 222.960 135.540 223.380 ;
        RECT 86.850 222.410 116.830 222.710 ;
        RECT 116.190 221.200 117.110 221.540 ;
        RECT 15.390 220.320 16.310 220.660 ;
        RECT 19.270 220.320 20.990 220.660 ;
        RECT 15.310 219.440 16.230 219.780 ;
        RECT 19.270 219.440 20.190 219.780 ;
        RECT 13.150 218.120 14.870 218.460 ;
        RECT 14.530 215.820 14.870 218.120 ;
        RECT 20.650 217.580 20.990 220.320 ;
        RECT 27.270 220.320 28.990 220.660 ;
        RECT 31.950 220.320 32.870 220.660 ;
        RECT 40.590 220.320 41.510 220.660 ;
        RECT 44.470 220.320 46.190 220.660 ;
        RECT 27.270 217.580 27.610 220.320 ;
        RECT 28.070 219.440 28.990 219.780 ;
        RECT 32.030 219.440 32.950 219.780 ;
        RECT 40.510 219.440 41.430 219.780 ;
        RECT 44.470 219.440 45.390 219.780 ;
        RECT 20.650 217.240 22.350 217.580 ;
        RECT 25.910 217.240 27.610 217.580 ;
        RECT 33.390 218.120 35.110 218.460 ;
        RECT 38.350 218.120 40.070 218.460 ;
        RECT 15.310 216.800 16.230 217.140 ;
        RECT 19.270 216.800 20.190 217.140 ;
        RECT 28.070 216.800 28.990 217.140 ;
        RECT 32.030 216.800 32.950 217.140 ;
        RECT 33.390 215.820 33.730 218.120 ;
        RECT 14.530 215.480 23.150 215.820 ;
        RECT 20.650 214.600 22.350 214.940 ;
        RECT 15.310 214.160 16.230 214.500 ;
        RECT 19.270 214.160 20.190 214.500 ;
        RECT 20.650 213.620 20.990 214.600 ;
        RECT 19.270 213.280 20.990 213.620 ;
        RECT 13.150 212.840 14.870 213.180 ;
        RECT 14.530 211.860 14.870 212.840 ;
        RECT 15.310 212.400 16.230 212.740 ;
        RECT 19.270 212.400 20.190 212.740 ;
        RECT 14.530 211.520 16.230 211.860 ;
        RECT 20.650 210.540 20.990 213.280 ;
        RECT 22.810 211.420 23.150 215.480 ;
        RECT 21.430 211.080 23.150 211.420 ;
        RECT 20.650 210.200 22.350 210.540 ;
        RECT 15.310 209.760 16.230 210.100 ;
        RECT 19.270 209.760 20.190 210.100 ;
        RECT 13.150 208.440 14.230 208.780 ;
        RECT 13.930 208.100 14.870 208.440 ;
        RECT 13.230 207.560 14.150 207.900 ;
        RECT 14.530 204.820 14.870 208.100 ;
        RECT 15.310 207.120 16.230 207.460 ;
        RECT 19.270 207.120 20.190 207.460 ;
        RECT 15.310 205.360 16.230 205.700 ;
        RECT 19.270 205.360 20.190 205.700 ;
        RECT 22.810 204.820 23.150 211.080 ;
        RECT 14.530 204.480 16.230 204.820 ;
        RECT 19.270 204.480 23.150 204.820 ;
        RECT 25.110 215.480 33.730 215.820 ;
        RECT 39.730 215.820 40.070 218.120 ;
        RECT 45.850 217.580 46.190 220.320 ;
        RECT 52.470 220.320 54.190 220.660 ;
        RECT 57.150 220.320 58.070 220.660 ;
        RECT 65.790 220.320 66.710 220.660 ;
        RECT 69.670 220.320 71.390 220.660 ;
        RECT 52.470 217.580 52.810 220.320 ;
        RECT 53.270 219.440 54.190 219.780 ;
        RECT 57.230 219.440 58.150 219.780 ;
        RECT 65.710 219.440 66.630 219.780 ;
        RECT 69.670 219.440 70.590 219.780 ;
        RECT 45.850 217.240 47.550 217.580 ;
        RECT 51.110 217.240 52.810 217.580 ;
        RECT 58.590 218.120 60.310 218.460 ;
        RECT 63.550 218.120 65.270 218.460 ;
        RECT 40.510 216.800 41.430 217.140 ;
        RECT 44.470 216.800 45.390 217.140 ;
        RECT 53.270 216.800 54.190 217.140 ;
        RECT 57.230 216.800 58.150 217.140 ;
        RECT 58.590 215.820 58.930 218.120 ;
        RECT 39.730 215.480 48.350 215.820 ;
        RECT 25.110 211.420 25.450 215.480 ;
        RECT 25.910 214.600 27.610 214.940 ;
        RECT 27.270 213.620 27.610 214.600 ;
        RECT 45.850 214.600 47.550 214.940 ;
        RECT 28.070 214.160 28.990 214.500 ;
        RECT 32.030 214.160 32.950 214.500 ;
        RECT 40.510 214.160 41.430 214.500 ;
        RECT 44.470 214.160 45.390 214.500 ;
        RECT 45.850 213.620 46.190 214.600 ;
        RECT 27.270 213.280 28.990 213.620 ;
        RECT 44.470 213.280 46.190 213.620 ;
        RECT 25.110 211.080 26.830 211.420 ;
        RECT 25.110 204.820 25.450 211.080 ;
        RECT 27.270 210.540 27.610 213.280 ;
        RECT 33.390 212.840 35.110 213.180 ;
        RECT 38.350 212.840 40.070 213.180 ;
        RECT 28.070 212.400 28.990 212.740 ;
        RECT 32.030 212.400 32.950 212.740 ;
        RECT 33.390 211.860 33.730 212.840 ;
        RECT 32.030 211.520 33.730 211.860 ;
        RECT 39.730 211.860 40.070 212.840 ;
        RECT 40.510 212.400 41.430 212.740 ;
        RECT 44.470 212.400 45.390 212.740 ;
        RECT 39.730 211.520 41.430 211.860 ;
        RECT 25.910 210.200 27.610 210.540 ;
        RECT 45.850 210.540 46.190 213.280 ;
        RECT 48.010 211.420 48.350 215.480 ;
        RECT 46.630 211.080 48.350 211.420 ;
        RECT 45.850 210.200 47.550 210.540 ;
        RECT 28.070 209.760 28.990 210.100 ;
        RECT 32.030 209.760 32.950 210.100 ;
        RECT 40.510 209.760 41.430 210.100 ;
        RECT 44.470 209.760 45.390 210.100 ;
        RECT 34.030 208.440 35.110 208.780 ;
        RECT 38.350 208.440 39.430 208.780 ;
        RECT 33.390 208.100 34.330 208.440 ;
        RECT 39.130 208.100 40.070 208.440 ;
        RECT 28.070 207.120 28.990 207.460 ;
        RECT 32.030 207.120 32.950 207.460 ;
        RECT 28.070 205.360 28.990 205.700 ;
        RECT 32.030 205.360 32.950 205.700 ;
        RECT 33.390 204.820 33.730 208.100 ;
        RECT 34.110 207.560 35.030 207.900 ;
        RECT 38.430 207.560 39.350 207.900 ;
        RECT 25.110 204.480 28.990 204.820 ;
        RECT 32.030 204.480 33.730 204.820 ;
        RECT 39.730 204.820 40.070 208.100 ;
        RECT 40.510 207.120 41.430 207.460 ;
        RECT 44.470 207.120 45.390 207.460 ;
        RECT 40.510 205.360 41.430 205.700 ;
        RECT 44.470 205.360 45.390 205.700 ;
        RECT 48.010 204.820 48.350 211.080 ;
        RECT 39.730 204.480 41.430 204.820 ;
        RECT 44.470 204.480 48.350 204.820 ;
        RECT 50.310 215.480 58.930 215.820 ;
        RECT 64.930 215.820 65.270 218.120 ;
        RECT 71.050 217.580 71.390 220.320 ;
        RECT 77.670 220.320 79.390 220.660 ;
        RECT 82.350 220.320 83.270 220.660 ;
        RECT 90.990 220.320 91.910 220.660 ;
        RECT 94.870 220.320 96.590 220.660 ;
        RECT 77.670 217.580 78.010 220.320 ;
        RECT 78.470 219.440 79.390 219.780 ;
        RECT 82.430 219.440 83.350 219.780 ;
        RECT 90.910 219.440 91.830 219.780 ;
        RECT 94.870 219.440 95.790 219.780 ;
        RECT 71.050 217.240 72.750 217.580 ;
        RECT 76.310 217.240 78.010 217.580 ;
        RECT 83.790 218.120 85.510 218.460 ;
        RECT 88.750 218.120 90.470 218.460 ;
        RECT 65.710 216.800 66.630 217.140 ;
        RECT 69.670 216.800 70.590 217.140 ;
        RECT 78.470 216.800 79.390 217.140 ;
        RECT 82.430 216.800 83.350 217.140 ;
        RECT 83.790 215.820 84.130 218.120 ;
        RECT 64.930 215.480 73.550 215.820 ;
        RECT 50.310 211.420 50.650 215.480 ;
        RECT 51.110 214.600 52.810 214.940 ;
        RECT 52.470 213.620 52.810 214.600 ;
        RECT 71.050 214.600 72.750 214.940 ;
        RECT 53.270 214.160 54.190 214.500 ;
        RECT 57.230 214.160 58.150 214.500 ;
        RECT 65.710 214.160 66.630 214.500 ;
        RECT 69.670 214.160 70.590 214.500 ;
        RECT 71.050 213.620 71.390 214.600 ;
        RECT 52.470 213.280 54.190 213.620 ;
        RECT 69.670 213.280 71.390 213.620 ;
        RECT 50.310 211.080 52.030 211.420 ;
        RECT 50.310 204.820 50.650 211.080 ;
        RECT 52.470 210.540 52.810 213.280 ;
        RECT 58.590 212.840 60.310 213.180 ;
        RECT 63.550 212.840 65.270 213.180 ;
        RECT 53.270 212.400 54.190 212.740 ;
        RECT 57.230 212.400 58.150 212.740 ;
        RECT 58.590 211.860 58.930 212.840 ;
        RECT 57.230 211.520 58.930 211.860 ;
        RECT 64.930 211.860 65.270 212.840 ;
        RECT 65.710 212.400 66.630 212.740 ;
        RECT 69.670 212.400 70.590 212.740 ;
        RECT 64.930 211.520 66.630 211.860 ;
        RECT 51.110 210.200 52.810 210.540 ;
        RECT 71.050 210.540 71.390 213.280 ;
        RECT 73.210 211.420 73.550 215.480 ;
        RECT 71.830 211.080 73.550 211.420 ;
        RECT 71.050 210.200 72.750 210.540 ;
        RECT 53.270 209.760 54.190 210.100 ;
        RECT 57.230 209.760 58.150 210.100 ;
        RECT 65.710 209.760 66.630 210.100 ;
        RECT 69.670 209.760 70.590 210.100 ;
        RECT 59.230 208.440 60.310 208.780 ;
        RECT 63.550 208.440 64.630 208.780 ;
        RECT 58.590 208.100 59.530 208.440 ;
        RECT 64.330 208.100 65.270 208.440 ;
        RECT 53.270 207.120 54.190 207.460 ;
        RECT 57.230 207.120 58.150 207.460 ;
        RECT 53.270 205.360 54.190 205.700 ;
        RECT 57.230 205.360 58.150 205.700 ;
        RECT 58.590 204.820 58.930 208.100 ;
        RECT 59.310 207.560 60.230 207.900 ;
        RECT 63.630 207.560 64.550 207.900 ;
        RECT 50.310 204.480 54.190 204.820 ;
        RECT 57.230 204.480 58.930 204.820 ;
        RECT 64.930 204.820 65.270 208.100 ;
        RECT 65.710 207.120 66.630 207.460 ;
        RECT 69.670 207.120 70.590 207.460 ;
        RECT 65.710 205.360 66.630 205.700 ;
        RECT 69.670 205.360 70.590 205.700 ;
        RECT 73.210 204.820 73.550 211.080 ;
        RECT 64.930 204.480 66.630 204.820 ;
        RECT 69.670 204.480 73.550 204.820 ;
        RECT 75.510 215.480 84.130 215.820 ;
        RECT 90.130 215.820 90.470 218.120 ;
        RECT 96.250 217.580 96.590 220.320 ;
        RECT 102.870 220.320 104.590 220.660 ;
        RECT 107.550 220.320 108.470 220.660 ;
        RECT 116.110 220.320 117.030 220.660 ;
        RECT 120.070 220.320 120.990 220.660 ;
        RECT 102.870 217.580 103.210 220.320 ;
        RECT 103.670 219.440 104.590 219.780 ;
        RECT 107.630 219.440 108.550 219.780 ;
        RECT 116.110 219.440 117.030 219.780 ;
        RECT 133.260 219.770 133.660 219.830 ;
        RECT 132.500 219.430 133.660 219.770 ;
        RECT 133.260 219.370 133.660 219.430 ;
        RECT 116.110 218.560 117.030 218.900 ;
        RECT 120.070 218.560 120.990 218.900 ;
        RECT 96.250 217.240 97.950 217.580 ;
        RECT 101.510 217.240 103.210 217.580 ;
        RECT 108.990 218.120 110.710 218.460 ;
        RECT 90.910 216.800 91.830 217.140 ;
        RECT 94.870 216.800 95.790 217.140 ;
        RECT 103.670 216.800 104.590 217.140 ;
        RECT 107.630 216.800 108.550 217.140 ;
        RECT 108.990 215.820 109.330 218.120 ;
        RECT 120.070 217.680 120.990 218.020 ;
        RECT 113.950 217.240 117.830 217.580 ;
        RECT 114.110 216.360 115.030 216.700 ;
        RECT 116.110 215.920 117.030 216.260 ;
        RECT 90.130 215.480 98.750 215.820 ;
        RECT 75.510 211.420 75.850 215.480 ;
        RECT 76.310 214.600 78.010 214.940 ;
        RECT 77.670 213.620 78.010 214.600 ;
        RECT 96.250 214.600 97.950 214.940 ;
        RECT 78.470 214.160 79.390 214.500 ;
        RECT 82.430 214.160 83.350 214.500 ;
        RECT 90.910 214.160 91.830 214.500 ;
        RECT 94.870 214.160 95.790 214.500 ;
        RECT 96.250 213.620 96.590 214.600 ;
        RECT 77.670 213.280 79.390 213.620 ;
        RECT 94.870 213.280 96.590 213.620 ;
        RECT 75.510 211.080 77.230 211.420 ;
        RECT 75.510 204.820 75.850 211.080 ;
        RECT 77.670 210.540 78.010 213.280 ;
        RECT 83.790 212.840 85.510 213.180 ;
        RECT 88.750 212.840 90.470 213.180 ;
        RECT 78.470 212.400 79.390 212.740 ;
        RECT 82.430 212.400 83.350 212.740 ;
        RECT 83.790 211.860 84.130 212.840 ;
        RECT 82.430 211.520 84.130 211.860 ;
        RECT 90.130 211.860 90.470 212.840 ;
        RECT 90.910 212.400 91.830 212.740 ;
        RECT 94.870 212.400 95.790 212.740 ;
        RECT 90.130 211.520 91.830 211.860 ;
        RECT 76.310 210.200 78.010 210.540 ;
        RECT 96.250 210.540 96.590 213.280 ;
        RECT 98.410 211.420 98.750 215.480 ;
        RECT 97.030 211.080 98.750 211.420 ;
        RECT 96.250 210.200 97.950 210.540 ;
        RECT 78.470 209.760 79.390 210.100 ;
        RECT 82.430 209.760 83.350 210.100 ;
        RECT 90.910 209.760 91.830 210.100 ;
        RECT 94.870 209.760 95.790 210.100 ;
        RECT 84.430 208.440 85.510 208.780 ;
        RECT 88.750 208.440 89.830 208.780 ;
        RECT 83.790 208.100 84.730 208.440 ;
        RECT 89.530 208.100 90.470 208.440 ;
        RECT 78.470 207.120 79.390 207.460 ;
        RECT 82.430 207.120 83.350 207.460 ;
        RECT 78.470 205.360 79.390 205.700 ;
        RECT 82.430 205.360 83.350 205.700 ;
        RECT 83.790 204.820 84.130 208.100 ;
        RECT 84.510 207.560 85.430 207.900 ;
        RECT 88.830 207.560 89.750 207.900 ;
        RECT 75.510 204.480 79.390 204.820 ;
        RECT 82.430 204.480 84.130 204.820 ;
        RECT 90.130 204.820 90.470 208.100 ;
        RECT 90.910 207.120 91.830 207.460 ;
        RECT 94.870 207.120 95.790 207.460 ;
        RECT 90.910 205.360 91.830 205.700 ;
        RECT 94.870 205.360 95.790 205.700 ;
        RECT 98.410 204.820 98.750 211.080 ;
        RECT 90.130 204.480 91.830 204.820 ;
        RECT 94.870 204.480 98.750 204.820 ;
        RECT 100.710 215.480 109.330 215.820 ;
        RECT 100.710 211.420 101.050 215.480 ;
        RECT 116.110 215.040 117.030 215.380 ;
        RECT 101.510 214.600 103.210 214.940 ;
        RECT 102.870 213.620 103.210 214.600 ;
        RECT 103.670 214.160 104.590 214.500 ;
        RECT 107.630 214.160 108.550 214.500 ;
        RECT 116.110 214.160 117.030 214.500 ;
        RECT 102.870 213.280 104.590 213.620 ;
        RECT 116.110 213.280 117.030 213.620 ;
        RECT 100.710 211.080 102.430 211.420 ;
        RECT 100.710 204.820 101.050 211.080 ;
        RECT 102.870 210.540 103.210 213.280 ;
        RECT 108.990 212.840 110.710 213.180 ;
        RECT 103.670 212.400 104.590 212.740 ;
        RECT 107.630 212.400 108.550 212.740 ;
        RECT 108.990 211.860 109.330 212.840 ;
        RECT 116.110 212.400 117.030 212.740 ;
        RECT 107.630 211.520 109.330 211.860 ;
        RECT 116.110 211.520 117.030 211.860 ;
        RECT 113.950 211.080 115.670 211.420 ;
        RECT 101.510 210.200 103.210 210.540 ;
        RECT 114.110 210.200 115.030 210.540 ;
        RECT 103.670 209.760 104.590 210.100 ;
        RECT 107.630 209.760 108.550 210.100 ;
        RECT 109.630 208.440 110.710 208.780 ;
        RECT 108.990 208.100 109.930 208.440 ;
        RECT 103.670 207.120 104.590 207.460 ;
        RECT 107.630 207.120 108.550 207.460 ;
        RECT 103.670 205.360 104.590 205.700 ;
        RECT 107.630 205.360 108.550 205.700 ;
        RECT 108.990 204.820 109.330 208.100 ;
        RECT 109.710 207.560 110.630 207.900 ;
        RECT 113.950 207.560 114.870 207.900 ;
        RECT 115.330 206.140 115.670 211.080 ;
        RECT 116.110 209.760 117.030 210.100 ;
        RECT 116.270 208.880 117.190 209.220 ;
        RECT 116.110 208.000 117.030 208.340 ;
        RECT 117.490 206.580 117.830 217.240 ;
        RECT 120.070 215.920 120.990 216.260 ;
        RECT 120.070 214.160 120.990 214.500 ;
        RECT 120.070 212.400 120.990 212.740 ;
        RECT 120.070 209.760 120.990 210.100 ;
        RECT 120.070 208.000 120.990 208.340 ;
        RECT 116.110 206.240 117.830 206.580 ;
        RECT 113.950 205.800 115.670 206.140 ;
        RECT 100.710 204.480 104.590 204.820 ;
        RECT 107.630 204.480 109.330 204.820 ;
        RECT 115.330 204.820 115.670 205.800 ;
        RECT 116.110 205.360 117.030 205.700 ;
        RECT 120.070 205.360 120.990 205.700 ;
        RECT 115.330 204.480 117.030 204.820 ;
        RECT 13.230 204.040 14.150 204.380 ;
        RECT 34.110 204.040 35.030 204.380 ;
        RECT 38.430 204.040 39.350 204.380 ;
        RECT 59.310 204.040 60.230 204.380 ;
        RECT 63.630 204.040 64.550 204.380 ;
        RECT 84.510 204.040 85.430 204.380 ;
        RECT 88.830 204.040 89.750 204.380 ;
        RECT 109.710 204.040 110.630 204.380 ;
        RECT 114.110 204.040 115.030 204.380 ;
        RECT 13.520 200.850 13.860 204.040 ;
        RECT 15.310 203.600 16.230 203.940 ;
        RECT 19.270 203.600 20.190 203.940 ;
        RECT 28.070 203.600 28.990 203.940 ;
        RECT 32.030 203.600 32.950 203.940 ;
        RECT 15.310 202.720 16.230 203.060 ;
        RECT 19.270 202.720 20.190 203.060 ;
        RECT 28.070 202.720 28.990 203.060 ;
        RECT 32.030 202.720 32.950 203.060 ;
        RECT 15.310 201.840 16.230 202.180 ;
        RECT 19.270 201.840 20.190 202.180 ;
        RECT 28.070 201.840 28.990 202.180 ;
        RECT 32.030 201.840 32.950 202.180 ;
        RECT 34.400 200.850 34.740 204.040 ;
        RECT 38.720 200.850 39.060 204.040 ;
        RECT 40.510 203.600 41.430 203.940 ;
        RECT 44.470 203.600 45.390 203.940 ;
        RECT 53.270 203.600 54.190 203.940 ;
        RECT 57.230 203.600 58.150 203.940 ;
        RECT 40.510 202.720 41.430 203.060 ;
        RECT 44.470 202.720 45.390 203.060 ;
        RECT 53.270 202.720 54.190 203.060 ;
        RECT 57.230 202.720 58.150 203.060 ;
        RECT 40.510 201.840 41.430 202.180 ;
        RECT 44.470 201.840 45.390 202.180 ;
        RECT 53.270 201.840 54.190 202.180 ;
        RECT 57.230 201.840 58.150 202.180 ;
        RECT 59.600 200.850 59.940 204.040 ;
        RECT 63.920 200.850 64.260 204.040 ;
        RECT 65.710 203.600 66.630 203.940 ;
        RECT 69.670 203.600 70.590 203.940 ;
        RECT 78.470 203.600 79.390 203.940 ;
        RECT 82.430 203.600 83.350 203.940 ;
        RECT 65.710 202.720 66.630 203.060 ;
        RECT 69.670 202.720 70.590 203.060 ;
        RECT 78.470 202.720 79.390 203.060 ;
        RECT 82.430 202.720 83.350 203.060 ;
        RECT 65.710 201.840 66.630 202.180 ;
        RECT 69.670 201.840 70.590 202.180 ;
        RECT 78.470 201.840 79.390 202.180 ;
        RECT 82.430 201.840 83.350 202.180 ;
        RECT 84.800 200.850 85.140 204.040 ;
        RECT 89.120 200.850 89.460 204.040 ;
        RECT 90.910 203.600 91.830 203.940 ;
        RECT 94.870 203.600 95.790 203.940 ;
        RECT 103.670 203.600 104.590 203.940 ;
        RECT 107.630 203.600 108.550 203.940 ;
        RECT 90.910 202.720 91.830 203.060 ;
        RECT 94.870 202.720 95.790 203.060 ;
        RECT 103.670 202.720 104.590 203.060 ;
        RECT 107.630 202.720 108.550 203.060 ;
        RECT 90.910 201.840 91.830 202.180 ;
        RECT 94.870 201.840 95.790 202.180 ;
        RECT 103.670 201.840 104.590 202.180 ;
        RECT 107.630 201.840 108.550 202.180 ;
        RECT 110.000 200.850 110.340 204.040 ;
        RECT 116.110 203.600 117.030 203.940 ;
        RECT 120.070 203.600 120.990 203.940 ;
        RECT 116.110 202.720 117.030 203.060 ;
        RECT 120.070 202.720 120.990 203.060 ;
        RECT 116.110 201.840 117.030 202.180 ;
        RECT 120.070 201.840 120.990 202.180 ;
        RECT 13.230 200.510 14.150 200.850 ;
        RECT 34.110 200.510 35.030 200.850 ;
        RECT 38.430 200.510 39.350 200.850 ;
        RECT 59.310 200.510 60.230 200.850 ;
        RECT 63.630 200.510 64.550 200.850 ;
        RECT 84.510 200.510 85.430 200.850 ;
        RECT 88.830 200.510 89.750 200.850 ;
        RECT 109.710 200.510 110.630 200.850 ;
        RECT 111.830 200.170 112.170 200.900 ;
        RECT 15.310 199.070 16.230 199.990 ;
        RECT 32.030 199.070 32.950 199.990 ;
        RECT 40.510 199.070 41.430 199.990 ;
        RECT 57.230 199.070 58.150 199.990 ;
        RECT 65.710 199.070 66.630 199.990 ;
        RECT 82.430 199.070 83.350 199.990 ;
        RECT 90.910 199.070 91.830 199.990 ;
        RECT 107.630 199.070 108.550 199.990 ;
        RECT 111.800 199.830 112.200 200.170 ;
        RECT 116.110 199.070 117.030 199.990 ;
        RECT 19.270 197.630 20.190 198.550 ;
        RECT 22.050 197.630 22.970 198.550 ;
        RECT 25.090 197.630 26.010 198.550 ;
        RECT 28.070 197.630 28.990 198.550 ;
        RECT 44.470 197.630 45.390 198.550 ;
        RECT 47.250 197.630 48.170 198.550 ;
        RECT 50.290 197.630 51.210 198.550 ;
        RECT 53.270 197.630 54.190 198.550 ;
        RECT 69.670 197.630 70.590 198.550 ;
        RECT 72.450 197.630 73.370 198.550 ;
        RECT 75.490 197.630 76.410 198.550 ;
        RECT 78.470 197.630 79.390 198.550 ;
        RECT 94.870 197.630 95.790 198.550 ;
        RECT 97.650 197.630 98.570 198.550 ;
        RECT 100.690 197.630 101.610 198.550 ;
        RECT 103.670 197.630 104.590 198.550 ;
        RECT 120.070 197.630 120.990 198.550 ;
        RECT 19.170 194.030 20.090 194.950 ;
        RECT 27.970 194.030 28.890 194.950 ;
        RECT 44.370 194.030 45.290 194.950 ;
        RECT 53.170 194.030 54.090 194.950 ;
        RECT 69.570 194.030 70.490 194.950 ;
        RECT 78.370 194.030 79.290 194.950 ;
        RECT 94.770 194.030 95.690 194.950 ;
        RECT 103.570 194.030 104.490 194.950 ;
        RECT 119.970 194.030 120.890 194.950 ;
        RECT 15.210 190.430 16.130 191.350 ;
        RECT 31.930 190.430 32.850 191.350 ;
        RECT 40.410 190.430 41.330 191.350 ;
        RECT 57.130 190.430 58.050 191.350 ;
        RECT 65.610 190.430 66.530 191.350 ;
        RECT 82.330 190.430 83.250 191.350 ;
        RECT 90.810 190.430 91.730 191.350 ;
        RECT 107.530 190.430 108.450 191.350 ;
        RECT 116.010 190.430 116.930 191.350 ;
        RECT 15.210 187.140 16.130 187.480 ;
        RECT 19.170 187.140 20.090 187.480 ;
        RECT 27.970 187.140 28.890 187.480 ;
        RECT 31.930 187.140 32.850 187.480 ;
        RECT 40.410 187.140 41.330 187.480 ;
        RECT 44.370 187.140 45.290 187.480 ;
        RECT 53.170 187.140 54.090 187.480 ;
        RECT 57.130 187.140 58.050 187.480 ;
        RECT 65.610 187.140 66.530 187.480 ;
        RECT 69.570 187.140 70.490 187.480 ;
        RECT 78.370 187.140 79.290 187.480 ;
        RECT 82.330 187.140 83.250 187.480 ;
        RECT 90.810 187.140 91.730 187.480 ;
        RECT 94.770 187.140 95.690 187.480 ;
        RECT 103.570 187.140 104.490 187.480 ;
        RECT 107.530 187.140 108.450 187.480 ;
        RECT 15.210 186.260 16.130 186.600 ;
        RECT 19.170 186.260 20.090 186.600 ;
        RECT 27.970 186.260 28.890 186.600 ;
        RECT 31.930 186.260 32.850 186.600 ;
        RECT 40.410 186.260 41.330 186.600 ;
        RECT 44.370 186.260 45.290 186.600 ;
        RECT 53.170 186.260 54.090 186.600 ;
        RECT 57.130 186.260 58.050 186.600 ;
        RECT 65.610 186.260 66.530 186.600 ;
        RECT 69.570 186.260 70.490 186.600 ;
        RECT 78.370 186.260 79.290 186.600 ;
        RECT 82.330 186.260 83.250 186.600 ;
        RECT 90.810 186.260 91.730 186.600 ;
        RECT 94.770 186.260 95.690 186.600 ;
        RECT 103.570 186.260 104.490 186.600 ;
        RECT 107.530 186.260 108.450 186.600 ;
        RECT 19.170 185.550 20.090 185.890 ;
        RECT 27.810 185.380 29.830 185.720 ;
        RECT 44.370 185.550 45.290 185.890 ;
        RECT 53.010 185.380 55.030 185.720 ;
        RECT 69.570 185.550 70.490 185.890 ;
        RECT 78.210 185.380 80.230 185.720 ;
        RECT 94.770 185.550 95.690 185.890 ;
        RECT 103.410 185.380 104.330 185.720 ;
        RECT 15.210 184.500 16.130 184.840 ;
        RECT 19.170 184.500 20.090 184.840 ;
        RECT 27.970 184.500 28.890 184.840 ;
        RECT 2.630 183.520 2.970 183.810 ;
        RECT 15.210 183.620 16.130 183.960 ;
        RECT 2.630 183.180 13.970 183.520 ;
        RECT 2.630 182.890 2.970 183.180 ;
        RECT 29.490 182.880 29.830 185.380 ;
        RECT 31.930 184.500 32.850 184.840 ;
        RECT 40.410 184.500 41.330 184.840 ;
        RECT 44.370 184.500 45.290 184.840 ;
        RECT 53.170 184.500 54.090 184.840 ;
        RECT 31.930 183.620 32.850 183.960 ;
        RECT 40.410 183.620 41.330 183.960 ;
        RECT 33.930 183.180 34.850 183.520 ;
        RECT 37.910 183.180 39.170 183.520 ;
        RECT 37.910 182.880 38.250 183.180 ;
        RECT 29.490 182.540 38.250 182.880 ;
        RECT 54.690 182.880 55.030 185.380 ;
        RECT 57.130 184.500 58.050 184.840 ;
        RECT 65.610 184.500 66.530 184.840 ;
        RECT 69.570 184.500 70.490 184.840 ;
        RECT 78.370 184.500 79.290 184.840 ;
        RECT 57.130 183.620 58.050 183.960 ;
        RECT 65.610 183.620 66.530 183.960 ;
        RECT 59.130 183.180 60.050 183.520 ;
        RECT 63.110 183.180 64.370 183.520 ;
        RECT 63.110 182.880 63.450 183.180 ;
        RECT 54.690 182.540 63.450 182.880 ;
        RECT 79.890 182.880 80.230 185.380 ;
        RECT 82.330 184.500 83.250 184.840 ;
        RECT 90.810 184.500 91.730 184.840 ;
        RECT 94.770 184.500 95.690 184.840 ;
        RECT 103.570 184.500 104.490 184.840 ;
        RECT 107.530 184.500 108.450 184.840 ;
        RECT 82.330 183.620 83.250 183.960 ;
        RECT 90.810 183.620 91.730 183.960 ;
        RECT 107.530 183.620 108.450 183.960 ;
        RECT 84.330 183.180 85.250 183.520 ;
        RECT 88.310 183.180 89.570 183.520 ;
        RECT 109.530 183.180 110.450 183.520 ;
        RECT 88.310 182.880 88.650 183.180 ;
        RECT 79.890 182.540 88.650 182.880 ;
        RECT 116.010 182.740 116.930 183.080 ;
        RECT 119.970 182.740 120.890 183.080 ;
        RECT 15.210 181.860 16.130 182.200 ;
        RECT 19.170 181.860 20.090 182.200 ;
        RECT 27.970 181.860 28.890 182.200 ;
        RECT 31.930 181.860 32.850 182.200 ;
        RECT 40.410 181.860 41.330 182.200 ;
        RECT 44.370 181.860 45.290 182.200 ;
        RECT 53.170 181.860 54.090 182.200 ;
        RECT 57.130 181.860 58.050 182.200 ;
        RECT 65.610 181.860 66.530 182.200 ;
        RECT 69.570 181.860 70.490 182.200 ;
        RECT 78.370 181.860 79.290 182.200 ;
        RECT 82.330 181.860 83.250 182.200 ;
        RECT 90.810 181.860 91.730 182.200 ;
        RECT 94.770 181.860 95.690 182.200 ;
        RECT 103.570 181.860 104.490 182.200 ;
        RECT 107.530 181.860 108.450 182.200 ;
        RECT 116.010 181.860 116.930 182.200 ;
        RECT 119.970 181.860 120.890 182.200 ;
        RECT 113.850 180.710 114.770 181.050 ;
        RECT 15.210 180.100 16.130 180.440 ;
        RECT 19.170 180.100 20.090 180.440 ;
        RECT 27.970 180.100 28.890 180.440 ;
        RECT 31.930 180.100 32.850 180.440 ;
        RECT 40.410 180.100 41.330 180.440 ;
        RECT 44.370 180.100 45.290 180.440 ;
        RECT 53.170 180.100 54.090 180.440 ;
        RECT 57.130 180.100 58.050 180.440 ;
        RECT 65.610 180.100 66.530 180.440 ;
        RECT 69.570 180.100 70.490 180.440 ;
        RECT 78.370 180.100 79.290 180.440 ;
        RECT 82.330 180.100 83.250 180.440 ;
        RECT 90.810 180.100 91.730 180.440 ;
        RECT 94.770 180.100 95.690 180.440 ;
        RECT 103.570 180.100 104.490 180.440 ;
        RECT 107.530 180.100 108.450 180.440 ;
        RECT 116.010 180.100 116.930 180.440 ;
        RECT 119.970 180.100 120.890 180.440 ;
        RECT 19.170 179.220 20.090 179.560 ;
        RECT 27.970 179.220 28.890 179.560 ;
        RECT 44.370 179.220 45.290 179.560 ;
        RECT 53.170 179.220 54.090 179.560 ;
        RECT 69.570 179.220 70.490 179.560 ;
        RECT 78.370 179.220 79.290 179.560 ;
        RECT 94.770 179.220 95.690 179.560 ;
        RECT 103.570 179.220 104.490 179.560 ;
        RECT 116.010 179.220 116.930 179.560 ;
        RECT 13.050 178.780 14.770 179.120 ;
        RECT 14.430 173.400 14.770 178.780 ;
        RECT 33.290 178.780 35.010 179.120 ;
        RECT 38.250 178.780 39.970 179.120 ;
        RECT 15.210 177.460 16.130 177.800 ;
        RECT 19.170 177.460 20.090 177.800 ;
        RECT 27.970 177.460 28.890 177.800 ;
        RECT 31.930 177.460 32.850 177.800 ;
        RECT 15.210 176.580 16.130 176.920 ;
        RECT 31.770 176.580 32.690 176.920 ;
        RECT 15.210 175.700 16.130 176.040 ;
        RECT 19.170 175.700 20.090 176.040 ;
        RECT 27.970 175.700 28.890 176.040 ;
        RECT 31.930 175.700 32.850 176.040 ;
        RECT 21.330 174.380 23.050 174.720 ;
        RECT 15.210 173.940 16.130 174.280 ;
        RECT 19.170 173.940 20.090 174.280 ;
        RECT 14.430 173.060 16.130 173.400 ;
        RECT 20.550 171.740 22.250 172.080 ;
        RECT 15.210 171.300 16.130 171.640 ;
        RECT 19.170 171.300 20.090 171.640 ;
        RECT 13.050 170.860 13.970 171.200 ;
        RECT 15.210 169.540 16.130 169.880 ;
        RECT 15.210 168.660 16.130 169.000 ;
        RECT 19.170 168.660 20.090 169.000 ;
        RECT 15.210 166.900 16.130 167.240 ;
        RECT 19.170 166.900 20.090 167.240 ;
        RECT 18.160 165.730 18.500 166.650 ;
        RECT 15.210 165.140 16.130 165.480 ;
        RECT 19.170 165.140 20.090 165.480 ;
        RECT 15.210 164.260 16.130 164.600 ;
        RECT 19.170 164.260 20.090 164.600 ;
        RECT 15.210 162.500 16.130 162.840 ;
        RECT 19.170 162.500 20.090 162.840 ;
        RECT 13.050 161.180 14.770 161.520 ;
        RECT 17.375 161.330 17.715 162.250 ;
        RECT 13.210 156.780 14.130 157.120 ;
        RECT 12.410 150.620 13.970 150.960 ;
        RECT 12.410 147.440 12.750 150.620 ;
        RECT 13.050 148.860 13.970 149.200 ;
        RECT 14.430 147.880 14.770 161.180 ;
        RECT 15.210 160.740 16.130 161.080 ;
        RECT 19.170 160.740 20.090 161.080 ;
        RECT 15.210 159.860 16.130 160.200 ;
        RECT 19.170 159.860 20.090 160.200 ;
        RECT 15.210 158.100 16.130 158.440 ;
        RECT 19.170 158.100 20.090 158.440 ;
        RECT 16.660 156.930 17.000 157.850 ;
        RECT 20.550 157.560 20.890 171.740 ;
        RECT 19.170 157.220 20.890 157.560 ;
        RECT 15.210 156.340 16.130 156.680 ;
        RECT 19.170 156.340 20.090 156.680 ;
        RECT 15.210 155.460 16.130 155.800 ;
        RECT 19.170 155.460 20.090 155.800 ;
        RECT 15.210 153.700 16.130 154.040 ;
        RECT 19.170 153.700 20.090 154.040 ;
        RECT 15.210 151.940 16.130 152.280 ;
        RECT 19.170 151.940 20.090 152.280 ;
        RECT 21.330 150.620 22.250 150.960 ;
        RECT 15.210 148.420 16.130 148.760 ;
        RECT 19.170 148.420 20.090 148.760 ;
        RECT 14.430 147.540 16.130 147.880 ;
        RECT 12.410 147.100 13.970 147.440 ;
        RECT 12.410 136.880 12.750 147.100 ;
        RECT 13.210 145.340 14.770 145.680 ;
        RECT 14.430 140.400 14.770 145.340 ;
        RECT 15.210 144.900 16.130 145.240 ;
        RECT 19.170 144.900 20.090 145.240 ;
        RECT 15.210 143.140 16.130 143.480 ;
        RECT 19.170 143.140 20.090 143.480 ;
        RECT 19.170 142.260 20.090 142.600 ;
        RECT 15.210 141.380 16.130 141.720 ;
        RECT 15.210 140.500 16.130 140.840 ;
        RECT 13.210 140.060 14.770 140.400 ;
        RECT 22.710 138.200 23.050 174.380 ;
        RECT 15.210 137.860 16.130 138.200 ;
        RECT 19.170 137.860 23.050 138.200 ;
        RECT 25.010 174.380 26.730 174.720 ;
        RECT 25.010 138.200 25.350 174.380 ;
        RECT 27.970 173.940 28.890 174.280 ;
        RECT 31.930 173.940 32.850 174.280 ;
        RECT 33.290 173.400 33.630 178.780 ;
        RECT 31.930 173.060 33.630 173.400 ;
        RECT 39.630 173.400 39.970 178.780 ;
        RECT 58.490 178.780 60.210 179.120 ;
        RECT 63.450 178.780 65.170 179.120 ;
        RECT 40.410 177.460 41.330 177.800 ;
        RECT 44.370 177.460 45.290 177.800 ;
        RECT 53.170 177.460 54.090 177.800 ;
        RECT 57.130 177.460 58.050 177.800 ;
        RECT 40.410 176.580 41.330 176.920 ;
        RECT 56.970 176.580 57.890 176.920 ;
        RECT 40.410 175.700 41.330 176.040 ;
        RECT 44.370 175.700 45.290 176.040 ;
        RECT 53.170 175.700 54.090 176.040 ;
        RECT 57.130 175.700 58.050 176.040 ;
        RECT 46.530 174.380 48.250 174.720 ;
        RECT 40.410 173.940 41.330 174.280 ;
        RECT 44.370 173.940 45.290 174.280 ;
        RECT 39.630 173.060 41.330 173.400 ;
        RECT 25.810 171.740 27.510 172.080 ;
        RECT 27.170 157.560 27.510 171.740 ;
        RECT 45.750 171.740 47.450 172.080 ;
        RECT 27.970 171.300 28.890 171.640 ;
        RECT 31.930 171.300 32.850 171.640 ;
        RECT 40.410 171.300 41.330 171.640 ;
        RECT 44.370 171.300 45.290 171.640 ;
        RECT 33.930 170.860 34.850 171.200 ;
        RECT 38.250 170.860 39.170 171.200 ;
        RECT 31.930 169.540 32.850 169.880 ;
        RECT 40.410 169.540 41.330 169.880 ;
        RECT 27.970 168.660 28.890 169.000 ;
        RECT 31.930 168.660 32.850 169.000 ;
        RECT 40.410 168.660 41.330 169.000 ;
        RECT 44.370 168.660 45.290 169.000 ;
        RECT 27.970 166.900 28.890 167.240 ;
        RECT 31.930 166.900 32.850 167.240 ;
        RECT 40.410 166.900 41.330 167.240 ;
        RECT 44.370 166.900 45.290 167.240 ;
        RECT 29.560 165.730 29.900 166.650 ;
        RECT 43.360 165.730 43.700 166.650 ;
        RECT 27.970 165.140 28.890 165.480 ;
        RECT 31.930 165.140 32.850 165.480 ;
        RECT 40.410 165.140 41.330 165.480 ;
        RECT 44.370 165.140 45.290 165.480 ;
        RECT 27.970 164.260 28.890 164.600 ;
        RECT 31.930 164.260 32.850 164.600 ;
        RECT 40.410 164.260 41.330 164.600 ;
        RECT 44.370 164.260 45.290 164.600 ;
        RECT 27.970 162.500 28.890 162.840 ;
        RECT 31.930 162.500 32.850 162.840 ;
        RECT 40.410 162.500 41.330 162.840 ;
        RECT 44.370 162.500 45.290 162.840 ;
        RECT 30.345 161.330 30.685 162.250 ;
        RECT 33.290 161.180 35.010 161.520 ;
        RECT 38.250 161.180 39.970 161.520 ;
        RECT 42.575 161.330 42.915 162.250 ;
        RECT 27.970 160.740 28.890 161.080 ;
        RECT 31.930 160.740 32.850 161.080 ;
        RECT 27.970 159.860 28.890 160.200 ;
        RECT 31.930 159.860 32.850 160.200 ;
        RECT 27.970 158.100 28.890 158.440 ;
        RECT 31.930 158.100 32.850 158.440 ;
        RECT 27.170 157.220 28.890 157.560 ;
        RECT 31.060 156.930 31.400 157.850 ;
        RECT 27.970 156.340 28.890 156.680 ;
        RECT 31.930 156.340 32.850 156.680 ;
        RECT 27.970 155.460 28.890 155.800 ;
        RECT 31.930 155.460 32.850 155.800 ;
        RECT 27.970 153.700 28.890 154.040 ;
        RECT 31.930 153.700 32.850 154.040 ;
        RECT 27.970 151.940 28.890 152.280 ;
        RECT 31.930 151.940 32.850 152.280 ;
        RECT 25.650 150.620 26.570 150.960 ;
        RECT 27.970 148.420 28.890 148.760 ;
        RECT 31.930 148.420 32.850 148.760 ;
        RECT 33.290 147.880 33.630 161.180 ;
        RECT 33.930 156.780 34.850 157.120 ;
        RECT 38.410 156.780 39.330 157.120 ;
        RECT 34.090 150.620 35.650 150.960 ;
        RECT 33.930 148.860 34.850 149.200 ;
        RECT 31.930 147.540 33.630 147.880 ;
        RECT 35.310 147.440 35.650 150.620 ;
        RECT 34.090 147.100 35.650 147.440 ;
        RECT 33.290 145.340 34.850 145.680 ;
        RECT 27.970 144.900 28.890 145.240 ;
        RECT 31.930 144.900 32.850 145.240 ;
        RECT 27.970 143.140 28.890 143.480 ;
        RECT 31.930 143.140 32.850 143.480 ;
        RECT 27.970 142.260 28.890 142.600 ;
        RECT 31.930 141.380 32.850 141.720 ;
        RECT 31.930 140.500 32.850 140.840 ;
        RECT 33.290 140.400 33.630 145.340 ;
        RECT 33.290 140.060 34.850 140.400 ;
        RECT 25.010 137.860 28.890 138.200 ;
        RECT 31.930 137.860 32.850 138.200 ;
        RECT 19.170 136.980 20.090 137.320 ;
        RECT 27.970 136.980 28.890 137.320 ;
        RECT 35.310 136.880 35.650 147.100 ;
        RECT 12.410 136.540 14.130 136.880 ;
        RECT 33.930 136.540 35.650 136.880 ;
        RECT 37.610 150.620 39.170 150.960 ;
        RECT 37.610 147.440 37.950 150.620 ;
        RECT 38.250 148.860 39.170 149.200 ;
        RECT 39.630 147.880 39.970 161.180 ;
        RECT 40.410 160.740 41.330 161.080 ;
        RECT 44.370 160.740 45.290 161.080 ;
        RECT 40.410 159.860 41.330 160.200 ;
        RECT 44.370 159.860 45.290 160.200 ;
        RECT 40.410 158.100 41.330 158.440 ;
        RECT 44.370 158.100 45.290 158.440 ;
        RECT 41.860 156.930 42.200 157.850 ;
        RECT 45.750 157.560 46.090 171.740 ;
        RECT 44.370 157.220 46.090 157.560 ;
        RECT 40.410 156.340 41.330 156.680 ;
        RECT 44.370 156.340 45.290 156.680 ;
        RECT 40.410 155.460 41.330 155.800 ;
        RECT 44.370 155.460 45.290 155.800 ;
        RECT 40.410 153.700 41.330 154.040 ;
        RECT 44.370 153.700 45.290 154.040 ;
        RECT 40.410 151.940 41.330 152.280 ;
        RECT 44.370 151.940 45.290 152.280 ;
        RECT 46.530 150.620 47.450 150.960 ;
        RECT 40.410 148.420 41.330 148.760 ;
        RECT 44.370 148.420 45.290 148.760 ;
        RECT 39.630 147.540 41.330 147.880 ;
        RECT 37.610 147.100 39.170 147.440 ;
        RECT 37.610 136.880 37.950 147.100 ;
        RECT 38.410 145.340 39.970 145.680 ;
        RECT 39.630 140.400 39.970 145.340 ;
        RECT 40.410 144.900 41.330 145.240 ;
        RECT 44.370 144.900 45.290 145.240 ;
        RECT 40.410 143.140 41.330 143.480 ;
        RECT 44.370 143.140 45.290 143.480 ;
        RECT 44.370 142.260 45.290 142.600 ;
        RECT 40.410 141.380 41.330 141.720 ;
        RECT 40.410 140.500 41.330 140.840 ;
        RECT 38.410 140.060 39.970 140.400 ;
        RECT 47.910 138.200 48.250 174.380 ;
        RECT 40.410 137.860 41.330 138.200 ;
        RECT 44.370 137.860 48.250 138.200 ;
        RECT 50.210 174.380 51.930 174.720 ;
        RECT 50.210 138.200 50.550 174.380 ;
        RECT 53.170 173.940 54.090 174.280 ;
        RECT 57.130 173.940 58.050 174.280 ;
        RECT 58.490 173.400 58.830 178.780 ;
        RECT 57.130 173.060 58.830 173.400 ;
        RECT 64.830 173.400 65.170 178.780 ;
        RECT 83.690 178.780 85.410 179.120 ;
        RECT 88.650 178.780 90.370 179.120 ;
        RECT 65.610 177.460 66.530 177.800 ;
        RECT 69.570 177.460 70.490 177.800 ;
        RECT 78.370 177.460 79.290 177.800 ;
        RECT 82.330 177.460 83.250 177.800 ;
        RECT 65.610 176.580 66.530 176.920 ;
        RECT 82.170 176.580 83.090 176.920 ;
        RECT 65.610 175.700 66.530 176.040 ;
        RECT 69.570 175.700 70.490 176.040 ;
        RECT 78.370 175.700 79.290 176.040 ;
        RECT 82.330 175.700 83.250 176.040 ;
        RECT 71.730 174.380 73.450 174.720 ;
        RECT 65.610 173.940 66.530 174.280 ;
        RECT 69.570 173.940 70.490 174.280 ;
        RECT 64.830 173.060 66.530 173.400 ;
        RECT 51.010 171.740 52.710 172.080 ;
        RECT 52.370 157.560 52.710 171.740 ;
        RECT 70.950 171.740 72.650 172.080 ;
        RECT 53.170 171.300 54.090 171.640 ;
        RECT 57.130 171.300 58.050 171.640 ;
        RECT 65.610 171.300 66.530 171.640 ;
        RECT 69.570 171.300 70.490 171.640 ;
        RECT 59.130 170.860 60.050 171.200 ;
        RECT 63.450 170.860 64.370 171.200 ;
        RECT 57.130 169.540 58.050 169.880 ;
        RECT 65.610 169.540 66.530 169.880 ;
        RECT 53.170 168.660 54.090 169.000 ;
        RECT 57.130 168.660 58.050 169.000 ;
        RECT 65.610 168.660 66.530 169.000 ;
        RECT 69.570 168.660 70.490 169.000 ;
        RECT 53.170 166.900 54.090 167.240 ;
        RECT 57.130 166.900 58.050 167.240 ;
        RECT 65.610 166.900 66.530 167.240 ;
        RECT 69.570 166.900 70.490 167.240 ;
        RECT 54.760 165.730 55.100 166.650 ;
        RECT 68.560 165.730 68.900 166.650 ;
        RECT 53.170 165.140 54.090 165.480 ;
        RECT 57.130 165.140 58.050 165.480 ;
        RECT 65.610 165.140 66.530 165.480 ;
        RECT 69.570 165.140 70.490 165.480 ;
        RECT 53.170 164.260 54.090 164.600 ;
        RECT 57.130 164.260 58.050 164.600 ;
        RECT 65.610 164.260 66.530 164.600 ;
        RECT 69.570 164.260 70.490 164.600 ;
        RECT 53.170 162.500 54.090 162.840 ;
        RECT 57.130 162.500 58.050 162.840 ;
        RECT 65.610 162.500 66.530 162.840 ;
        RECT 69.570 162.500 70.490 162.840 ;
        RECT 55.545 161.330 55.885 162.250 ;
        RECT 58.490 161.180 60.210 161.520 ;
        RECT 63.450 161.180 65.170 161.520 ;
        RECT 67.775 161.330 68.115 162.250 ;
        RECT 53.170 160.740 54.090 161.080 ;
        RECT 57.130 160.740 58.050 161.080 ;
        RECT 53.170 159.860 54.090 160.200 ;
        RECT 57.130 159.860 58.050 160.200 ;
        RECT 53.170 158.100 54.090 158.440 ;
        RECT 57.130 158.100 58.050 158.440 ;
        RECT 52.370 157.220 54.090 157.560 ;
        RECT 56.260 156.930 56.600 157.850 ;
        RECT 53.170 156.340 54.090 156.680 ;
        RECT 57.130 156.340 58.050 156.680 ;
        RECT 53.170 155.460 54.090 155.800 ;
        RECT 57.130 155.460 58.050 155.800 ;
        RECT 53.170 153.700 54.090 154.040 ;
        RECT 57.130 153.700 58.050 154.040 ;
        RECT 53.170 151.940 54.090 152.280 ;
        RECT 57.130 151.940 58.050 152.280 ;
        RECT 50.850 150.620 51.770 150.960 ;
        RECT 53.170 148.420 54.090 148.760 ;
        RECT 57.130 148.420 58.050 148.760 ;
        RECT 58.490 147.880 58.830 161.180 ;
        RECT 59.130 156.780 60.050 157.120 ;
        RECT 63.610 156.780 64.530 157.120 ;
        RECT 59.290 150.620 60.850 150.960 ;
        RECT 59.130 148.860 60.050 149.200 ;
        RECT 57.130 147.540 58.830 147.880 ;
        RECT 60.510 147.440 60.850 150.620 ;
        RECT 59.290 147.100 60.850 147.440 ;
        RECT 58.490 145.340 60.050 145.680 ;
        RECT 53.170 144.900 54.090 145.240 ;
        RECT 57.130 144.900 58.050 145.240 ;
        RECT 53.170 143.140 54.090 143.480 ;
        RECT 57.130 143.140 58.050 143.480 ;
        RECT 53.170 142.260 54.090 142.600 ;
        RECT 57.130 141.380 58.050 141.720 ;
        RECT 57.130 140.500 58.050 140.840 ;
        RECT 58.490 140.400 58.830 145.340 ;
        RECT 58.490 140.060 60.050 140.400 ;
        RECT 50.210 137.860 54.090 138.200 ;
        RECT 57.130 137.860 58.050 138.200 ;
        RECT 44.370 136.980 45.290 137.320 ;
        RECT 53.170 136.980 54.090 137.320 ;
        RECT 60.510 136.880 60.850 147.100 ;
        RECT 37.610 136.540 39.330 136.880 ;
        RECT 59.130 136.540 60.850 136.880 ;
        RECT 62.810 150.620 64.370 150.960 ;
        RECT 62.810 147.440 63.150 150.620 ;
        RECT 63.450 148.860 64.370 149.200 ;
        RECT 64.830 147.880 65.170 161.180 ;
        RECT 65.610 160.740 66.530 161.080 ;
        RECT 69.570 160.740 70.490 161.080 ;
        RECT 65.610 159.860 66.530 160.200 ;
        RECT 69.570 159.860 70.490 160.200 ;
        RECT 65.610 158.100 66.530 158.440 ;
        RECT 69.570 158.100 70.490 158.440 ;
        RECT 67.060 156.930 67.400 157.850 ;
        RECT 70.950 157.560 71.290 171.740 ;
        RECT 69.570 157.220 71.290 157.560 ;
        RECT 65.610 156.340 66.530 156.680 ;
        RECT 69.570 156.340 70.490 156.680 ;
        RECT 65.610 155.460 66.530 155.800 ;
        RECT 69.570 155.460 70.490 155.800 ;
        RECT 65.610 153.700 66.530 154.040 ;
        RECT 69.570 153.700 70.490 154.040 ;
        RECT 65.610 151.940 66.530 152.280 ;
        RECT 69.570 151.940 70.490 152.280 ;
        RECT 71.730 150.620 72.650 150.960 ;
        RECT 65.610 148.420 66.530 148.760 ;
        RECT 69.570 148.420 70.490 148.760 ;
        RECT 64.830 147.540 66.530 147.880 ;
        RECT 62.810 147.100 64.370 147.440 ;
        RECT 62.810 136.880 63.150 147.100 ;
        RECT 63.610 145.340 65.170 145.680 ;
        RECT 64.830 140.400 65.170 145.340 ;
        RECT 65.610 144.900 66.530 145.240 ;
        RECT 69.570 144.900 70.490 145.240 ;
        RECT 65.610 143.140 66.530 143.480 ;
        RECT 69.570 143.140 70.490 143.480 ;
        RECT 69.570 142.260 70.490 142.600 ;
        RECT 65.610 141.380 66.530 141.720 ;
        RECT 65.610 140.500 66.530 140.840 ;
        RECT 63.610 140.060 65.170 140.400 ;
        RECT 73.110 138.200 73.450 174.380 ;
        RECT 65.610 137.860 66.530 138.200 ;
        RECT 69.570 137.860 73.450 138.200 ;
        RECT 75.410 174.380 77.130 174.720 ;
        RECT 75.410 138.200 75.750 174.380 ;
        RECT 78.370 173.940 79.290 174.280 ;
        RECT 82.330 173.940 83.250 174.280 ;
        RECT 83.690 173.400 84.030 178.780 ;
        RECT 82.330 173.060 84.030 173.400 ;
        RECT 90.030 173.400 90.370 178.780 ;
        RECT 108.890 178.780 110.610 179.120 ;
        RECT 113.850 178.780 114.770 179.120 ;
        RECT 90.810 177.460 91.730 177.800 ;
        RECT 94.770 177.460 95.690 177.800 ;
        RECT 103.570 177.460 104.490 177.800 ;
        RECT 107.530 177.460 108.450 177.800 ;
        RECT 90.810 176.580 91.730 176.920 ;
        RECT 107.370 176.580 108.290 176.920 ;
        RECT 90.810 175.700 91.730 176.040 ;
        RECT 94.770 175.700 95.690 176.040 ;
        RECT 103.570 175.700 104.490 176.040 ;
        RECT 107.530 175.700 108.450 176.040 ;
        RECT 96.930 174.380 98.650 174.720 ;
        RECT 90.810 173.940 91.730 174.280 ;
        RECT 94.770 173.940 95.690 174.280 ;
        RECT 90.030 173.060 91.730 173.400 ;
        RECT 76.210 171.740 77.910 172.080 ;
        RECT 77.570 157.560 77.910 171.740 ;
        RECT 96.150 171.740 97.850 172.080 ;
        RECT 78.370 171.300 79.290 171.640 ;
        RECT 82.330 171.300 83.250 171.640 ;
        RECT 90.810 171.300 91.730 171.640 ;
        RECT 94.770 171.300 95.690 171.640 ;
        RECT 84.330 170.860 85.250 171.200 ;
        RECT 88.650 170.860 89.570 171.200 ;
        RECT 82.330 169.540 83.250 169.880 ;
        RECT 90.810 169.540 91.730 169.880 ;
        RECT 78.370 168.660 79.290 169.000 ;
        RECT 82.330 168.660 83.250 169.000 ;
        RECT 90.810 168.660 91.730 169.000 ;
        RECT 94.770 168.660 95.690 169.000 ;
        RECT 78.370 166.900 79.290 167.240 ;
        RECT 82.330 166.900 83.250 167.240 ;
        RECT 90.810 166.900 91.730 167.240 ;
        RECT 94.770 166.900 95.690 167.240 ;
        RECT 79.960 165.730 80.300 166.650 ;
        RECT 93.760 165.730 94.100 166.650 ;
        RECT 78.370 165.140 79.290 165.480 ;
        RECT 82.330 165.140 83.250 165.480 ;
        RECT 90.810 165.140 91.730 165.480 ;
        RECT 94.770 165.140 95.690 165.480 ;
        RECT 78.370 164.260 79.290 164.600 ;
        RECT 82.330 164.260 83.250 164.600 ;
        RECT 90.810 164.260 91.730 164.600 ;
        RECT 94.770 164.260 95.690 164.600 ;
        RECT 78.370 162.500 79.290 162.840 ;
        RECT 82.330 162.500 83.250 162.840 ;
        RECT 90.810 162.500 91.730 162.840 ;
        RECT 94.770 162.500 95.690 162.840 ;
        RECT 80.745 161.330 81.085 162.250 ;
        RECT 83.690 161.180 85.410 161.520 ;
        RECT 88.650 161.180 90.370 161.520 ;
        RECT 92.975 161.330 93.315 162.250 ;
        RECT 78.370 160.740 79.290 161.080 ;
        RECT 82.330 160.740 83.250 161.080 ;
        RECT 78.370 159.860 79.290 160.200 ;
        RECT 82.330 159.860 83.250 160.200 ;
        RECT 78.370 158.100 79.290 158.440 ;
        RECT 82.330 158.100 83.250 158.440 ;
        RECT 77.570 157.220 79.290 157.560 ;
        RECT 81.460 156.930 81.800 157.850 ;
        RECT 78.370 156.340 79.290 156.680 ;
        RECT 82.330 156.340 83.250 156.680 ;
        RECT 78.370 155.460 79.290 155.800 ;
        RECT 82.330 155.460 83.250 155.800 ;
        RECT 78.370 153.700 79.290 154.040 ;
        RECT 82.330 153.700 83.250 154.040 ;
        RECT 78.370 151.940 79.290 152.280 ;
        RECT 82.330 151.940 83.250 152.280 ;
        RECT 76.050 150.620 76.970 150.960 ;
        RECT 78.370 148.420 79.290 148.760 ;
        RECT 82.330 148.420 83.250 148.760 ;
        RECT 83.690 147.880 84.030 161.180 ;
        RECT 84.330 156.780 85.250 157.120 ;
        RECT 88.810 156.780 89.730 157.120 ;
        RECT 84.490 150.620 86.050 150.960 ;
        RECT 84.330 148.860 85.250 149.200 ;
        RECT 82.330 147.540 84.030 147.880 ;
        RECT 85.710 147.440 86.050 150.620 ;
        RECT 84.490 147.100 86.050 147.440 ;
        RECT 83.690 145.340 85.250 145.680 ;
        RECT 78.370 144.900 79.290 145.240 ;
        RECT 82.330 144.900 83.250 145.240 ;
        RECT 78.370 143.140 79.290 143.480 ;
        RECT 82.330 143.140 83.250 143.480 ;
        RECT 78.370 142.260 79.290 142.600 ;
        RECT 82.330 141.380 83.250 141.720 ;
        RECT 82.330 140.500 83.250 140.840 ;
        RECT 83.690 140.400 84.030 145.340 ;
        RECT 83.690 140.060 85.250 140.400 ;
        RECT 75.410 137.860 79.290 138.200 ;
        RECT 82.330 137.860 83.250 138.200 ;
        RECT 69.570 136.980 70.490 137.320 ;
        RECT 78.370 136.980 79.290 137.320 ;
        RECT 85.710 136.880 86.050 147.100 ;
        RECT 62.810 136.540 64.530 136.880 ;
        RECT 84.330 136.540 86.050 136.880 ;
        RECT 88.010 150.620 89.570 150.960 ;
        RECT 88.010 147.440 88.350 150.620 ;
        RECT 88.650 148.860 89.570 149.200 ;
        RECT 90.030 147.880 90.370 161.180 ;
        RECT 90.810 160.740 91.730 161.080 ;
        RECT 94.770 160.740 95.690 161.080 ;
        RECT 90.810 159.860 91.730 160.200 ;
        RECT 94.770 159.860 95.690 160.200 ;
        RECT 90.810 158.100 91.730 158.440 ;
        RECT 94.770 158.100 95.690 158.440 ;
        RECT 92.260 156.930 92.600 157.850 ;
        RECT 96.150 157.560 96.490 171.740 ;
        RECT 94.770 157.220 96.490 157.560 ;
        RECT 90.810 156.340 91.730 156.680 ;
        RECT 94.770 156.340 95.690 156.680 ;
        RECT 90.810 155.460 91.730 155.800 ;
        RECT 94.770 155.460 95.690 155.800 ;
        RECT 90.810 153.700 91.730 154.040 ;
        RECT 94.770 153.700 95.690 154.040 ;
        RECT 90.810 151.940 91.730 152.280 ;
        RECT 94.770 151.940 95.690 152.280 ;
        RECT 96.930 150.620 97.850 150.960 ;
        RECT 90.810 148.420 91.730 148.760 ;
        RECT 94.770 148.420 95.690 148.760 ;
        RECT 90.030 147.540 91.730 147.880 ;
        RECT 88.010 147.100 89.570 147.440 ;
        RECT 88.010 136.880 88.350 147.100 ;
        RECT 88.810 145.340 90.370 145.680 ;
        RECT 90.030 140.400 90.370 145.340 ;
        RECT 90.810 144.900 91.730 145.240 ;
        RECT 94.770 144.900 95.690 145.240 ;
        RECT 90.810 143.140 91.730 143.480 ;
        RECT 94.770 143.140 95.690 143.480 ;
        RECT 94.770 142.260 95.690 142.600 ;
        RECT 90.810 141.380 91.730 141.720 ;
        RECT 90.810 140.500 91.730 140.840 ;
        RECT 88.810 140.060 90.370 140.400 ;
        RECT 98.310 138.200 98.650 174.380 ;
        RECT 90.810 137.860 91.730 138.200 ;
        RECT 94.770 137.860 98.650 138.200 ;
        RECT 100.610 174.380 102.330 174.720 ;
        RECT 100.610 138.200 100.950 174.380 ;
        RECT 103.570 173.940 104.490 174.280 ;
        RECT 107.530 173.940 108.450 174.280 ;
        RECT 108.890 173.400 109.230 178.780 ;
        RECT 122.130 177.900 123.050 178.240 ;
        RECT 116.010 177.460 116.930 177.800 ;
        RECT 119.970 177.460 120.890 177.800 ;
        RECT 115.230 176.580 116.930 176.920 ;
        RECT 119.970 176.580 120.890 176.920 ;
        RECT 115.230 173.840 115.570 176.580 ;
        RECT 116.010 174.820 116.930 175.160 ;
        RECT 119.970 174.820 120.890 175.160 ;
        RECT 107.530 173.060 109.230 173.400 ;
        RECT 113.210 173.500 115.570 173.840 ;
        RECT 109.530 172.620 110.450 172.960 ;
        RECT 101.410 171.740 103.110 172.080 ;
        RECT 102.770 157.560 103.110 171.740 ;
        RECT 103.570 171.300 104.490 171.640 ;
        RECT 107.530 171.300 108.450 171.640 ;
        RECT 109.530 170.860 110.450 171.200 ;
        RECT 107.530 169.540 108.450 169.880 ;
        RECT 103.570 168.660 104.490 169.000 ;
        RECT 107.530 168.660 108.450 169.000 ;
        RECT 103.570 166.900 104.490 167.240 ;
        RECT 107.530 166.900 108.450 167.240 ;
        RECT 113.210 166.800 113.550 173.500 ;
        RECT 116.010 173.060 116.930 173.400 ;
        RECT 119.970 173.060 120.890 173.400 ;
        RECT 126.710 170.190 127.050 213.600 ;
        RECT 135.210 207.985 135.510 222.960 ;
        RECT 136.440 203.095 136.740 223.960 ;
        RECT 146.520 208.025 146.880 208.445 ;
        RECT 140.035 206.315 140.955 206.655 ;
        RECT 143.995 206.315 144.915 206.655 ;
        RECT 140.035 205.435 140.955 205.775 ;
        RECT 143.995 205.435 144.915 205.775 ;
        RECT 144.155 204.855 145.075 204.895 ;
        RECT 146.550 204.855 146.850 208.025 ;
        RECT 143.395 204.555 148.855 204.855 ;
        RECT 146.550 204.550 146.850 204.555 ;
        RECT 140.035 203.675 140.955 204.015 ;
        RECT 143.995 203.675 144.915 204.015 ;
        RECT 140.195 203.095 141.115 203.135 ;
        RECT 136.255 202.795 141.115 203.095 ;
        RECT 136.440 202.790 136.740 202.795 ;
        RECT 140.035 201.915 140.955 202.255 ;
        RECT 143.995 201.915 144.915 202.255 ;
        RECT 140.035 201.035 140.955 201.375 ;
        RECT 143.995 201.035 144.915 201.375 ;
        RECT 132.080 200.850 132.480 200.910 ;
        RECT 138.035 200.895 138.955 200.935 ;
        RECT 136.255 200.850 138.955 200.895 ;
        RECT 132.080 200.595 138.955 200.850 ;
        RECT 132.080 200.510 136.680 200.595 ;
        RECT 132.080 200.450 132.480 200.510 ;
        RECT 114.010 167.340 115.570 167.680 ;
        RECT 105.160 165.730 105.500 166.650 ;
        RECT 113.210 166.460 114.770 166.800 ;
        RECT 103.570 165.140 104.490 165.480 ;
        RECT 107.530 165.140 108.450 165.480 ;
        RECT 103.570 164.260 104.490 164.600 ;
        RECT 107.530 164.260 108.450 164.600 ;
        RECT 103.570 162.500 104.490 162.840 ;
        RECT 107.530 162.500 108.450 162.840 ;
        RECT 105.945 161.330 106.285 162.250 ;
        RECT 108.890 161.180 110.610 161.520 ;
        RECT 103.570 160.740 104.490 161.080 ;
        RECT 107.530 160.740 108.450 161.080 ;
        RECT 103.570 159.860 104.490 160.200 ;
        RECT 107.530 159.860 108.450 160.200 ;
        RECT 103.570 158.100 104.490 158.440 ;
        RECT 107.530 158.100 108.450 158.440 ;
        RECT 102.770 157.220 104.490 157.560 ;
        RECT 106.660 156.930 107.000 157.850 ;
        RECT 103.570 156.340 104.490 156.680 ;
        RECT 107.530 156.340 108.450 156.680 ;
        RECT 103.570 155.460 104.490 155.800 ;
        RECT 107.530 155.460 108.450 155.800 ;
        RECT 103.570 153.700 104.490 154.040 ;
        RECT 107.530 153.700 108.450 154.040 ;
        RECT 103.570 151.940 104.490 152.280 ;
        RECT 107.530 151.940 108.450 152.280 ;
        RECT 101.250 150.620 102.170 150.960 ;
        RECT 103.570 148.420 104.490 148.760 ;
        RECT 107.530 148.420 108.450 148.760 ;
        RECT 108.890 147.880 109.230 161.180 ;
        RECT 109.530 156.780 110.450 157.120 ;
        RECT 109.690 150.620 111.250 150.960 ;
        RECT 109.530 148.860 110.450 149.200 ;
        RECT 107.530 147.540 109.230 147.880 ;
        RECT 110.910 147.440 111.250 150.620 ;
        RECT 109.690 147.100 111.250 147.440 ;
        RECT 108.890 145.340 110.450 145.680 ;
        RECT 103.570 144.900 104.490 145.240 ;
        RECT 107.530 144.900 108.450 145.240 ;
        RECT 103.570 143.140 104.490 143.480 ;
        RECT 107.530 143.140 108.450 143.480 ;
        RECT 103.570 142.260 104.490 142.600 ;
        RECT 107.530 141.380 108.450 141.720 ;
        RECT 107.530 140.500 108.450 140.840 ;
        RECT 108.890 140.400 109.230 145.340 ;
        RECT 108.890 140.060 110.450 140.400 ;
        RECT 100.610 137.860 104.490 138.200 ;
        RECT 107.530 137.860 108.450 138.200 ;
        RECT 94.770 136.980 95.690 137.320 ;
        RECT 103.570 136.980 104.490 137.320 ;
        RECT 110.910 136.880 111.250 147.100 ;
        RECT 88.010 136.540 89.730 136.880 ;
        RECT 109.530 136.540 111.250 136.880 ;
        RECT 113.210 136.880 113.550 166.460 ;
        RECT 115.230 164.160 115.570 167.340 ;
        RECT 119.970 166.900 120.890 167.240 ;
        RECT 116.010 166.020 116.930 166.360 ;
        RECT 119.970 165.140 120.890 165.480 ;
        RECT 113.850 163.820 115.570 164.160 ;
        RECT 119.970 163.380 120.890 163.720 ;
        RECT 119.970 162.500 121.690 162.840 ;
        RECT 119.970 161.620 120.890 161.960 ;
        RECT 119.970 159.860 120.890 160.200 ;
        RECT 116.010 158.980 116.930 159.320 ;
        RECT 116.010 158.100 116.930 158.440 ;
        RECT 119.970 158.100 120.890 158.440 ;
        RECT 116.010 156.340 116.930 156.680 ;
        RECT 119.970 156.340 120.890 156.680 ;
        RECT 119.970 155.460 120.890 155.800 ;
        RECT 116.010 154.580 116.930 154.920 ;
        RECT 119.970 154.580 120.890 154.920 ;
        RECT 116.010 153.700 116.930 154.040 ;
        RECT 119.970 153.700 120.890 154.040 ;
        RECT 116.010 151.940 116.930 152.280 ;
        RECT 119.970 151.940 120.890 152.280 ;
        RECT 116.170 151.230 117.090 151.570 ;
        RECT 121.350 150.960 121.690 162.500 ;
        RECT 122.130 161.180 123.050 161.520 ;
        RECT 121.350 150.620 123.050 150.960 ;
        RECT 116.010 150.180 116.930 150.520 ;
        RECT 119.970 150.180 120.890 150.520 ;
        RECT 119.970 149.300 120.890 149.640 ;
        RECT 121.350 148.320 121.690 150.620 ;
        RECT 121.350 147.980 123.050 148.320 ;
        RECT 119.970 147.540 120.890 147.880 ;
        RECT 119.970 145.780 120.890 146.120 ;
        RECT 122.130 145.340 123.050 145.680 ;
        RECT 114.010 144.460 115.570 144.800 ;
        RECT 115.230 141.280 115.570 144.460 ;
        RECT 119.970 144.020 120.890 144.360 ;
        RECT 116.010 143.140 116.930 143.480 ;
        RECT 113.850 140.940 115.570 141.280 ;
        RECT 119.970 136.980 120.890 137.320 ;
        RECT 113.210 136.540 114.770 136.880 ;
        RECT 116.010 136.100 116.930 136.440 ;
        RECT 15.210 135.220 16.130 135.560 ;
        RECT 19.170 135.220 20.090 135.560 ;
        RECT 27.970 135.220 28.890 135.560 ;
        RECT 31.930 135.220 32.850 135.560 ;
        RECT 40.410 135.220 41.330 135.560 ;
        RECT 44.370 135.220 45.290 135.560 ;
        RECT 53.170 135.220 54.090 135.560 ;
        RECT 57.130 135.220 58.050 135.560 ;
        RECT 65.610 135.220 66.530 135.560 ;
        RECT 69.570 135.220 70.490 135.560 ;
        RECT 78.370 135.220 79.290 135.560 ;
        RECT 82.330 135.220 83.250 135.560 ;
        RECT 90.810 135.220 91.730 135.560 ;
        RECT 94.770 135.220 95.690 135.560 ;
        RECT 103.570 135.220 104.490 135.560 ;
        RECT 107.530 135.220 108.450 135.560 ;
        RECT 116.010 135.220 116.930 135.560 ;
        RECT 119.970 135.220 120.890 135.560 ;
        RECT 15.210 134.340 16.130 134.680 ;
        RECT 19.170 134.340 20.090 134.680 ;
        RECT 27.970 134.340 28.890 134.680 ;
        RECT 31.930 134.340 32.850 134.680 ;
        RECT 40.410 134.340 41.330 134.680 ;
        RECT 44.370 134.340 45.290 134.680 ;
        RECT 53.170 134.340 54.090 134.680 ;
        RECT 57.130 134.340 58.050 134.680 ;
        RECT 65.610 134.340 66.530 134.680 ;
        RECT 69.570 134.340 70.490 134.680 ;
        RECT 78.370 134.340 79.290 134.680 ;
        RECT 82.330 134.340 83.250 134.680 ;
        RECT 90.810 134.340 91.730 134.680 ;
        RECT 94.770 134.340 95.690 134.680 ;
        RECT 103.570 134.340 104.490 134.680 ;
        RECT 107.530 134.340 108.450 134.680 ;
        RECT 116.010 134.340 116.930 134.680 ;
        RECT 119.970 134.340 120.890 134.680 ;
        RECT 12.240 106.170 55.480 106.510 ;
        RECT 7.290 89.510 8.210 90.430 ;
        RECT 12.240 89.510 12.580 106.170 ;
        RECT 12.900 89.510 13.240 106.170 ;
        RECT 13.560 94.070 13.900 106.170 ;
        RECT 13.560 92.850 13.900 93.770 ;
        RECT 13.560 89.510 13.900 92.550 ;
        RECT 14.220 89.510 14.560 106.170 ;
        RECT 14.880 94.070 15.220 106.170 ;
        RECT 14.880 92.850 15.220 93.770 ;
        RECT 14.880 89.510 15.220 92.550 ;
        RECT 15.540 89.510 15.880 106.170 ;
        RECT 16.200 94.070 16.540 106.170 ;
        RECT 16.200 92.850 16.540 93.770 ;
        RECT 16.200 89.510 16.540 92.550 ;
        RECT 16.860 89.510 17.200 106.170 ;
        RECT 17.520 94.070 17.860 106.170 ;
        RECT 17.520 92.850 17.860 93.770 ;
        RECT 17.520 89.510 17.860 92.550 ;
        RECT 18.180 89.510 18.520 106.170 ;
        RECT 18.840 100.110 19.180 106.170 ;
        RECT 18.840 98.890 19.180 99.810 ;
        RECT 18.840 89.510 19.180 98.590 ;
        RECT 19.500 89.510 19.840 106.170 ;
        RECT 20.160 100.110 20.500 106.170 ;
        RECT 20.160 98.890 20.500 99.810 ;
        RECT 20.160 89.510 20.500 98.590 ;
        RECT 20.820 89.510 21.160 106.170 ;
        RECT 21.480 103.130 21.820 106.170 ;
        RECT 21.480 101.910 21.820 102.830 ;
        RECT 21.480 89.510 21.820 101.610 ;
        RECT 22.140 89.510 22.480 106.170 ;
        RECT 22.800 104.930 23.140 105.850 ;
        RECT 22.800 89.510 23.140 104.630 ;
        RECT 23.460 89.510 23.800 106.170 ;
        RECT 24.120 97.090 24.460 106.170 ;
        RECT 24.120 95.870 24.460 96.790 ;
        RECT 24.120 89.510 24.460 95.570 ;
        RECT 24.780 89.510 25.120 106.170 ;
        RECT 25.440 103.130 25.780 106.170 ;
        RECT 25.440 101.910 25.780 102.830 ;
        RECT 25.440 89.510 25.780 101.610 ;
        RECT 26.100 89.510 26.440 106.170 ;
        RECT 26.760 100.110 27.100 106.170 ;
        RECT 26.760 98.890 27.100 99.810 ;
        RECT 26.760 89.510 27.100 98.590 ;
        RECT 27.420 89.510 27.760 106.170 ;
        RECT 28.080 100.110 28.420 106.170 ;
        RECT 28.080 98.890 28.420 99.810 ;
        RECT 28.080 89.510 28.420 98.590 ;
        RECT 28.740 89.510 29.080 106.170 ;
        RECT 29.400 94.070 29.740 106.170 ;
        RECT 29.400 92.850 29.740 93.770 ;
        RECT 29.400 89.510 29.740 92.550 ;
        RECT 30.060 89.510 30.400 106.170 ;
        RECT 30.720 94.070 31.060 106.170 ;
        RECT 30.720 92.850 31.060 93.770 ;
        RECT 30.720 89.510 31.060 92.550 ;
        RECT 31.380 89.510 31.720 106.170 ;
        RECT 32.040 94.070 32.380 106.170 ;
        RECT 32.040 92.850 32.380 93.770 ;
        RECT 32.040 89.510 32.380 92.550 ;
        RECT 32.700 89.510 33.040 106.170 ;
        RECT 33.360 94.070 33.700 106.170 ;
        RECT 33.360 92.850 33.700 93.770 ;
        RECT 33.360 89.510 33.700 92.550 ;
        RECT 34.020 89.510 34.360 106.170 ;
        RECT 34.680 94.070 35.020 106.170 ;
        RECT 34.680 92.850 35.020 93.770 ;
        RECT 34.680 89.510 35.020 92.550 ;
        RECT 35.340 89.510 35.680 106.170 ;
        RECT 36.000 94.070 36.340 106.170 ;
        RECT 36.000 92.850 36.340 93.770 ;
        RECT 36.000 89.510 36.340 92.550 ;
        RECT 36.660 89.510 37.000 106.170 ;
        RECT 37.320 94.070 37.660 106.170 ;
        RECT 37.320 92.850 37.660 93.770 ;
        RECT 37.320 89.510 37.660 92.550 ;
        RECT 37.980 89.510 38.320 106.170 ;
        RECT 38.640 94.070 38.980 106.170 ;
        RECT 38.640 92.850 38.980 93.770 ;
        RECT 38.640 89.510 38.980 92.550 ;
        RECT 39.300 89.510 39.640 106.170 ;
        RECT 39.960 100.110 40.300 106.170 ;
        RECT 39.960 98.890 40.300 99.810 ;
        RECT 39.960 89.510 40.300 98.590 ;
        RECT 40.620 89.510 40.960 106.170 ;
        RECT 41.280 100.110 41.620 106.170 ;
        RECT 41.280 98.890 41.620 99.810 ;
        RECT 41.280 89.510 41.620 98.590 ;
        RECT 41.940 89.510 42.280 106.170 ;
        RECT 42.600 103.130 42.940 106.170 ;
        RECT 42.600 101.910 42.940 102.830 ;
        RECT 42.600 89.510 42.940 101.610 ;
        RECT 43.260 89.510 43.600 106.170 ;
        RECT 43.920 97.090 44.260 106.170 ;
        RECT 43.920 95.870 44.260 96.790 ;
        RECT 43.920 89.510 44.260 95.570 ;
        RECT 44.580 89.510 44.920 106.170 ;
        RECT 45.240 91.050 45.580 106.170 ;
        RECT 45.240 89.830 45.580 90.750 ;
        RECT 45.900 89.510 46.240 106.170 ;
        RECT 46.560 103.130 46.900 106.170 ;
        RECT 46.560 101.910 46.900 102.830 ;
        RECT 46.560 89.510 46.900 101.610 ;
        RECT 47.220 89.510 47.560 106.170 ;
        RECT 47.880 100.110 48.220 106.170 ;
        RECT 47.880 98.890 48.220 99.810 ;
        RECT 47.880 89.510 48.220 98.590 ;
        RECT 48.540 89.510 48.880 106.170 ;
        RECT 49.200 100.110 49.540 106.170 ;
        RECT 49.200 98.890 49.540 99.810 ;
        RECT 49.200 89.510 49.540 98.590 ;
        RECT 49.860 89.510 50.200 106.170 ;
        RECT 50.520 94.070 50.860 106.170 ;
        RECT 50.520 92.850 50.860 93.770 ;
        RECT 50.520 89.510 50.860 92.550 ;
        RECT 51.180 89.510 51.520 106.170 ;
        RECT 51.840 94.070 52.180 106.170 ;
        RECT 51.840 92.850 52.180 93.770 ;
        RECT 51.840 89.510 52.180 92.550 ;
        RECT 52.500 89.510 52.840 106.170 ;
        RECT 53.160 94.070 53.500 106.170 ;
        RECT 53.160 92.850 53.500 93.770 ;
        RECT 53.160 89.510 53.500 92.550 ;
        RECT 53.820 89.510 54.160 106.170 ;
        RECT 54.480 94.070 54.820 106.170 ;
        RECT 54.480 92.850 54.820 93.770 ;
        RECT 54.480 89.510 54.820 92.550 ;
        RECT 55.140 89.510 55.480 106.170 ;
        RECT 56.120 105.220 57.040 105.560 ;
        RECT 56.120 102.200 57.040 102.540 ;
        RECT 56.120 99.180 57.040 99.520 ;
        RECT 56.120 96.160 57.040 96.500 ;
        RECT 56.120 93.140 57.040 93.480 ;
        RECT 56.120 90.120 57.040 90.460 ;
        RECT 57.900 89.830 58.240 116.100 ;
        RECT 7.290 89.170 55.480 89.510 ;
        RECT 7.290 72.510 8.210 73.430 ;
        RECT 12.240 72.510 12.580 89.170 ;
        RECT 12.900 72.510 13.240 89.170 ;
        RECT 13.560 77.070 13.900 89.170 ;
        RECT 13.560 75.850 13.900 76.770 ;
        RECT 13.560 72.510 13.900 75.550 ;
        RECT 14.220 72.510 14.560 89.170 ;
        RECT 14.880 77.070 15.220 89.170 ;
        RECT 14.880 75.850 15.220 76.770 ;
        RECT 14.880 72.510 15.220 75.550 ;
        RECT 15.540 72.510 15.880 89.170 ;
        RECT 16.200 77.070 16.540 89.170 ;
        RECT 16.200 75.850 16.540 76.770 ;
        RECT 16.200 72.510 16.540 75.550 ;
        RECT 16.860 72.510 17.200 89.170 ;
        RECT 17.520 77.070 17.860 89.170 ;
        RECT 17.520 75.850 17.860 76.770 ;
        RECT 17.520 72.510 17.860 75.550 ;
        RECT 18.180 72.510 18.520 89.170 ;
        RECT 18.840 83.110 19.180 89.170 ;
        RECT 18.840 81.890 19.180 82.810 ;
        RECT 18.840 72.510 19.180 81.590 ;
        RECT 19.500 72.510 19.840 89.170 ;
        RECT 20.160 83.110 20.500 89.170 ;
        RECT 20.160 81.890 20.500 82.810 ;
        RECT 20.160 72.510 20.500 81.590 ;
        RECT 20.820 72.510 21.160 89.170 ;
        RECT 21.480 86.130 21.820 89.170 ;
        RECT 21.480 84.910 21.820 85.830 ;
        RECT 21.480 72.510 21.820 84.610 ;
        RECT 22.140 72.510 22.480 89.170 ;
        RECT 22.800 87.930 23.140 88.850 ;
        RECT 22.800 72.510 23.140 87.630 ;
        RECT 23.460 72.510 23.800 89.170 ;
        RECT 24.120 80.090 24.460 89.170 ;
        RECT 24.120 78.870 24.460 79.790 ;
        RECT 24.120 72.510 24.460 78.570 ;
        RECT 24.780 72.510 25.120 89.170 ;
        RECT 25.440 86.130 25.780 89.170 ;
        RECT 25.440 84.910 25.780 85.830 ;
        RECT 25.440 72.510 25.780 84.610 ;
        RECT 26.100 72.510 26.440 89.170 ;
        RECT 26.760 83.110 27.100 89.170 ;
        RECT 26.760 81.890 27.100 82.810 ;
        RECT 26.760 72.510 27.100 81.590 ;
        RECT 27.420 72.510 27.760 89.170 ;
        RECT 28.080 83.110 28.420 89.170 ;
        RECT 28.080 81.890 28.420 82.810 ;
        RECT 28.080 72.510 28.420 81.590 ;
        RECT 28.740 72.510 29.080 89.170 ;
        RECT 29.400 77.070 29.740 89.170 ;
        RECT 29.400 75.850 29.740 76.770 ;
        RECT 29.400 72.510 29.740 75.550 ;
        RECT 30.060 72.510 30.400 89.170 ;
        RECT 30.720 77.070 31.060 89.170 ;
        RECT 30.720 75.850 31.060 76.770 ;
        RECT 30.720 72.510 31.060 75.550 ;
        RECT 31.380 72.510 31.720 89.170 ;
        RECT 32.040 77.070 32.380 89.170 ;
        RECT 32.040 75.850 32.380 76.770 ;
        RECT 32.040 72.510 32.380 75.550 ;
        RECT 32.700 72.510 33.040 89.170 ;
        RECT 33.360 77.070 33.700 89.170 ;
        RECT 33.360 75.850 33.700 76.770 ;
        RECT 33.360 72.510 33.700 75.550 ;
        RECT 34.020 72.510 34.360 89.170 ;
        RECT 34.680 77.070 35.020 89.170 ;
        RECT 34.680 75.850 35.020 76.770 ;
        RECT 34.680 72.510 35.020 75.550 ;
        RECT 35.340 72.510 35.680 89.170 ;
        RECT 36.000 77.070 36.340 89.170 ;
        RECT 36.000 75.850 36.340 76.770 ;
        RECT 36.000 72.510 36.340 75.550 ;
        RECT 36.660 72.510 37.000 89.170 ;
        RECT 37.320 77.070 37.660 89.170 ;
        RECT 37.320 75.850 37.660 76.770 ;
        RECT 37.320 72.510 37.660 75.550 ;
        RECT 37.980 72.510 38.320 89.170 ;
        RECT 38.640 77.070 38.980 89.170 ;
        RECT 38.640 75.850 38.980 76.770 ;
        RECT 38.640 72.510 38.980 75.550 ;
        RECT 39.300 72.510 39.640 89.170 ;
        RECT 39.960 83.110 40.300 89.170 ;
        RECT 39.960 81.890 40.300 82.810 ;
        RECT 39.960 72.510 40.300 81.590 ;
        RECT 40.620 72.510 40.960 89.170 ;
        RECT 41.280 83.110 41.620 89.170 ;
        RECT 41.280 81.890 41.620 82.810 ;
        RECT 41.280 72.510 41.620 81.590 ;
        RECT 41.940 72.510 42.280 89.170 ;
        RECT 42.600 86.130 42.940 89.170 ;
        RECT 42.600 84.910 42.940 85.830 ;
        RECT 42.600 72.510 42.940 84.610 ;
        RECT 43.260 72.510 43.600 89.170 ;
        RECT 43.920 80.090 44.260 89.170 ;
        RECT 43.920 78.870 44.260 79.790 ;
        RECT 43.920 72.510 44.260 78.570 ;
        RECT 44.580 72.510 44.920 89.170 ;
        RECT 45.240 74.050 45.580 89.170 ;
        RECT 45.240 72.830 45.580 73.750 ;
        RECT 45.900 72.510 46.240 89.170 ;
        RECT 46.560 86.130 46.900 89.170 ;
        RECT 46.560 84.910 46.900 85.830 ;
        RECT 46.560 72.510 46.900 84.610 ;
        RECT 47.220 72.510 47.560 89.170 ;
        RECT 47.880 83.110 48.220 89.170 ;
        RECT 47.880 81.890 48.220 82.810 ;
        RECT 47.880 72.510 48.220 81.590 ;
        RECT 48.540 72.510 48.880 89.170 ;
        RECT 49.200 83.110 49.540 89.170 ;
        RECT 49.200 81.890 49.540 82.810 ;
        RECT 49.200 72.510 49.540 81.590 ;
        RECT 49.860 72.510 50.200 89.170 ;
        RECT 50.520 77.070 50.860 89.170 ;
        RECT 50.520 75.850 50.860 76.770 ;
        RECT 50.520 72.510 50.860 75.550 ;
        RECT 51.180 72.510 51.520 89.170 ;
        RECT 51.840 77.070 52.180 89.170 ;
        RECT 51.840 75.850 52.180 76.770 ;
        RECT 51.840 72.510 52.180 75.550 ;
        RECT 52.500 72.510 52.840 89.170 ;
        RECT 53.160 77.070 53.500 89.170 ;
        RECT 53.160 75.850 53.500 76.770 ;
        RECT 53.160 72.510 53.500 75.550 ;
        RECT 53.820 72.510 54.160 89.170 ;
        RECT 54.480 77.070 54.820 89.170 ;
        RECT 54.480 75.850 54.820 76.770 ;
        RECT 54.480 72.510 54.820 75.550 ;
        RECT 55.140 72.510 55.480 89.170 ;
        RECT 56.120 88.220 57.040 88.560 ;
        RECT 56.120 85.200 57.040 85.540 ;
        RECT 56.120 82.180 57.040 82.520 ;
        RECT 56.120 79.160 57.040 79.500 ;
        RECT 56.120 76.140 57.040 76.480 ;
        RECT 56.120 73.120 57.040 73.460 ;
        RECT 7.290 72.170 55.480 72.510 ;
        RECT 7.290 55.510 8.210 56.430 ;
        RECT 12.240 55.510 12.580 72.170 ;
        RECT 12.900 55.510 13.240 72.170 ;
        RECT 13.560 60.070 13.900 72.170 ;
        RECT 13.560 58.850 13.900 59.770 ;
        RECT 13.560 55.510 13.900 58.550 ;
        RECT 14.220 55.510 14.560 72.170 ;
        RECT 14.880 60.070 15.220 72.170 ;
        RECT 14.880 58.850 15.220 59.770 ;
        RECT 14.880 55.510 15.220 58.550 ;
        RECT 15.540 55.510 15.880 72.170 ;
        RECT 16.200 60.070 16.540 72.170 ;
        RECT 16.200 58.850 16.540 59.770 ;
        RECT 16.200 55.510 16.540 58.550 ;
        RECT 16.860 55.510 17.200 72.170 ;
        RECT 17.520 60.070 17.860 72.170 ;
        RECT 17.520 58.850 17.860 59.770 ;
        RECT 17.520 55.510 17.860 58.550 ;
        RECT 18.180 55.510 18.520 72.170 ;
        RECT 18.840 66.110 19.180 72.170 ;
        RECT 18.840 64.890 19.180 65.810 ;
        RECT 18.840 55.510 19.180 64.590 ;
        RECT 19.500 55.510 19.840 72.170 ;
        RECT 20.160 66.110 20.500 72.170 ;
        RECT 20.160 64.890 20.500 65.810 ;
        RECT 20.160 55.510 20.500 64.590 ;
        RECT 20.820 55.510 21.160 72.170 ;
        RECT 21.480 69.130 21.820 72.170 ;
        RECT 21.480 67.910 21.820 68.830 ;
        RECT 21.480 55.510 21.820 67.610 ;
        RECT 22.140 55.510 22.480 72.170 ;
        RECT 22.800 70.930 23.140 71.850 ;
        RECT 22.800 55.510 23.140 70.630 ;
        RECT 23.460 55.510 23.800 72.170 ;
        RECT 24.120 63.090 24.460 72.170 ;
        RECT 24.120 61.870 24.460 62.790 ;
        RECT 24.120 55.510 24.460 61.570 ;
        RECT 24.780 55.510 25.120 72.170 ;
        RECT 25.440 69.130 25.780 72.170 ;
        RECT 25.440 67.910 25.780 68.830 ;
        RECT 25.440 55.510 25.780 67.610 ;
        RECT 26.100 55.510 26.440 72.170 ;
        RECT 26.760 66.110 27.100 72.170 ;
        RECT 26.760 64.890 27.100 65.810 ;
        RECT 26.760 55.510 27.100 64.590 ;
        RECT 27.420 55.510 27.760 72.170 ;
        RECT 28.080 66.110 28.420 72.170 ;
        RECT 28.080 64.890 28.420 65.810 ;
        RECT 28.080 55.510 28.420 64.590 ;
        RECT 28.740 55.510 29.080 72.170 ;
        RECT 29.400 60.070 29.740 72.170 ;
        RECT 29.400 58.850 29.740 59.770 ;
        RECT 29.400 55.510 29.740 58.550 ;
        RECT 30.060 55.510 30.400 72.170 ;
        RECT 30.720 60.070 31.060 72.170 ;
        RECT 30.720 58.850 31.060 59.770 ;
        RECT 30.720 55.510 31.060 58.550 ;
        RECT 31.380 55.510 31.720 72.170 ;
        RECT 32.040 60.070 32.380 72.170 ;
        RECT 32.040 58.850 32.380 59.770 ;
        RECT 32.040 55.510 32.380 58.550 ;
        RECT 32.700 55.510 33.040 72.170 ;
        RECT 33.360 60.070 33.700 72.170 ;
        RECT 33.360 58.850 33.700 59.770 ;
        RECT 33.360 55.510 33.700 58.550 ;
        RECT 34.020 55.510 34.360 72.170 ;
        RECT 34.680 60.070 35.020 72.170 ;
        RECT 34.680 58.850 35.020 59.770 ;
        RECT 34.680 55.510 35.020 58.550 ;
        RECT 35.340 55.510 35.680 72.170 ;
        RECT 36.000 60.070 36.340 72.170 ;
        RECT 36.000 58.850 36.340 59.770 ;
        RECT 36.000 55.510 36.340 58.550 ;
        RECT 36.660 55.510 37.000 72.170 ;
        RECT 37.320 60.070 37.660 72.170 ;
        RECT 37.320 58.850 37.660 59.770 ;
        RECT 37.320 55.510 37.660 58.550 ;
        RECT 37.980 55.510 38.320 72.170 ;
        RECT 38.640 60.070 38.980 72.170 ;
        RECT 38.640 58.850 38.980 59.770 ;
        RECT 38.640 55.510 38.980 58.550 ;
        RECT 39.300 55.510 39.640 72.170 ;
        RECT 39.960 66.110 40.300 72.170 ;
        RECT 39.960 64.890 40.300 65.810 ;
        RECT 39.960 55.510 40.300 64.590 ;
        RECT 40.620 55.510 40.960 72.170 ;
        RECT 41.280 66.110 41.620 72.170 ;
        RECT 41.280 64.890 41.620 65.810 ;
        RECT 41.280 55.510 41.620 64.590 ;
        RECT 41.940 55.510 42.280 72.170 ;
        RECT 42.600 69.130 42.940 72.170 ;
        RECT 42.600 67.910 42.940 68.830 ;
        RECT 42.600 55.510 42.940 67.610 ;
        RECT 43.260 55.510 43.600 72.170 ;
        RECT 43.920 63.090 44.260 72.170 ;
        RECT 43.920 61.870 44.260 62.790 ;
        RECT 43.920 55.510 44.260 61.570 ;
        RECT 44.580 55.510 44.920 72.170 ;
        RECT 45.240 57.050 45.580 72.170 ;
        RECT 45.240 55.830 45.580 56.750 ;
        RECT 45.900 55.510 46.240 72.170 ;
        RECT 46.560 69.130 46.900 72.170 ;
        RECT 46.560 67.910 46.900 68.830 ;
        RECT 46.560 55.510 46.900 67.610 ;
        RECT 47.220 55.510 47.560 72.170 ;
        RECT 47.880 66.110 48.220 72.170 ;
        RECT 47.880 64.890 48.220 65.810 ;
        RECT 47.880 55.510 48.220 64.590 ;
        RECT 48.540 55.510 48.880 72.170 ;
        RECT 49.200 66.110 49.540 72.170 ;
        RECT 49.200 64.890 49.540 65.810 ;
        RECT 49.200 55.510 49.540 64.590 ;
        RECT 49.860 55.510 50.200 72.170 ;
        RECT 50.520 60.070 50.860 72.170 ;
        RECT 50.520 58.850 50.860 59.770 ;
        RECT 50.520 55.510 50.860 58.550 ;
        RECT 51.180 55.510 51.520 72.170 ;
        RECT 51.840 60.070 52.180 72.170 ;
        RECT 51.840 58.850 52.180 59.770 ;
        RECT 51.840 55.510 52.180 58.550 ;
        RECT 52.500 55.510 52.840 72.170 ;
        RECT 53.160 60.070 53.500 72.170 ;
        RECT 53.160 58.850 53.500 59.770 ;
        RECT 53.160 55.510 53.500 58.550 ;
        RECT 53.820 55.510 54.160 72.170 ;
        RECT 54.480 60.070 54.820 72.170 ;
        RECT 54.480 58.850 54.820 59.770 ;
        RECT 54.480 55.510 54.820 58.550 ;
        RECT 55.140 56.460 55.480 72.170 ;
        RECT 56.120 71.220 57.040 71.560 ;
        RECT 56.120 68.200 57.040 68.540 ;
        RECT 56.120 65.180 57.040 65.520 ;
        RECT 56.120 62.160 57.040 62.500 ;
        RECT 56.120 59.140 57.040 59.480 ;
        RECT 56.700 56.460 57.040 56.750 ;
        RECT 55.140 56.120 57.040 56.460 ;
        RECT 55.140 55.510 55.480 56.120 ;
        RECT 56.700 55.830 57.040 56.120 ;
        RECT 7.290 55.170 55.480 55.510 ;
        RECT 7.290 38.510 8.210 39.430 ;
        RECT 12.240 38.510 12.580 55.170 ;
        RECT 12.900 38.510 13.240 55.170 ;
        RECT 13.560 43.070 13.900 55.170 ;
        RECT 13.560 41.850 13.900 42.770 ;
        RECT 13.560 38.510 13.900 41.550 ;
        RECT 14.220 38.510 14.560 55.170 ;
        RECT 14.880 43.070 15.220 55.170 ;
        RECT 14.880 41.850 15.220 42.770 ;
        RECT 14.880 38.510 15.220 41.550 ;
        RECT 15.540 38.510 15.880 55.170 ;
        RECT 16.200 43.070 16.540 55.170 ;
        RECT 16.200 41.850 16.540 42.770 ;
        RECT 16.200 38.510 16.540 41.550 ;
        RECT 16.860 38.510 17.200 55.170 ;
        RECT 17.520 43.070 17.860 55.170 ;
        RECT 17.520 41.850 17.860 42.770 ;
        RECT 17.520 38.510 17.860 41.550 ;
        RECT 18.180 38.510 18.520 55.170 ;
        RECT 18.840 49.110 19.180 55.170 ;
        RECT 18.840 47.890 19.180 48.810 ;
        RECT 18.840 38.510 19.180 47.590 ;
        RECT 19.500 38.510 19.840 55.170 ;
        RECT 20.160 49.110 20.500 55.170 ;
        RECT 20.160 47.890 20.500 48.810 ;
        RECT 20.160 38.510 20.500 47.590 ;
        RECT 20.820 38.510 21.160 55.170 ;
        RECT 21.480 52.130 21.820 55.170 ;
        RECT 21.480 50.910 21.820 51.830 ;
        RECT 21.480 38.510 21.820 50.610 ;
        RECT 22.140 38.510 22.480 55.170 ;
        RECT 22.800 53.930 23.140 54.850 ;
        RECT 22.800 38.510 23.140 53.630 ;
        RECT 23.460 38.510 23.800 55.170 ;
        RECT 24.120 46.090 24.460 55.170 ;
        RECT 24.120 44.870 24.460 45.790 ;
        RECT 24.120 38.510 24.460 44.570 ;
        RECT 24.780 38.510 25.120 55.170 ;
        RECT 25.440 52.130 25.780 55.170 ;
        RECT 25.440 50.910 25.780 51.830 ;
        RECT 25.440 38.510 25.780 50.610 ;
        RECT 26.100 38.510 26.440 55.170 ;
        RECT 26.760 49.110 27.100 55.170 ;
        RECT 26.760 47.890 27.100 48.810 ;
        RECT 26.760 38.510 27.100 47.590 ;
        RECT 27.420 38.510 27.760 55.170 ;
        RECT 28.080 49.110 28.420 55.170 ;
        RECT 28.080 47.890 28.420 48.810 ;
        RECT 28.080 38.510 28.420 47.590 ;
        RECT 28.740 38.510 29.080 55.170 ;
        RECT 29.400 43.070 29.740 55.170 ;
        RECT 29.400 41.850 29.740 42.770 ;
        RECT 29.400 38.510 29.740 41.550 ;
        RECT 30.060 38.510 30.400 55.170 ;
        RECT 30.720 43.070 31.060 55.170 ;
        RECT 30.720 41.850 31.060 42.770 ;
        RECT 30.720 38.510 31.060 41.550 ;
        RECT 31.380 38.510 31.720 55.170 ;
        RECT 32.040 43.070 32.380 55.170 ;
        RECT 32.040 41.850 32.380 42.770 ;
        RECT 32.040 38.510 32.380 41.550 ;
        RECT 32.700 38.510 33.040 55.170 ;
        RECT 33.360 43.070 33.700 55.170 ;
        RECT 33.360 41.850 33.700 42.770 ;
        RECT 33.360 38.510 33.700 41.550 ;
        RECT 34.020 38.510 34.360 55.170 ;
        RECT 34.680 43.070 35.020 55.170 ;
        RECT 34.680 41.850 35.020 42.770 ;
        RECT 34.680 38.510 35.020 41.550 ;
        RECT 35.340 38.510 35.680 55.170 ;
        RECT 36.000 43.070 36.340 55.170 ;
        RECT 36.000 41.850 36.340 42.770 ;
        RECT 36.000 38.510 36.340 41.550 ;
        RECT 36.660 38.510 37.000 55.170 ;
        RECT 37.320 43.070 37.660 55.170 ;
        RECT 37.320 41.850 37.660 42.770 ;
        RECT 37.320 38.510 37.660 41.550 ;
        RECT 37.980 38.510 38.320 55.170 ;
        RECT 38.640 43.070 38.980 55.170 ;
        RECT 38.640 41.850 38.980 42.770 ;
        RECT 38.640 38.510 38.980 41.550 ;
        RECT 39.300 38.510 39.640 55.170 ;
        RECT 39.960 49.110 40.300 55.170 ;
        RECT 39.960 47.890 40.300 48.810 ;
        RECT 39.960 38.510 40.300 47.590 ;
        RECT 40.620 38.510 40.960 55.170 ;
        RECT 41.280 49.110 41.620 55.170 ;
        RECT 41.280 47.890 41.620 48.810 ;
        RECT 41.280 38.510 41.620 47.590 ;
        RECT 41.940 38.510 42.280 55.170 ;
        RECT 42.600 52.130 42.940 55.170 ;
        RECT 42.600 50.910 42.940 51.830 ;
        RECT 42.600 38.510 42.940 50.610 ;
        RECT 43.260 38.510 43.600 55.170 ;
        RECT 43.920 46.090 44.260 55.170 ;
        RECT 43.920 44.870 44.260 45.790 ;
        RECT 43.920 38.510 44.260 44.570 ;
        RECT 44.580 38.510 44.920 55.170 ;
        RECT 45.240 40.050 45.580 55.170 ;
        RECT 45.240 38.830 45.580 39.750 ;
        RECT 45.900 38.510 46.240 55.170 ;
        RECT 46.560 52.130 46.900 55.170 ;
        RECT 46.560 50.910 46.900 51.830 ;
        RECT 46.560 38.510 46.900 50.610 ;
        RECT 47.220 38.510 47.560 55.170 ;
        RECT 47.880 49.110 48.220 55.170 ;
        RECT 47.880 47.890 48.220 48.810 ;
        RECT 47.880 38.510 48.220 47.590 ;
        RECT 48.540 38.510 48.880 55.170 ;
        RECT 49.200 49.110 49.540 55.170 ;
        RECT 49.200 47.890 49.540 48.810 ;
        RECT 49.200 38.510 49.540 47.590 ;
        RECT 49.860 38.510 50.200 55.170 ;
        RECT 50.520 43.070 50.860 55.170 ;
        RECT 50.520 41.850 50.860 42.770 ;
        RECT 50.520 38.510 50.860 41.550 ;
        RECT 51.180 38.510 51.520 55.170 ;
        RECT 51.840 43.070 52.180 55.170 ;
        RECT 51.840 41.850 52.180 42.770 ;
        RECT 51.840 38.510 52.180 41.550 ;
        RECT 52.500 38.510 52.840 55.170 ;
        RECT 53.160 43.070 53.500 55.170 ;
        RECT 53.160 41.850 53.500 42.770 ;
        RECT 53.160 38.510 53.500 41.550 ;
        RECT 53.820 38.510 54.160 55.170 ;
        RECT 54.480 43.070 54.820 55.170 ;
        RECT 54.480 41.850 54.820 42.770 ;
        RECT 54.480 38.510 54.820 41.550 ;
        RECT 55.140 38.510 55.480 55.170 ;
        RECT 56.120 54.220 57.040 54.560 ;
        RECT 56.120 51.200 57.040 51.540 ;
        RECT 56.120 48.180 57.040 48.520 ;
        RECT 56.120 45.160 57.040 45.500 ;
        RECT 56.120 42.140 57.040 42.480 ;
        RECT 56.120 39.120 57.040 39.460 ;
        RECT 58.840 38.830 59.180 122.610 ;
        RECT 59.780 58.850 60.120 117.030 ;
        RECT 60.720 75.850 61.060 123.540 ;
        RECT 61.660 72.830 62.000 117.960 ;
        RECT 62.600 81.890 62.940 124.470 ;
        RECT 63.540 64.890 63.880 118.890 ;
        RECT 64.480 67.910 64.820 119.820 ;
        RECT 65.420 61.870 65.760 120.750 ;
        RECT 66.360 70.930 66.700 121.680 ;
        RECT 69.560 70.930 69.900 130.980 ;
        RECT 70.500 61.870 70.840 130.050 ;
        RECT 71.440 67.910 71.780 129.120 ;
        RECT 72.380 64.890 72.720 128.190 ;
        RECT 73.320 81.890 73.660 127.260 ;
        RECT 74.260 72.830 74.600 115.170 ;
        RECT 75.200 75.850 75.540 126.330 ;
        RECT 76.140 58.850 76.480 114.240 ;
        RECT 77.080 38.830 77.420 125.400 ;
        RECT 78.020 89.830 78.360 113.310 ;
        RECT 80.780 106.170 124.020 106.510 ;
        RECT 79.220 105.220 80.140 105.560 ;
        RECT 79.220 102.200 80.140 102.540 ;
        RECT 79.220 99.180 80.140 99.520 ;
        RECT 79.220 96.160 80.140 96.500 ;
        RECT 79.220 93.140 80.140 93.480 ;
        RECT 79.220 90.120 80.140 90.460 ;
        RECT 80.780 89.510 81.120 106.170 ;
        RECT 81.440 94.070 81.780 106.170 ;
        RECT 81.440 92.850 81.780 93.770 ;
        RECT 81.440 89.510 81.780 92.550 ;
        RECT 82.100 89.510 82.440 106.170 ;
        RECT 82.760 94.070 83.100 106.170 ;
        RECT 82.760 92.850 83.100 93.770 ;
        RECT 82.760 89.510 83.100 92.550 ;
        RECT 83.420 89.510 83.760 106.170 ;
        RECT 84.080 94.070 84.420 106.170 ;
        RECT 84.080 92.850 84.420 93.770 ;
        RECT 84.080 89.510 84.420 92.550 ;
        RECT 84.740 89.510 85.080 106.170 ;
        RECT 85.400 94.070 85.740 106.170 ;
        RECT 85.400 92.850 85.740 93.770 ;
        RECT 85.400 89.510 85.740 92.550 ;
        RECT 86.060 89.510 86.400 106.170 ;
        RECT 86.720 100.110 87.060 106.170 ;
        RECT 86.720 98.890 87.060 99.810 ;
        RECT 86.720 89.510 87.060 98.590 ;
        RECT 87.380 89.510 87.720 106.170 ;
        RECT 88.040 100.110 88.380 106.170 ;
        RECT 88.040 98.890 88.380 99.810 ;
        RECT 88.040 89.510 88.380 98.590 ;
        RECT 88.700 89.510 89.040 106.170 ;
        RECT 89.360 103.130 89.700 106.170 ;
        RECT 89.360 101.910 89.700 102.830 ;
        RECT 89.360 89.510 89.700 101.610 ;
        RECT 90.020 89.510 90.360 106.170 ;
        RECT 90.680 91.050 91.020 106.170 ;
        RECT 90.680 89.830 91.020 90.750 ;
        RECT 91.340 89.510 91.680 106.170 ;
        RECT 92.000 97.090 92.340 106.170 ;
        RECT 92.000 95.870 92.340 96.790 ;
        RECT 92.000 89.510 92.340 95.570 ;
        RECT 92.660 89.510 93.000 106.170 ;
        RECT 93.320 103.130 93.660 106.170 ;
        RECT 93.320 101.910 93.660 102.830 ;
        RECT 93.320 89.510 93.660 101.610 ;
        RECT 93.980 89.510 94.320 106.170 ;
        RECT 94.640 100.110 94.980 106.170 ;
        RECT 94.640 98.890 94.980 99.810 ;
        RECT 94.640 89.510 94.980 98.590 ;
        RECT 95.300 89.510 95.640 106.170 ;
        RECT 95.960 100.110 96.300 106.170 ;
        RECT 95.960 98.890 96.300 99.810 ;
        RECT 95.960 89.510 96.300 98.590 ;
        RECT 96.620 89.510 96.960 106.170 ;
        RECT 97.280 94.070 97.620 106.170 ;
        RECT 97.280 92.850 97.620 93.770 ;
        RECT 97.280 89.510 97.620 92.550 ;
        RECT 97.940 89.510 98.280 106.170 ;
        RECT 98.600 94.070 98.940 106.170 ;
        RECT 98.600 92.850 98.940 93.770 ;
        RECT 98.600 89.510 98.940 92.550 ;
        RECT 99.260 89.510 99.600 106.170 ;
        RECT 99.920 94.070 100.260 106.170 ;
        RECT 99.920 92.850 100.260 93.770 ;
        RECT 99.920 89.510 100.260 92.550 ;
        RECT 100.580 89.510 100.920 106.170 ;
        RECT 101.240 94.070 101.580 106.170 ;
        RECT 101.240 92.850 101.580 93.770 ;
        RECT 101.240 89.510 101.580 92.550 ;
        RECT 101.900 89.510 102.240 106.170 ;
        RECT 102.560 94.070 102.900 106.170 ;
        RECT 102.560 92.850 102.900 93.770 ;
        RECT 102.560 89.510 102.900 92.550 ;
        RECT 103.220 89.510 103.560 106.170 ;
        RECT 103.880 94.070 104.220 106.170 ;
        RECT 103.880 92.850 104.220 93.770 ;
        RECT 103.880 89.510 104.220 92.550 ;
        RECT 104.540 89.510 104.880 106.170 ;
        RECT 105.200 94.070 105.540 106.170 ;
        RECT 105.200 92.850 105.540 93.770 ;
        RECT 105.200 89.510 105.540 92.550 ;
        RECT 105.860 89.510 106.200 106.170 ;
        RECT 106.520 94.070 106.860 106.170 ;
        RECT 106.520 92.850 106.860 93.770 ;
        RECT 106.520 89.510 106.860 92.550 ;
        RECT 107.180 89.510 107.520 106.170 ;
        RECT 107.840 100.110 108.180 106.170 ;
        RECT 107.840 98.890 108.180 99.810 ;
        RECT 107.840 89.510 108.180 98.590 ;
        RECT 108.500 89.510 108.840 106.170 ;
        RECT 109.160 100.110 109.500 106.170 ;
        RECT 109.160 98.890 109.500 99.810 ;
        RECT 109.160 89.510 109.500 98.590 ;
        RECT 109.820 89.510 110.160 106.170 ;
        RECT 110.480 103.130 110.820 106.170 ;
        RECT 110.480 101.910 110.820 102.830 ;
        RECT 110.480 89.510 110.820 101.610 ;
        RECT 111.140 89.510 111.480 106.170 ;
        RECT 111.800 97.090 112.140 106.170 ;
        RECT 111.800 95.870 112.140 96.790 ;
        RECT 111.800 89.510 112.140 95.570 ;
        RECT 112.460 89.510 112.800 106.170 ;
        RECT 113.120 104.930 113.460 105.850 ;
        RECT 113.120 89.510 113.460 104.630 ;
        RECT 113.780 89.510 114.120 106.170 ;
        RECT 114.440 103.130 114.780 106.170 ;
        RECT 114.440 101.910 114.780 102.830 ;
        RECT 114.440 89.510 114.780 101.610 ;
        RECT 115.100 89.510 115.440 106.170 ;
        RECT 115.760 100.110 116.100 106.170 ;
        RECT 115.760 98.890 116.100 99.810 ;
        RECT 115.760 89.510 116.100 98.590 ;
        RECT 116.420 89.510 116.760 106.170 ;
        RECT 117.080 100.110 117.420 106.170 ;
        RECT 117.080 98.890 117.420 99.810 ;
        RECT 117.080 89.510 117.420 98.590 ;
        RECT 117.740 89.510 118.080 106.170 ;
        RECT 118.400 94.070 118.740 106.170 ;
        RECT 118.400 92.850 118.740 93.770 ;
        RECT 118.400 89.510 118.740 92.550 ;
        RECT 119.060 89.510 119.400 106.170 ;
        RECT 119.720 94.070 120.060 106.170 ;
        RECT 119.720 92.850 120.060 93.770 ;
        RECT 119.720 89.510 120.060 92.550 ;
        RECT 120.380 89.510 120.720 106.170 ;
        RECT 121.040 94.070 121.380 106.170 ;
        RECT 121.040 92.850 121.380 93.770 ;
        RECT 121.040 89.510 121.380 92.550 ;
        RECT 121.700 89.510 122.040 106.170 ;
        RECT 122.360 94.070 122.700 106.170 ;
        RECT 122.360 92.850 122.700 93.770 ;
        RECT 122.360 89.510 122.700 92.550 ;
        RECT 123.020 89.510 123.360 106.170 ;
        RECT 123.680 89.510 124.020 106.170 ;
        RECT 128.630 89.510 128.970 90.090 ;
        RECT 80.780 89.170 128.970 89.510 ;
        RECT 79.220 88.220 80.140 88.560 ;
        RECT 79.220 85.200 80.140 85.540 ;
        RECT 79.220 82.180 80.140 82.520 ;
        RECT 79.220 79.160 80.140 79.500 ;
        RECT 79.220 76.140 80.140 76.480 ;
        RECT 79.220 73.120 80.140 73.460 ;
        RECT 80.780 72.510 81.120 89.170 ;
        RECT 81.440 77.070 81.780 89.170 ;
        RECT 81.440 75.850 81.780 76.770 ;
        RECT 81.440 72.510 81.780 75.550 ;
        RECT 82.100 72.510 82.440 89.170 ;
        RECT 82.760 77.070 83.100 89.170 ;
        RECT 82.760 75.850 83.100 76.770 ;
        RECT 82.760 72.510 83.100 75.550 ;
        RECT 83.420 72.510 83.760 89.170 ;
        RECT 84.080 77.070 84.420 89.170 ;
        RECT 84.080 75.850 84.420 76.770 ;
        RECT 84.080 72.510 84.420 75.550 ;
        RECT 84.740 72.510 85.080 89.170 ;
        RECT 85.400 77.070 85.740 89.170 ;
        RECT 85.400 75.850 85.740 76.770 ;
        RECT 85.400 72.510 85.740 75.550 ;
        RECT 86.060 72.510 86.400 89.170 ;
        RECT 86.720 83.110 87.060 89.170 ;
        RECT 86.720 81.890 87.060 82.810 ;
        RECT 86.720 72.510 87.060 81.590 ;
        RECT 87.380 72.510 87.720 89.170 ;
        RECT 88.040 83.110 88.380 89.170 ;
        RECT 88.040 81.890 88.380 82.810 ;
        RECT 88.040 72.510 88.380 81.590 ;
        RECT 88.700 72.510 89.040 89.170 ;
        RECT 89.360 86.130 89.700 89.170 ;
        RECT 89.360 84.910 89.700 85.830 ;
        RECT 89.360 72.510 89.700 84.610 ;
        RECT 90.020 72.510 90.360 89.170 ;
        RECT 90.680 74.050 91.020 89.170 ;
        RECT 90.680 72.830 91.020 73.750 ;
        RECT 91.340 72.510 91.680 89.170 ;
        RECT 92.000 80.090 92.340 89.170 ;
        RECT 92.000 78.870 92.340 79.790 ;
        RECT 92.000 72.510 92.340 78.570 ;
        RECT 92.660 72.510 93.000 89.170 ;
        RECT 93.320 86.130 93.660 89.170 ;
        RECT 93.320 84.910 93.660 85.830 ;
        RECT 93.320 72.510 93.660 84.610 ;
        RECT 93.980 72.510 94.320 89.170 ;
        RECT 94.640 83.110 94.980 89.170 ;
        RECT 94.640 81.890 94.980 82.810 ;
        RECT 94.640 72.510 94.980 81.590 ;
        RECT 95.300 72.510 95.640 89.170 ;
        RECT 95.960 83.110 96.300 89.170 ;
        RECT 95.960 81.890 96.300 82.810 ;
        RECT 95.960 72.510 96.300 81.590 ;
        RECT 96.620 72.510 96.960 89.170 ;
        RECT 97.280 77.070 97.620 89.170 ;
        RECT 97.280 75.850 97.620 76.770 ;
        RECT 97.280 72.510 97.620 75.550 ;
        RECT 97.940 72.510 98.280 89.170 ;
        RECT 98.600 77.070 98.940 89.170 ;
        RECT 98.600 75.850 98.940 76.770 ;
        RECT 98.600 72.510 98.940 75.550 ;
        RECT 99.260 72.510 99.600 89.170 ;
        RECT 99.920 77.070 100.260 89.170 ;
        RECT 99.920 75.850 100.260 76.770 ;
        RECT 99.920 72.510 100.260 75.550 ;
        RECT 100.580 72.510 100.920 89.170 ;
        RECT 101.240 77.070 101.580 89.170 ;
        RECT 101.240 75.850 101.580 76.770 ;
        RECT 101.240 72.510 101.580 75.550 ;
        RECT 101.900 72.510 102.240 89.170 ;
        RECT 102.560 77.070 102.900 89.170 ;
        RECT 102.560 75.850 102.900 76.770 ;
        RECT 102.560 72.510 102.900 75.550 ;
        RECT 103.220 72.510 103.560 89.170 ;
        RECT 103.880 77.070 104.220 89.170 ;
        RECT 103.880 75.850 104.220 76.770 ;
        RECT 103.880 72.510 104.220 75.550 ;
        RECT 104.540 72.510 104.880 89.170 ;
        RECT 105.200 77.070 105.540 89.170 ;
        RECT 105.200 75.850 105.540 76.770 ;
        RECT 105.200 72.510 105.540 75.550 ;
        RECT 105.860 72.510 106.200 89.170 ;
        RECT 106.520 77.070 106.860 89.170 ;
        RECT 106.520 75.850 106.860 76.770 ;
        RECT 106.520 72.510 106.860 75.550 ;
        RECT 107.180 72.510 107.520 89.170 ;
        RECT 107.840 83.110 108.180 89.170 ;
        RECT 107.840 81.890 108.180 82.810 ;
        RECT 107.840 72.510 108.180 81.590 ;
        RECT 108.500 72.510 108.840 89.170 ;
        RECT 109.160 83.110 109.500 89.170 ;
        RECT 109.160 81.890 109.500 82.810 ;
        RECT 109.160 72.510 109.500 81.590 ;
        RECT 109.820 72.510 110.160 89.170 ;
        RECT 110.480 86.130 110.820 89.170 ;
        RECT 110.480 84.910 110.820 85.830 ;
        RECT 110.480 72.510 110.820 84.610 ;
        RECT 111.140 72.510 111.480 89.170 ;
        RECT 111.800 80.090 112.140 89.170 ;
        RECT 111.800 78.870 112.140 79.790 ;
        RECT 111.800 72.510 112.140 78.570 ;
        RECT 112.460 72.510 112.800 89.170 ;
        RECT 113.120 87.930 113.460 88.850 ;
        RECT 113.120 72.510 113.460 87.630 ;
        RECT 113.780 72.510 114.120 89.170 ;
        RECT 114.440 86.130 114.780 89.170 ;
        RECT 114.440 84.910 114.780 85.830 ;
        RECT 114.440 72.510 114.780 84.610 ;
        RECT 115.100 72.510 115.440 89.170 ;
        RECT 115.760 83.110 116.100 89.170 ;
        RECT 115.760 81.890 116.100 82.810 ;
        RECT 115.760 72.510 116.100 81.590 ;
        RECT 116.420 72.510 116.760 89.170 ;
        RECT 117.080 83.110 117.420 89.170 ;
        RECT 117.080 81.890 117.420 82.810 ;
        RECT 117.080 72.510 117.420 81.590 ;
        RECT 117.740 72.510 118.080 89.170 ;
        RECT 118.400 77.070 118.740 89.170 ;
        RECT 118.400 75.850 118.740 76.770 ;
        RECT 118.400 72.510 118.740 75.550 ;
        RECT 119.060 72.510 119.400 89.170 ;
        RECT 119.720 77.070 120.060 89.170 ;
        RECT 119.720 75.850 120.060 76.770 ;
        RECT 119.720 72.510 120.060 75.550 ;
        RECT 120.380 72.510 120.720 89.170 ;
        RECT 121.040 77.070 121.380 89.170 ;
        RECT 121.040 75.850 121.380 76.770 ;
        RECT 121.040 72.510 121.380 75.550 ;
        RECT 121.700 72.510 122.040 89.170 ;
        RECT 122.360 77.070 122.700 89.170 ;
        RECT 122.360 75.850 122.700 76.770 ;
        RECT 122.360 72.510 122.700 75.550 ;
        RECT 123.020 72.510 123.360 89.170 ;
        RECT 123.680 72.510 124.020 89.170 ;
        RECT 128.630 72.510 128.970 73.090 ;
        RECT 80.780 72.170 128.970 72.510 ;
        RECT 79.220 71.220 80.140 71.560 ;
        RECT 79.220 68.200 80.140 68.540 ;
        RECT 79.220 65.180 80.140 65.520 ;
        RECT 79.220 62.160 80.140 62.500 ;
        RECT 79.220 59.140 80.140 59.480 ;
        RECT 79.220 56.460 79.560 56.750 ;
        RECT 80.780 56.460 81.120 72.170 ;
        RECT 81.440 60.070 81.780 72.170 ;
        RECT 81.440 58.850 81.780 59.770 ;
        RECT 79.220 56.120 81.120 56.460 ;
        RECT 79.220 55.830 79.560 56.120 ;
        RECT 80.780 55.510 81.120 56.120 ;
        RECT 81.440 55.510 81.780 58.550 ;
        RECT 82.100 55.510 82.440 72.170 ;
        RECT 82.760 60.070 83.100 72.170 ;
        RECT 82.760 58.850 83.100 59.770 ;
        RECT 82.760 55.510 83.100 58.550 ;
        RECT 83.420 55.510 83.760 72.170 ;
        RECT 84.080 60.070 84.420 72.170 ;
        RECT 84.080 58.850 84.420 59.770 ;
        RECT 84.080 55.510 84.420 58.550 ;
        RECT 84.740 55.510 85.080 72.170 ;
        RECT 85.400 60.070 85.740 72.170 ;
        RECT 85.400 58.850 85.740 59.770 ;
        RECT 85.400 55.510 85.740 58.550 ;
        RECT 86.060 55.510 86.400 72.170 ;
        RECT 86.720 66.110 87.060 72.170 ;
        RECT 86.720 64.890 87.060 65.810 ;
        RECT 86.720 55.510 87.060 64.590 ;
        RECT 87.380 55.510 87.720 72.170 ;
        RECT 88.040 66.110 88.380 72.170 ;
        RECT 88.040 64.890 88.380 65.810 ;
        RECT 88.040 55.510 88.380 64.590 ;
        RECT 88.700 55.510 89.040 72.170 ;
        RECT 89.360 69.130 89.700 72.170 ;
        RECT 89.360 67.910 89.700 68.830 ;
        RECT 89.360 55.510 89.700 67.610 ;
        RECT 90.020 55.510 90.360 72.170 ;
        RECT 90.680 57.050 91.020 72.170 ;
        RECT 90.680 55.830 91.020 56.750 ;
        RECT 91.340 55.510 91.680 72.170 ;
        RECT 92.000 63.090 92.340 72.170 ;
        RECT 92.000 61.870 92.340 62.790 ;
        RECT 92.000 55.510 92.340 61.570 ;
        RECT 92.660 55.510 93.000 72.170 ;
        RECT 93.320 69.130 93.660 72.170 ;
        RECT 93.320 67.910 93.660 68.830 ;
        RECT 93.320 55.510 93.660 67.610 ;
        RECT 93.980 55.510 94.320 72.170 ;
        RECT 94.640 66.110 94.980 72.170 ;
        RECT 94.640 64.890 94.980 65.810 ;
        RECT 94.640 55.510 94.980 64.590 ;
        RECT 95.300 55.510 95.640 72.170 ;
        RECT 95.960 66.110 96.300 72.170 ;
        RECT 95.960 64.890 96.300 65.810 ;
        RECT 95.960 55.510 96.300 64.590 ;
        RECT 96.620 55.510 96.960 72.170 ;
        RECT 97.280 60.070 97.620 72.170 ;
        RECT 97.280 58.850 97.620 59.770 ;
        RECT 97.280 55.510 97.620 58.550 ;
        RECT 97.940 55.510 98.280 72.170 ;
        RECT 98.600 60.070 98.940 72.170 ;
        RECT 98.600 58.850 98.940 59.770 ;
        RECT 98.600 55.510 98.940 58.550 ;
        RECT 99.260 55.510 99.600 72.170 ;
        RECT 99.920 60.070 100.260 72.170 ;
        RECT 99.920 58.850 100.260 59.770 ;
        RECT 99.920 55.510 100.260 58.550 ;
        RECT 100.580 55.510 100.920 72.170 ;
        RECT 101.240 60.070 101.580 72.170 ;
        RECT 101.240 58.850 101.580 59.770 ;
        RECT 101.240 55.510 101.580 58.550 ;
        RECT 101.900 55.510 102.240 72.170 ;
        RECT 102.560 60.070 102.900 72.170 ;
        RECT 102.560 58.850 102.900 59.770 ;
        RECT 102.560 55.510 102.900 58.550 ;
        RECT 103.220 55.510 103.560 72.170 ;
        RECT 103.880 60.070 104.220 72.170 ;
        RECT 103.880 58.850 104.220 59.770 ;
        RECT 103.880 55.510 104.220 58.550 ;
        RECT 104.540 55.510 104.880 72.170 ;
        RECT 105.200 60.070 105.540 72.170 ;
        RECT 105.200 58.850 105.540 59.770 ;
        RECT 105.200 55.510 105.540 58.550 ;
        RECT 105.860 55.510 106.200 72.170 ;
        RECT 106.520 60.070 106.860 72.170 ;
        RECT 106.520 58.850 106.860 59.770 ;
        RECT 106.520 55.510 106.860 58.550 ;
        RECT 107.180 55.510 107.520 72.170 ;
        RECT 107.840 66.110 108.180 72.170 ;
        RECT 107.840 64.890 108.180 65.810 ;
        RECT 107.840 55.510 108.180 64.590 ;
        RECT 108.500 55.510 108.840 72.170 ;
        RECT 109.160 66.110 109.500 72.170 ;
        RECT 109.160 64.890 109.500 65.810 ;
        RECT 109.160 55.510 109.500 64.590 ;
        RECT 109.820 55.510 110.160 72.170 ;
        RECT 110.480 69.130 110.820 72.170 ;
        RECT 110.480 67.910 110.820 68.830 ;
        RECT 110.480 55.510 110.820 67.610 ;
        RECT 111.140 55.510 111.480 72.170 ;
        RECT 111.800 63.090 112.140 72.170 ;
        RECT 111.800 61.870 112.140 62.790 ;
        RECT 111.800 55.510 112.140 61.570 ;
        RECT 112.460 55.510 112.800 72.170 ;
        RECT 113.120 70.930 113.460 71.850 ;
        RECT 113.120 55.510 113.460 70.630 ;
        RECT 113.780 55.510 114.120 72.170 ;
        RECT 114.440 69.130 114.780 72.170 ;
        RECT 114.440 67.910 114.780 68.830 ;
        RECT 114.440 55.510 114.780 67.610 ;
        RECT 115.100 55.510 115.440 72.170 ;
        RECT 115.760 66.110 116.100 72.170 ;
        RECT 115.760 64.890 116.100 65.810 ;
        RECT 115.760 55.510 116.100 64.590 ;
        RECT 116.420 55.510 116.760 72.170 ;
        RECT 117.080 66.110 117.420 72.170 ;
        RECT 117.080 64.890 117.420 65.810 ;
        RECT 117.080 55.510 117.420 64.590 ;
        RECT 117.740 55.510 118.080 72.170 ;
        RECT 118.400 60.070 118.740 72.170 ;
        RECT 118.400 58.850 118.740 59.770 ;
        RECT 118.400 55.510 118.740 58.550 ;
        RECT 119.060 55.510 119.400 72.170 ;
        RECT 119.720 60.070 120.060 72.170 ;
        RECT 119.720 58.850 120.060 59.770 ;
        RECT 119.720 55.510 120.060 58.550 ;
        RECT 120.380 55.510 120.720 72.170 ;
        RECT 121.040 60.070 121.380 72.170 ;
        RECT 121.040 58.850 121.380 59.770 ;
        RECT 121.040 55.510 121.380 58.550 ;
        RECT 121.700 55.510 122.040 72.170 ;
        RECT 122.360 60.070 122.700 72.170 ;
        RECT 122.360 58.850 122.700 59.770 ;
        RECT 122.360 55.510 122.700 58.550 ;
        RECT 123.020 55.510 123.360 72.170 ;
        RECT 123.680 55.510 124.020 72.170 ;
        RECT 128.630 55.510 128.970 56.090 ;
        RECT 80.780 55.170 128.970 55.510 ;
        RECT 79.220 54.220 80.140 54.560 ;
        RECT 79.220 51.200 80.140 51.540 ;
        RECT 79.220 48.180 80.140 48.520 ;
        RECT 79.220 45.160 80.140 45.500 ;
        RECT 79.220 42.140 80.140 42.480 ;
        RECT 79.220 39.120 80.140 39.460 ;
        RECT 7.290 38.170 55.480 38.510 ;
        RECT 80.780 38.510 81.120 55.170 ;
        RECT 81.440 43.070 81.780 55.170 ;
        RECT 81.440 41.850 81.780 42.770 ;
        RECT 81.440 38.510 81.780 41.550 ;
        RECT 82.100 38.510 82.440 55.170 ;
        RECT 82.760 43.070 83.100 55.170 ;
        RECT 82.760 41.850 83.100 42.770 ;
        RECT 82.760 38.510 83.100 41.550 ;
        RECT 83.420 38.510 83.760 55.170 ;
        RECT 84.080 43.070 84.420 55.170 ;
        RECT 84.080 41.850 84.420 42.770 ;
        RECT 84.080 38.510 84.420 41.550 ;
        RECT 84.740 38.510 85.080 55.170 ;
        RECT 85.400 43.070 85.740 55.170 ;
        RECT 85.400 41.850 85.740 42.770 ;
        RECT 85.400 38.510 85.740 41.550 ;
        RECT 86.060 38.510 86.400 55.170 ;
        RECT 86.720 49.110 87.060 55.170 ;
        RECT 86.720 47.890 87.060 48.810 ;
        RECT 86.720 38.510 87.060 47.590 ;
        RECT 87.380 38.510 87.720 55.170 ;
        RECT 88.040 49.110 88.380 55.170 ;
        RECT 88.040 47.890 88.380 48.810 ;
        RECT 88.040 38.510 88.380 47.590 ;
        RECT 88.700 38.510 89.040 55.170 ;
        RECT 89.360 52.130 89.700 55.170 ;
        RECT 89.360 50.910 89.700 51.830 ;
        RECT 89.360 38.510 89.700 50.610 ;
        RECT 90.020 38.510 90.360 55.170 ;
        RECT 90.680 40.050 91.020 55.170 ;
        RECT 90.680 38.830 91.020 39.750 ;
        RECT 91.340 38.510 91.680 55.170 ;
        RECT 92.000 46.090 92.340 55.170 ;
        RECT 92.000 44.870 92.340 45.790 ;
        RECT 92.000 38.510 92.340 44.570 ;
        RECT 92.660 38.510 93.000 55.170 ;
        RECT 93.320 52.130 93.660 55.170 ;
        RECT 93.320 50.910 93.660 51.830 ;
        RECT 93.320 38.510 93.660 50.610 ;
        RECT 93.980 38.510 94.320 55.170 ;
        RECT 94.640 49.110 94.980 55.170 ;
        RECT 94.640 47.890 94.980 48.810 ;
        RECT 94.640 38.510 94.980 47.590 ;
        RECT 95.300 38.510 95.640 55.170 ;
        RECT 95.960 49.110 96.300 55.170 ;
        RECT 95.960 47.890 96.300 48.810 ;
        RECT 95.960 38.510 96.300 47.590 ;
        RECT 96.620 38.510 96.960 55.170 ;
        RECT 97.280 43.070 97.620 55.170 ;
        RECT 97.280 41.850 97.620 42.770 ;
        RECT 97.280 38.510 97.620 41.550 ;
        RECT 97.940 38.510 98.280 55.170 ;
        RECT 98.600 43.070 98.940 55.170 ;
        RECT 98.600 41.850 98.940 42.770 ;
        RECT 98.600 38.510 98.940 41.550 ;
        RECT 99.260 38.510 99.600 55.170 ;
        RECT 99.920 43.070 100.260 55.170 ;
        RECT 99.920 41.850 100.260 42.770 ;
        RECT 99.920 38.510 100.260 41.550 ;
        RECT 100.580 38.510 100.920 55.170 ;
        RECT 101.240 43.070 101.580 55.170 ;
        RECT 101.240 41.850 101.580 42.770 ;
        RECT 101.240 38.510 101.580 41.550 ;
        RECT 101.900 38.510 102.240 55.170 ;
        RECT 102.560 43.070 102.900 55.170 ;
        RECT 102.560 41.850 102.900 42.770 ;
        RECT 102.560 38.510 102.900 41.550 ;
        RECT 103.220 38.510 103.560 55.170 ;
        RECT 103.880 43.070 104.220 55.170 ;
        RECT 103.880 41.850 104.220 42.770 ;
        RECT 103.880 38.510 104.220 41.550 ;
        RECT 104.540 38.510 104.880 55.170 ;
        RECT 105.200 43.070 105.540 55.170 ;
        RECT 105.200 41.850 105.540 42.770 ;
        RECT 105.200 38.510 105.540 41.550 ;
        RECT 105.860 38.510 106.200 55.170 ;
        RECT 106.520 43.070 106.860 55.170 ;
        RECT 106.520 41.850 106.860 42.770 ;
        RECT 106.520 38.510 106.860 41.550 ;
        RECT 107.180 38.510 107.520 55.170 ;
        RECT 107.840 49.110 108.180 55.170 ;
        RECT 107.840 47.890 108.180 48.810 ;
        RECT 107.840 38.510 108.180 47.590 ;
        RECT 108.500 38.510 108.840 55.170 ;
        RECT 109.160 49.110 109.500 55.170 ;
        RECT 109.160 47.890 109.500 48.810 ;
        RECT 109.160 38.510 109.500 47.590 ;
        RECT 109.820 38.510 110.160 55.170 ;
        RECT 110.480 52.130 110.820 55.170 ;
        RECT 110.480 50.910 110.820 51.830 ;
        RECT 110.480 38.510 110.820 50.610 ;
        RECT 111.140 38.510 111.480 55.170 ;
        RECT 111.800 46.090 112.140 55.170 ;
        RECT 111.800 44.870 112.140 45.790 ;
        RECT 111.800 38.510 112.140 44.570 ;
        RECT 112.460 38.510 112.800 55.170 ;
        RECT 113.120 53.930 113.460 54.850 ;
        RECT 113.120 38.510 113.460 53.630 ;
        RECT 113.780 38.510 114.120 55.170 ;
        RECT 114.440 52.130 114.780 55.170 ;
        RECT 114.440 50.910 114.780 51.830 ;
        RECT 114.440 38.510 114.780 50.610 ;
        RECT 115.100 38.510 115.440 55.170 ;
        RECT 115.760 49.110 116.100 55.170 ;
        RECT 115.760 47.890 116.100 48.810 ;
        RECT 115.760 38.510 116.100 47.590 ;
        RECT 116.420 38.510 116.760 55.170 ;
        RECT 117.080 49.110 117.420 55.170 ;
        RECT 117.080 47.890 117.420 48.810 ;
        RECT 117.080 38.510 117.420 47.590 ;
        RECT 117.740 38.510 118.080 55.170 ;
        RECT 118.400 43.070 118.740 55.170 ;
        RECT 118.400 41.850 118.740 42.770 ;
        RECT 118.400 38.510 118.740 41.550 ;
        RECT 119.060 38.510 119.400 55.170 ;
        RECT 119.720 43.070 120.060 55.170 ;
        RECT 119.720 41.850 120.060 42.770 ;
        RECT 119.720 38.510 120.060 41.550 ;
        RECT 120.380 38.510 120.720 55.170 ;
        RECT 121.040 43.070 121.380 55.170 ;
        RECT 121.040 41.850 121.380 42.770 ;
        RECT 121.040 38.510 121.380 41.550 ;
        RECT 121.700 38.510 122.040 55.170 ;
        RECT 122.360 43.070 122.700 55.170 ;
        RECT 122.360 41.850 122.700 42.770 ;
        RECT 122.360 38.510 122.700 41.550 ;
        RECT 123.020 38.510 123.360 55.170 ;
        RECT 123.680 38.510 124.020 55.170 ;
        RECT 128.630 38.510 128.970 39.090 ;
        RECT 80.780 38.170 128.970 38.510 ;
        RECT 11.070 36.240 46.710 36.640 ;
        RECT 11.070 35.440 45.990 35.840 ;
        RECT 11.070 34.240 11.430 35.440 ;
        RECT 46.350 35.040 46.710 36.240 ;
        RECT 11.790 34.640 46.710 35.040 ;
        RECT 11.070 33.840 45.990 34.240 ;
        RECT 11.070 32.640 11.430 33.840 ;
        RECT 46.350 33.440 46.710 34.640 ;
        RECT 11.790 33.040 46.710 33.440 ;
        RECT 89.550 36.240 125.190 36.640 ;
        RECT 89.550 35.040 89.910 36.240 ;
        RECT 90.270 35.440 125.190 35.840 ;
        RECT 89.550 34.640 124.470 35.040 ;
        RECT 89.550 33.440 89.910 34.640 ;
        RECT 124.830 34.240 125.190 35.440 ;
        RECT 90.270 33.840 125.190 34.240 ;
        RECT 89.550 33.040 124.470 33.440 ;
        RECT 124.830 32.640 125.190 33.840 ;
        RECT 11.070 32.240 46.710 32.640 ;
        RECT 89.550 32.240 125.190 32.640 ;
        RECT 11.070 31.440 46.710 31.840 ;
        RECT 11.070 30.640 45.990 31.040 ;
        RECT 11.070 29.440 11.430 30.640 ;
        RECT 46.350 30.240 46.710 31.440 ;
        RECT 11.790 29.840 46.710 30.240 ;
        RECT 11.070 29.040 45.990 29.440 ;
        RECT 11.070 27.840 11.430 29.040 ;
        RECT 46.350 28.640 46.710 29.840 ;
        RECT 89.550 31.440 125.190 31.840 ;
        RECT 89.550 30.240 89.910 31.440 ;
        RECT 90.270 30.640 125.190 31.040 ;
        RECT 89.550 29.840 124.470 30.240 ;
        RECT 52.270 29.350 53.190 29.690 ;
        RECT 56.230 29.350 57.150 29.690 ;
        RECT 79.110 29.350 80.030 29.690 ;
        RECT 83.070 29.350 83.990 29.690 ;
        RECT 11.790 28.240 46.710 28.640 ;
        RECT 52.270 28.470 53.190 28.810 ;
        RECT 56.230 28.470 57.150 28.810 ;
        RECT 79.110 28.470 80.030 28.810 ;
        RECT 83.070 28.470 83.990 28.810 ;
        RECT 89.550 28.640 89.910 29.840 ;
        RECT 124.830 29.440 125.190 30.640 ;
        RECT 90.270 29.040 125.190 29.440 ;
        RECT 89.550 28.240 124.470 28.640 ;
        RECT 11.070 27.440 46.710 27.840 ;
        RECT 56.230 27.590 65.130 27.930 ;
        RECT 11.070 26.640 46.710 27.040 ;
        RECT 52.270 26.710 53.190 27.050 ;
        RECT 56.230 26.710 57.150 27.050 ;
        RECT 11.070 25.840 45.990 26.240 ;
        RECT 11.070 24.640 11.430 25.840 ;
        RECT 46.350 25.440 46.710 26.640 ;
        RECT 64.790 26.610 65.130 27.590 ;
        RECT 71.130 27.590 80.030 27.930 ;
        RECT 124.830 27.840 125.190 29.040 ;
        RECT 71.130 26.610 71.470 27.590 ;
        RECT 89.550 27.440 125.190 27.840 ;
        RECT 79.110 26.710 80.030 27.050 ;
        RECT 83.070 26.710 83.990 27.050 ;
        RECT 64.790 26.270 66.510 26.610 ;
        RECT 69.750 26.270 71.470 26.610 ;
        RECT 89.550 26.640 125.190 27.040 ;
        RECT 52.270 25.830 53.190 26.170 ;
        RECT 56.230 25.830 57.150 26.170 ;
        RECT 63.270 25.830 64.190 26.170 ;
        RECT 71.910 25.830 72.830 26.170 ;
        RECT 79.110 25.830 80.030 26.170 ;
        RECT 83.070 25.830 83.990 26.170 ;
        RECT 11.790 25.040 46.710 25.440 ;
        RECT 89.550 25.440 89.910 26.640 ;
        RECT 90.270 25.840 125.190 26.240 ;
        RECT 11.070 24.240 45.990 24.640 ;
        RECT 11.070 23.040 11.430 24.240 ;
        RECT 46.350 23.840 46.710 25.040 ;
        RECT 52.270 24.950 53.190 25.290 ;
        RECT 56.230 24.950 57.150 25.290 ;
        RECT 79.110 24.950 80.030 25.290 ;
        RECT 83.070 24.950 83.990 25.290 ;
        RECT 89.550 25.040 124.470 25.440 ;
        RECT 52.270 24.240 57.930 24.580 ;
        RECT 11.790 23.440 46.710 23.840 ;
        RECT 52.270 23.190 53.190 23.530 ;
        RECT 56.230 23.190 57.150 23.530 ;
        RECT 11.070 22.640 46.710 23.040 ;
        RECT 52.270 22.310 53.190 22.650 ;
        RECT 56.070 22.310 56.990 22.650 ;
        RECT 11.070 21.840 46.710 22.240 ;
        RECT 57.590 22.210 57.930 24.240 ;
        RECT 78.330 24.240 83.990 24.580 ;
        RECT 78.330 22.210 78.670 24.240 ;
        RECT 89.550 23.840 89.910 25.040 ;
        RECT 124.830 24.640 125.190 25.840 ;
        RECT 90.270 24.240 125.190 24.640 ;
        RECT 79.110 23.190 80.030 23.530 ;
        RECT 83.070 23.190 83.990 23.530 ;
        RECT 89.550 23.440 124.470 23.840 ;
        RECT 124.830 23.040 125.190 24.240 ;
        RECT 79.270 22.310 80.190 22.650 ;
        RECT 83.070 22.310 83.990 22.650 ;
        RECT 89.550 22.640 125.190 23.040 ;
        RECT 57.590 21.870 59.310 22.210 ;
        RECT 76.950 21.870 78.670 22.210 ;
        RECT 11.070 21.040 45.990 21.440 ;
        RECT 11.070 19.840 11.430 21.040 ;
        RECT 46.350 20.640 46.710 21.840 ;
        RECT 89.550 21.840 125.190 22.240 ;
        RECT 50.110 21.430 53.190 21.770 ;
        RECT 83.070 21.430 86.150 21.770 ;
        RECT 58.390 20.990 59.310 21.330 ;
        RECT 76.950 20.990 77.870 21.330 ;
        RECT 11.790 20.240 46.710 20.640 ;
        RECT 56.230 20.550 57.150 20.890 ;
        RECT 79.110 20.550 80.030 20.890 ;
        RECT 89.550 20.640 89.910 21.840 ;
        RECT 90.270 21.040 125.190 21.440 ;
        RECT 11.070 19.440 45.990 19.840 ;
        RECT 11.070 18.240 11.430 19.440 ;
        RECT 46.350 19.040 46.710 20.240 ;
        RECT 89.550 20.240 124.470 20.640 ;
        RECT 56.230 19.670 62.970 20.010 ;
        RECT 11.790 18.640 46.710 19.040 ;
        RECT 52.270 18.790 53.190 19.130 ;
        RECT 50.110 18.350 51.030 18.690 ;
        RECT 62.630 18.250 62.970 19.670 ;
        RECT 73.290 19.670 80.030 20.010 ;
        RECT 63.270 18.790 64.190 19.130 ;
        RECT 71.910 18.790 72.830 19.130 ;
        RECT 73.290 18.250 73.630 19.670 ;
        RECT 83.070 18.790 83.990 19.130 ;
        RECT 89.550 19.040 89.910 20.240 ;
        RECT 124.830 19.840 125.190 21.040 ;
        RECT 90.270 19.440 125.190 19.840 ;
        RECT 85.230 18.350 86.150 18.690 ;
        RECT 89.550 18.640 124.470 19.040 ;
        RECT 11.070 17.840 46.710 18.240 ;
        RECT 52.270 17.910 53.190 18.250 ;
        RECT 56.230 17.910 57.150 18.250 ;
        RECT 62.630 17.910 64.350 18.250 ;
        RECT 71.910 17.910 73.630 18.250 ;
        RECT 79.110 17.910 80.030 18.250 ;
        RECT 83.070 17.910 83.990 18.250 ;
        RECT 124.830 18.240 125.190 19.440 ;
        RECT 89.550 17.840 125.190 18.240 ;
        RECT 50.110 17.470 51.810 17.810 ;
        RECT 65.430 17.470 66.350 17.810 ;
        RECT 69.910 17.470 70.830 17.810 ;
        RECT 84.450 17.470 86.150 17.810 ;
        RECT 11.070 17.040 46.710 17.440 ;
        RECT 11.070 16.240 45.990 16.640 ;
        RECT 11.070 15.040 11.430 16.240 ;
        RECT 46.350 15.840 46.710 17.040 ;
        RECT 51.470 16.490 51.810 17.470 ;
        RECT 51.470 16.150 53.190 16.490 ;
        RECT 56.230 16.320 57.150 16.660 ;
        RECT 79.110 16.320 80.030 16.660 ;
        RECT 84.450 16.490 84.790 17.470 ;
        RECT 83.070 16.150 84.790 16.490 ;
        RECT 89.550 17.040 125.190 17.440 ;
        RECT 11.790 15.440 46.710 15.840 ;
        RECT 58.310 15.710 59.230 16.050 ;
        RECT 77.030 15.710 77.950 16.050 ;
        RECT 89.550 15.840 89.910 17.040 ;
        RECT 90.270 16.240 125.190 16.640 ;
        RECT 11.070 14.640 45.990 15.040 ;
        RECT 11.070 13.440 11.430 14.640 ;
        RECT 46.350 14.240 46.710 15.440 ;
        RECT 52.270 15.270 53.190 15.610 ;
        RECT 56.230 15.270 57.150 15.610 ;
        RECT 52.270 14.390 53.190 14.730 ;
        RECT 56.230 14.390 57.150 14.730 ;
        RECT 11.790 13.840 46.710 14.240 ;
        RECT 52.270 13.510 53.190 13.850 ;
        RECT 56.230 13.510 57.150 13.850 ;
        RECT 11.070 13.040 46.710 13.440 ;
        RECT 56.230 9.640 57.150 10.560 ;
        RECT 52.270 6.040 53.190 6.960 ;
        RECT 58.600 5.320 58.940 15.710 ;
        RECT 63.270 14.390 64.190 14.730 ;
        RECT 72.070 14.390 72.990 14.730 ;
        RECT 77.320 5.320 77.660 15.710 ;
        RECT 79.110 15.270 80.030 15.610 ;
        RECT 83.070 15.270 83.990 15.610 ;
        RECT 89.550 15.440 124.470 15.840 ;
        RECT 79.110 14.390 80.030 14.730 ;
        RECT 83.070 14.390 83.990 14.730 ;
        RECT 89.550 14.240 89.910 15.440 ;
        RECT 124.830 15.040 125.190 16.240 ;
        RECT 90.270 14.640 125.190 15.040 ;
        RECT 79.110 13.510 80.030 13.850 ;
        RECT 83.070 13.510 83.990 13.850 ;
        RECT 89.550 13.840 124.470 14.240 ;
        RECT 124.830 13.440 125.190 14.640 ;
        RECT 89.550 13.040 125.190 13.440 ;
        RECT 79.110 9.640 80.030 10.560 ;
        RECT 83.070 6.040 83.990 6.960 ;
        RECT 58.310 4.980 59.230 5.320 ;
        RECT 77.030 4.980 77.950 5.320 ;
        RECT 58.830 3.920 59.750 4.260 ;
        RECT 76.510 3.920 77.430 4.260 ;
      LAYER via ;
        RECT 59.695 224.020 59.995 224.320 ;
        RECT 61.210 224.160 61.510 224.460 ;
        RECT 86.880 222.410 87.180 222.710 ;
        RECT 116.500 222.410 116.800 222.710 ;
        RECT 116.250 221.230 116.530 221.510 ;
        RECT 116.770 221.230 117.050 221.510 ;
        RECT 15.450 220.350 15.730 220.630 ;
        RECT 15.970 220.350 16.250 220.630 ;
        RECT 15.370 219.470 15.650 219.750 ;
        RECT 15.890 219.470 16.170 219.750 ;
        RECT 19.330 219.470 19.610 219.750 ;
        RECT 19.850 219.470 20.130 219.750 ;
        RECT 32.010 220.350 32.290 220.630 ;
        RECT 32.530 220.350 32.810 220.630 ;
        RECT 40.650 220.350 40.930 220.630 ;
        RECT 41.170 220.350 41.450 220.630 ;
        RECT 28.130 219.470 28.410 219.750 ;
        RECT 28.650 219.470 28.930 219.750 ;
        RECT 32.090 219.470 32.370 219.750 ;
        RECT 32.610 219.470 32.890 219.750 ;
        RECT 40.570 219.470 40.850 219.750 ;
        RECT 41.090 219.470 41.370 219.750 ;
        RECT 44.530 219.470 44.810 219.750 ;
        RECT 45.050 219.470 45.330 219.750 ;
        RECT 15.370 216.830 15.650 217.110 ;
        RECT 15.890 216.830 16.170 217.110 ;
        RECT 19.330 216.830 19.610 217.110 ;
        RECT 19.850 216.830 20.130 217.110 ;
        RECT 28.130 216.830 28.410 217.110 ;
        RECT 28.650 216.830 28.930 217.110 ;
        RECT 32.090 216.830 32.370 217.110 ;
        RECT 32.610 216.830 32.890 217.110 ;
        RECT 15.370 214.190 15.650 214.470 ;
        RECT 15.890 214.190 16.170 214.470 ;
        RECT 19.330 214.190 19.610 214.470 ;
        RECT 19.850 214.190 20.130 214.470 ;
        RECT 15.370 212.430 15.650 212.710 ;
        RECT 15.890 212.430 16.170 212.710 ;
        RECT 19.330 212.430 19.610 212.710 ;
        RECT 19.850 212.430 20.130 212.710 ;
        RECT 15.370 209.790 15.650 210.070 ;
        RECT 15.890 209.790 16.170 210.070 ;
        RECT 19.330 209.790 19.610 210.070 ;
        RECT 19.850 209.790 20.130 210.070 ;
        RECT 13.290 207.590 13.570 207.870 ;
        RECT 13.810 207.590 14.090 207.870 ;
        RECT 15.370 207.150 15.650 207.430 ;
        RECT 15.890 207.150 16.170 207.430 ;
        RECT 19.330 207.150 19.610 207.430 ;
        RECT 19.850 207.150 20.130 207.430 ;
        RECT 15.370 205.390 15.650 205.670 ;
        RECT 15.890 205.390 16.170 205.670 ;
        RECT 19.330 205.390 19.610 205.670 ;
        RECT 19.850 205.390 20.130 205.670 ;
        RECT 57.210 220.350 57.490 220.630 ;
        RECT 57.730 220.350 58.010 220.630 ;
        RECT 65.850 220.350 66.130 220.630 ;
        RECT 66.370 220.350 66.650 220.630 ;
        RECT 53.330 219.470 53.610 219.750 ;
        RECT 53.850 219.470 54.130 219.750 ;
        RECT 57.290 219.470 57.570 219.750 ;
        RECT 57.810 219.470 58.090 219.750 ;
        RECT 65.770 219.470 66.050 219.750 ;
        RECT 66.290 219.470 66.570 219.750 ;
        RECT 69.730 219.470 70.010 219.750 ;
        RECT 70.250 219.470 70.530 219.750 ;
        RECT 40.570 216.830 40.850 217.110 ;
        RECT 41.090 216.830 41.370 217.110 ;
        RECT 44.530 216.830 44.810 217.110 ;
        RECT 45.050 216.830 45.330 217.110 ;
        RECT 53.330 216.830 53.610 217.110 ;
        RECT 53.850 216.830 54.130 217.110 ;
        RECT 57.290 216.830 57.570 217.110 ;
        RECT 57.810 216.830 58.090 217.110 ;
        RECT 28.130 214.190 28.410 214.470 ;
        RECT 28.650 214.190 28.930 214.470 ;
        RECT 32.090 214.190 32.370 214.470 ;
        RECT 32.610 214.190 32.890 214.470 ;
        RECT 40.570 214.190 40.850 214.470 ;
        RECT 41.090 214.190 41.370 214.470 ;
        RECT 44.530 214.190 44.810 214.470 ;
        RECT 45.050 214.190 45.330 214.470 ;
        RECT 28.130 212.430 28.410 212.710 ;
        RECT 28.650 212.430 28.930 212.710 ;
        RECT 32.090 212.430 32.370 212.710 ;
        RECT 32.610 212.430 32.890 212.710 ;
        RECT 40.570 212.430 40.850 212.710 ;
        RECT 41.090 212.430 41.370 212.710 ;
        RECT 44.530 212.430 44.810 212.710 ;
        RECT 45.050 212.430 45.330 212.710 ;
        RECT 28.130 209.790 28.410 210.070 ;
        RECT 28.650 209.790 28.930 210.070 ;
        RECT 32.090 209.790 32.370 210.070 ;
        RECT 32.610 209.790 32.890 210.070 ;
        RECT 40.570 209.790 40.850 210.070 ;
        RECT 41.090 209.790 41.370 210.070 ;
        RECT 44.530 209.790 44.810 210.070 ;
        RECT 45.050 209.790 45.330 210.070 ;
        RECT 28.130 207.150 28.410 207.430 ;
        RECT 28.650 207.150 28.930 207.430 ;
        RECT 32.090 207.150 32.370 207.430 ;
        RECT 32.610 207.150 32.890 207.430 ;
        RECT 28.130 205.390 28.410 205.670 ;
        RECT 28.650 205.390 28.930 205.670 ;
        RECT 32.090 205.390 32.370 205.670 ;
        RECT 32.610 205.390 32.890 205.670 ;
        RECT 34.170 207.590 34.450 207.870 ;
        RECT 34.690 207.590 34.970 207.870 ;
        RECT 38.490 207.590 38.770 207.870 ;
        RECT 39.010 207.590 39.290 207.870 ;
        RECT 40.570 207.150 40.850 207.430 ;
        RECT 41.090 207.150 41.370 207.430 ;
        RECT 44.530 207.150 44.810 207.430 ;
        RECT 45.050 207.150 45.330 207.430 ;
        RECT 40.570 205.390 40.850 205.670 ;
        RECT 41.090 205.390 41.370 205.670 ;
        RECT 44.530 205.390 44.810 205.670 ;
        RECT 45.050 205.390 45.330 205.670 ;
        RECT 82.410 220.350 82.690 220.630 ;
        RECT 82.930 220.350 83.210 220.630 ;
        RECT 91.050 220.350 91.330 220.630 ;
        RECT 91.570 220.350 91.850 220.630 ;
        RECT 78.530 219.470 78.810 219.750 ;
        RECT 79.050 219.470 79.330 219.750 ;
        RECT 82.490 219.470 82.770 219.750 ;
        RECT 83.010 219.470 83.290 219.750 ;
        RECT 90.970 219.470 91.250 219.750 ;
        RECT 91.490 219.470 91.770 219.750 ;
        RECT 94.930 219.470 95.210 219.750 ;
        RECT 95.450 219.470 95.730 219.750 ;
        RECT 65.770 216.830 66.050 217.110 ;
        RECT 66.290 216.830 66.570 217.110 ;
        RECT 69.730 216.830 70.010 217.110 ;
        RECT 70.250 216.830 70.530 217.110 ;
        RECT 78.530 216.830 78.810 217.110 ;
        RECT 79.050 216.830 79.330 217.110 ;
        RECT 82.490 216.830 82.770 217.110 ;
        RECT 83.010 216.830 83.290 217.110 ;
        RECT 53.330 214.190 53.610 214.470 ;
        RECT 53.850 214.190 54.130 214.470 ;
        RECT 57.290 214.190 57.570 214.470 ;
        RECT 57.810 214.190 58.090 214.470 ;
        RECT 65.770 214.190 66.050 214.470 ;
        RECT 66.290 214.190 66.570 214.470 ;
        RECT 69.730 214.190 70.010 214.470 ;
        RECT 70.250 214.190 70.530 214.470 ;
        RECT 53.330 212.430 53.610 212.710 ;
        RECT 53.850 212.430 54.130 212.710 ;
        RECT 57.290 212.430 57.570 212.710 ;
        RECT 57.810 212.430 58.090 212.710 ;
        RECT 65.770 212.430 66.050 212.710 ;
        RECT 66.290 212.430 66.570 212.710 ;
        RECT 69.730 212.430 70.010 212.710 ;
        RECT 70.250 212.430 70.530 212.710 ;
        RECT 53.330 209.790 53.610 210.070 ;
        RECT 53.850 209.790 54.130 210.070 ;
        RECT 57.290 209.790 57.570 210.070 ;
        RECT 57.810 209.790 58.090 210.070 ;
        RECT 65.770 209.790 66.050 210.070 ;
        RECT 66.290 209.790 66.570 210.070 ;
        RECT 69.730 209.790 70.010 210.070 ;
        RECT 70.250 209.790 70.530 210.070 ;
        RECT 53.330 207.150 53.610 207.430 ;
        RECT 53.850 207.150 54.130 207.430 ;
        RECT 57.290 207.150 57.570 207.430 ;
        RECT 57.810 207.150 58.090 207.430 ;
        RECT 53.330 205.390 53.610 205.670 ;
        RECT 53.850 205.390 54.130 205.670 ;
        RECT 57.290 205.390 57.570 205.670 ;
        RECT 57.810 205.390 58.090 205.670 ;
        RECT 59.370 207.590 59.650 207.870 ;
        RECT 59.890 207.590 60.170 207.870 ;
        RECT 63.690 207.590 63.970 207.870 ;
        RECT 64.210 207.590 64.490 207.870 ;
        RECT 65.770 207.150 66.050 207.430 ;
        RECT 66.290 207.150 66.570 207.430 ;
        RECT 69.730 207.150 70.010 207.430 ;
        RECT 70.250 207.150 70.530 207.430 ;
        RECT 65.770 205.390 66.050 205.670 ;
        RECT 66.290 205.390 66.570 205.670 ;
        RECT 69.730 205.390 70.010 205.670 ;
        RECT 70.250 205.390 70.530 205.670 ;
        RECT 107.610 220.350 107.890 220.630 ;
        RECT 108.130 220.350 108.410 220.630 ;
        RECT 116.170 220.350 116.450 220.630 ;
        RECT 116.690 220.350 116.970 220.630 ;
        RECT 120.130 220.350 120.410 220.630 ;
        RECT 120.650 220.350 120.930 220.630 ;
        RECT 103.730 219.470 104.010 219.750 ;
        RECT 104.250 219.470 104.530 219.750 ;
        RECT 107.690 219.470 107.970 219.750 ;
        RECT 108.210 219.470 108.490 219.750 ;
        RECT 116.170 219.470 116.450 219.750 ;
        RECT 116.690 219.470 116.970 219.750 ;
        RECT 132.530 219.430 132.870 219.770 ;
        RECT 116.170 218.590 116.450 218.870 ;
        RECT 116.690 218.590 116.970 218.870 ;
        RECT 120.130 218.590 120.410 218.870 ;
        RECT 120.650 218.590 120.930 218.870 ;
        RECT 90.970 216.830 91.250 217.110 ;
        RECT 91.490 216.830 91.770 217.110 ;
        RECT 94.930 216.830 95.210 217.110 ;
        RECT 95.450 216.830 95.730 217.110 ;
        RECT 103.730 216.830 104.010 217.110 ;
        RECT 104.250 216.830 104.530 217.110 ;
        RECT 107.690 216.830 107.970 217.110 ;
        RECT 108.210 216.830 108.490 217.110 ;
        RECT 120.130 217.710 120.410 217.990 ;
        RECT 120.650 217.710 120.930 217.990 ;
        RECT 114.170 216.390 114.450 216.670 ;
        RECT 114.690 216.390 114.970 216.670 ;
        RECT 116.170 215.950 116.450 216.230 ;
        RECT 116.690 215.950 116.970 216.230 ;
        RECT 78.530 214.190 78.810 214.470 ;
        RECT 79.050 214.190 79.330 214.470 ;
        RECT 82.490 214.190 82.770 214.470 ;
        RECT 83.010 214.190 83.290 214.470 ;
        RECT 90.970 214.190 91.250 214.470 ;
        RECT 91.490 214.190 91.770 214.470 ;
        RECT 94.930 214.190 95.210 214.470 ;
        RECT 95.450 214.190 95.730 214.470 ;
        RECT 78.530 212.430 78.810 212.710 ;
        RECT 79.050 212.430 79.330 212.710 ;
        RECT 82.490 212.430 82.770 212.710 ;
        RECT 83.010 212.430 83.290 212.710 ;
        RECT 90.970 212.430 91.250 212.710 ;
        RECT 91.490 212.430 91.770 212.710 ;
        RECT 94.930 212.430 95.210 212.710 ;
        RECT 95.450 212.430 95.730 212.710 ;
        RECT 78.530 209.790 78.810 210.070 ;
        RECT 79.050 209.790 79.330 210.070 ;
        RECT 82.490 209.790 82.770 210.070 ;
        RECT 83.010 209.790 83.290 210.070 ;
        RECT 90.970 209.790 91.250 210.070 ;
        RECT 91.490 209.790 91.770 210.070 ;
        RECT 94.930 209.790 95.210 210.070 ;
        RECT 95.450 209.790 95.730 210.070 ;
        RECT 78.530 207.150 78.810 207.430 ;
        RECT 79.050 207.150 79.330 207.430 ;
        RECT 82.490 207.150 82.770 207.430 ;
        RECT 83.010 207.150 83.290 207.430 ;
        RECT 78.530 205.390 78.810 205.670 ;
        RECT 79.050 205.390 79.330 205.670 ;
        RECT 82.490 205.390 82.770 205.670 ;
        RECT 83.010 205.390 83.290 205.670 ;
        RECT 84.570 207.590 84.850 207.870 ;
        RECT 85.090 207.590 85.370 207.870 ;
        RECT 88.890 207.590 89.170 207.870 ;
        RECT 89.410 207.590 89.690 207.870 ;
        RECT 90.970 207.150 91.250 207.430 ;
        RECT 91.490 207.150 91.770 207.430 ;
        RECT 94.930 207.150 95.210 207.430 ;
        RECT 95.450 207.150 95.730 207.430 ;
        RECT 90.970 205.390 91.250 205.670 ;
        RECT 91.490 205.390 91.770 205.670 ;
        RECT 94.930 205.390 95.210 205.670 ;
        RECT 95.450 205.390 95.730 205.670 ;
        RECT 116.170 215.070 116.450 215.350 ;
        RECT 116.690 215.070 116.970 215.350 ;
        RECT 103.730 214.190 104.010 214.470 ;
        RECT 104.250 214.190 104.530 214.470 ;
        RECT 107.690 214.190 107.970 214.470 ;
        RECT 108.210 214.190 108.490 214.470 ;
        RECT 116.170 214.190 116.450 214.470 ;
        RECT 116.690 214.190 116.970 214.470 ;
        RECT 116.170 213.310 116.450 213.590 ;
        RECT 116.690 213.310 116.970 213.590 ;
        RECT 103.730 212.430 104.010 212.710 ;
        RECT 104.250 212.430 104.530 212.710 ;
        RECT 107.690 212.430 107.970 212.710 ;
        RECT 108.210 212.430 108.490 212.710 ;
        RECT 116.170 212.430 116.450 212.710 ;
        RECT 116.690 212.430 116.970 212.710 ;
        RECT 116.170 211.550 116.450 211.830 ;
        RECT 116.690 211.550 116.970 211.830 ;
        RECT 114.170 210.230 114.450 210.510 ;
        RECT 114.690 210.230 114.970 210.510 ;
        RECT 103.730 209.790 104.010 210.070 ;
        RECT 104.250 209.790 104.530 210.070 ;
        RECT 107.690 209.790 107.970 210.070 ;
        RECT 108.210 209.790 108.490 210.070 ;
        RECT 103.730 207.150 104.010 207.430 ;
        RECT 104.250 207.150 104.530 207.430 ;
        RECT 107.690 207.150 107.970 207.430 ;
        RECT 108.210 207.150 108.490 207.430 ;
        RECT 103.730 205.390 104.010 205.670 ;
        RECT 104.250 205.390 104.530 205.670 ;
        RECT 107.690 205.390 107.970 205.670 ;
        RECT 108.210 205.390 108.490 205.670 ;
        RECT 109.770 207.590 110.050 207.870 ;
        RECT 110.290 207.590 110.570 207.870 ;
        RECT 114.010 207.590 114.290 207.870 ;
        RECT 114.530 207.590 114.810 207.870 ;
        RECT 116.170 209.790 116.450 210.070 ;
        RECT 116.690 209.790 116.970 210.070 ;
        RECT 116.330 208.910 116.610 209.190 ;
        RECT 116.850 208.910 117.130 209.190 ;
        RECT 116.170 208.030 116.450 208.310 ;
        RECT 116.690 208.030 116.970 208.310 ;
        RECT 120.130 215.950 120.410 216.230 ;
        RECT 120.650 215.950 120.930 216.230 ;
        RECT 120.130 214.190 120.410 214.470 ;
        RECT 120.650 214.190 120.930 214.470 ;
        RECT 126.710 213.230 127.050 213.570 ;
        RECT 120.130 212.430 120.410 212.710 ;
        RECT 120.650 212.430 120.930 212.710 ;
        RECT 120.130 209.790 120.410 210.070 ;
        RECT 120.650 209.790 120.930 210.070 ;
        RECT 120.130 208.030 120.410 208.310 ;
        RECT 120.650 208.030 120.930 208.310 ;
        RECT 116.170 205.390 116.450 205.670 ;
        RECT 116.690 205.390 116.970 205.670 ;
        RECT 120.130 205.390 120.410 205.670 ;
        RECT 120.650 205.390 120.930 205.670 ;
        RECT 114.170 204.070 114.450 204.350 ;
        RECT 114.690 204.070 114.970 204.350 ;
        RECT 15.370 203.630 15.650 203.910 ;
        RECT 15.890 203.630 16.170 203.910 ;
        RECT 19.330 203.630 19.610 203.910 ;
        RECT 19.850 203.630 20.130 203.910 ;
        RECT 28.130 203.630 28.410 203.910 ;
        RECT 28.650 203.630 28.930 203.910 ;
        RECT 32.090 203.630 32.370 203.910 ;
        RECT 32.610 203.630 32.890 203.910 ;
        RECT 15.370 202.750 15.650 203.030 ;
        RECT 15.890 202.750 16.170 203.030 ;
        RECT 19.330 202.750 19.610 203.030 ;
        RECT 19.850 202.750 20.130 203.030 ;
        RECT 28.130 202.750 28.410 203.030 ;
        RECT 28.650 202.750 28.930 203.030 ;
        RECT 32.090 202.750 32.370 203.030 ;
        RECT 32.610 202.750 32.890 203.030 ;
        RECT 15.370 201.870 15.650 202.150 ;
        RECT 15.890 201.870 16.170 202.150 ;
        RECT 19.330 201.870 19.610 202.150 ;
        RECT 19.850 201.870 20.130 202.150 ;
        RECT 28.130 201.870 28.410 202.150 ;
        RECT 28.650 201.870 28.930 202.150 ;
        RECT 32.090 201.870 32.370 202.150 ;
        RECT 32.610 201.870 32.890 202.150 ;
        RECT 40.570 203.630 40.850 203.910 ;
        RECT 41.090 203.630 41.370 203.910 ;
        RECT 44.530 203.630 44.810 203.910 ;
        RECT 45.050 203.630 45.330 203.910 ;
        RECT 53.330 203.630 53.610 203.910 ;
        RECT 53.850 203.630 54.130 203.910 ;
        RECT 57.290 203.630 57.570 203.910 ;
        RECT 57.810 203.630 58.090 203.910 ;
        RECT 40.570 202.750 40.850 203.030 ;
        RECT 41.090 202.750 41.370 203.030 ;
        RECT 44.530 202.750 44.810 203.030 ;
        RECT 45.050 202.750 45.330 203.030 ;
        RECT 53.330 202.750 53.610 203.030 ;
        RECT 53.850 202.750 54.130 203.030 ;
        RECT 57.290 202.750 57.570 203.030 ;
        RECT 57.810 202.750 58.090 203.030 ;
        RECT 40.570 201.870 40.850 202.150 ;
        RECT 41.090 201.870 41.370 202.150 ;
        RECT 44.530 201.870 44.810 202.150 ;
        RECT 45.050 201.870 45.330 202.150 ;
        RECT 53.330 201.870 53.610 202.150 ;
        RECT 53.850 201.870 54.130 202.150 ;
        RECT 57.290 201.870 57.570 202.150 ;
        RECT 57.810 201.870 58.090 202.150 ;
        RECT 65.770 203.630 66.050 203.910 ;
        RECT 66.290 203.630 66.570 203.910 ;
        RECT 69.730 203.630 70.010 203.910 ;
        RECT 70.250 203.630 70.530 203.910 ;
        RECT 78.530 203.630 78.810 203.910 ;
        RECT 79.050 203.630 79.330 203.910 ;
        RECT 82.490 203.630 82.770 203.910 ;
        RECT 83.010 203.630 83.290 203.910 ;
        RECT 65.770 202.750 66.050 203.030 ;
        RECT 66.290 202.750 66.570 203.030 ;
        RECT 69.730 202.750 70.010 203.030 ;
        RECT 70.250 202.750 70.530 203.030 ;
        RECT 78.530 202.750 78.810 203.030 ;
        RECT 79.050 202.750 79.330 203.030 ;
        RECT 82.490 202.750 82.770 203.030 ;
        RECT 83.010 202.750 83.290 203.030 ;
        RECT 65.770 201.870 66.050 202.150 ;
        RECT 66.290 201.870 66.570 202.150 ;
        RECT 69.730 201.870 70.010 202.150 ;
        RECT 70.250 201.870 70.530 202.150 ;
        RECT 78.530 201.870 78.810 202.150 ;
        RECT 79.050 201.870 79.330 202.150 ;
        RECT 82.490 201.870 82.770 202.150 ;
        RECT 83.010 201.870 83.290 202.150 ;
        RECT 90.970 203.630 91.250 203.910 ;
        RECT 91.490 203.630 91.770 203.910 ;
        RECT 94.930 203.630 95.210 203.910 ;
        RECT 95.450 203.630 95.730 203.910 ;
        RECT 103.730 203.630 104.010 203.910 ;
        RECT 104.250 203.630 104.530 203.910 ;
        RECT 107.690 203.630 107.970 203.910 ;
        RECT 108.210 203.630 108.490 203.910 ;
        RECT 90.970 202.750 91.250 203.030 ;
        RECT 91.490 202.750 91.770 203.030 ;
        RECT 94.930 202.750 95.210 203.030 ;
        RECT 95.450 202.750 95.730 203.030 ;
        RECT 103.730 202.750 104.010 203.030 ;
        RECT 104.250 202.750 104.530 203.030 ;
        RECT 107.690 202.750 107.970 203.030 ;
        RECT 108.210 202.750 108.490 203.030 ;
        RECT 90.970 201.870 91.250 202.150 ;
        RECT 91.490 201.870 91.770 202.150 ;
        RECT 94.930 201.870 95.210 202.150 ;
        RECT 95.450 201.870 95.730 202.150 ;
        RECT 103.730 201.870 104.010 202.150 ;
        RECT 104.250 201.870 104.530 202.150 ;
        RECT 107.690 201.870 107.970 202.150 ;
        RECT 108.210 201.870 108.490 202.150 ;
        RECT 116.170 203.630 116.450 203.910 ;
        RECT 116.690 203.630 116.970 203.910 ;
        RECT 120.130 203.630 120.410 203.910 ;
        RECT 120.650 203.630 120.930 203.910 ;
        RECT 116.170 202.750 116.450 203.030 ;
        RECT 116.690 202.750 116.970 203.030 ;
        RECT 120.130 202.750 120.410 203.030 ;
        RECT 120.650 202.750 120.930 203.030 ;
        RECT 116.170 201.870 116.450 202.150 ;
        RECT 116.690 201.870 116.970 202.150 ;
        RECT 120.130 201.870 120.410 202.150 ;
        RECT 120.650 201.870 120.930 202.150 ;
        RECT 15.370 199.650 15.650 199.930 ;
        RECT 15.890 199.650 16.170 199.930 ;
        RECT 15.370 199.130 15.650 199.410 ;
        RECT 15.890 199.130 16.170 199.410 ;
        RECT 32.090 199.650 32.370 199.930 ;
        RECT 32.610 199.650 32.890 199.930 ;
        RECT 32.090 199.130 32.370 199.410 ;
        RECT 32.610 199.130 32.890 199.410 ;
        RECT 40.570 199.650 40.850 199.930 ;
        RECT 41.090 199.650 41.370 199.930 ;
        RECT 40.570 199.130 40.850 199.410 ;
        RECT 41.090 199.130 41.370 199.410 ;
        RECT 57.290 199.650 57.570 199.930 ;
        RECT 57.810 199.650 58.090 199.930 ;
        RECT 57.290 199.130 57.570 199.410 ;
        RECT 57.810 199.130 58.090 199.410 ;
        RECT 65.770 199.650 66.050 199.930 ;
        RECT 66.290 199.650 66.570 199.930 ;
        RECT 65.770 199.130 66.050 199.410 ;
        RECT 66.290 199.130 66.570 199.410 ;
        RECT 82.490 199.650 82.770 199.930 ;
        RECT 83.010 199.650 83.290 199.930 ;
        RECT 82.490 199.130 82.770 199.410 ;
        RECT 83.010 199.130 83.290 199.410 ;
        RECT 90.970 199.650 91.250 199.930 ;
        RECT 91.490 199.650 91.770 199.930 ;
        RECT 90.970 199.130 91.250 199.410 ;
        RECT 91.490 199.130 91.770 199.410 ;
        RECT 107.690 199.650 107.970 199.930 ;
        RECT 108.210 199.650 108.490 199.930 ;
        RECT 111.830 199.830 112.170 200.170 ;
        RECT 107.690 199.130 107.970 199.410 ;
        RECT 108.210 199.130 108.490 199.410 ;
        RECT 116.170 199.650 116.450 199.930 ;
        RECT 116.690 199.650 116.970 199.930 ;
        RECT 116.170 199.130 116.450 199.410 ;
        RECT 116.690 199.130 116.970 199.410 ;
        RECT 19.330 198.210 19.610 198.490 ;
        RECT 19.850 198.210 20.130 198.490 ;
        RECT 19.330 197.690 19.610 197.970 ;
        RECT 19.850 197.690 20.130 197.970 ;
        RECT 22.110 198.210 22.390 198.490 ;
        RECT 22.630 198.210 22.910 198.490 ;
        RECT 22.110 197.690 22.390 197.970 ;
        RECT 22.630 197.690 22.910 197.970 ;
        RECT 25.150 198.210 25.430 198.490 ;
        RECT 25.670 198.210 25.950 198.490 ;
        RECT 25.150 197.690 25.430 197.970 ;
        RECT 25.670 197.690 25.950 197.970 ;
        RECT 28.130 198.210 28.410 198.490 ;
        RECT 28.650 198.210 28.930 198.490 ;
        RECT 28.130 197.690 28.410 197.970 ;
        RECT 28.650 197.690 28.930 197.970 ;
        RECT 44.530 198.210 44.810 198.490 ;
        RECT 45.050 198.210 45.330 198.490 ;
        RECT 44.530 197.690 44.810 197.970 ;
        RECT 45.050 197.690 45.330 197.970 ;
        RECT 47.310 198.210 47.590 198.490 ;
        RECT 47.830 198.210 48.110 198.490 ;
        RECT 47.310 197.690 47.590 197.970 ;
        RECT 47.830 197.690 48.110 197.970 ;
        RECT 50.350 198.210 50.630 198.490 ;
        RECT 50.870 198.210 51.150 198.490 ;
        RECT 50.350 197.690 50.630 197.970 ;
        RECT 50.870 197.690 51.150 197.970 ;
        RECT 53.330 198.210 53.610 198.490 ;
        RECT 53.850 198.210 54.130 198.490 ;
        RECT 53.330 197.690 53.610 197.970 ;
        RECT 53.850 197.690 54.130 197.970 ;
        RECT 69.730 198.210 70.010 198.490 ;
        RECT 70.250 198.210 70.530 198.490 ;
        RECT 69.730 197.690 70.010 197.970 ;
        RECT 70.250 197.690 70.530 197.970 ;
        RECT 72.510 198.210 72.790 198.490 ;
        RECT 73.030 198.210 73.310 198.490 ;
        RECT 72.510 197.690 72.790 197.970 ;
        RECT 73.030 197.690 73.310 197.970 ;
        RECT 75.550 198.210 75.830 198.490 ;
        RECT 76.070 198.210 76.350 198.490 ;
        RECT 75.550 197.690 75.830 197.970 ;
        RECT 76.070 197.690 76.350 197.970 ;
        RECT 78.530 198.210 78.810 198.490 ;
        RECT 79.050 198.210 79.330 198.490 ;
        RECT 78.530 197.690 78.810 197.970 ;
        RECT 79.050 197.690 79.330 197.970 ;
        RECT 94.930 198.210 95.210 198.490 ;
        RECT 95.450 198.210 95.730 198.490 ;
        RECT 94.930 197.690 95.210 197.970 ;
        RECT 95.450 197.690 95.730 197.970 ;
        RECT 97.710 198.210 97.990 198.490 ;
        RECT 98.230 198.210 98.510 198.490 ;
        RECT 97.710 197.690 97.990 197.970 ;
        RECT 98.230 197.690 98.510 197.970 ;
        RECT 100.750 198.210 101.030 198.490 ;
        RECT 101.270 198.210 101.550 198.490 ;
        RECT 100.750 197.690 101.030 197.970 ;
        RECT 101.270 197.690 101.550 197.970 ;
        RECT 103.730 198.210 104.010 198.490 ;
        RECT 104.250 198.210 104.530 198.490 ;
        RECT 103.730 197.690 104.010 197.970 ;
        RECT 104.250 197.690 104.530 197.970 ;
        RECT 120.130 198.210 120.410 198.490 ;
        RECT 120.650 198.210 120.930 198.490 ;
        RECT 120.130 197.690 120.410 197.970 ;
        RECT 120.650 197.690 120.930 197.970 ;
        RECT 19.230 194.610 19.510 194.890 ;
        RECT 19.750 194.610 20.030 194.890 ;
        RECT 19.230 194.090 19.510 194.370 ;
        RECT 19.750 194.090 20.030 194.370 ;
        RECT 28.030 194.610 28.310 194.890 ;
        RECT 28.550 194.610 28.830 194.890 ;
        RECT 28.030 194.090 28.310 194.370 ;
        RECT 28.550 194.090 28.830 194.370 ;
        RECT 44.430 194.610 44.710 194.890 ;
        RECT 44.950 194.610 45.230 194.890 ;
        RECT 44.430 194.090 44.710 194.370 ;
        RECT 44.950 194.090 45.230 194.370 ;
        RECT 53.230 194.610 53.510 194.890 ;
        RECT 53.750 194.610 54.030 194.890 ;
        RECT 53.230 194.090 53.510 194.370 ;
        RECT 53.750 194.090 54.030 194.370 ;
        RECT 69.630 194.610 69.910 194.890 ;
        RECT 70.150 194.610 70.430 194.890 ;
        RECT 69.630 194.090 69.910 194.370 ;
        RECT 70.150 194.090 70.430 194.370 ;
        RECT 78.430 194.610 78.710 194.890 ;
        RECT 78.950 194.610 79.230 194.890 ;
        RECT 78.430 194.090 78.710 194.370 ;
        RECT 78.950 194.090 79.230 194.370 ;
        RECT 94.830 194.610 95.110 194.890 ;
        RECT 95.350 194.610 95.630 194.890 ;
        RECT 94.830 194.090 95.110 194.370 ;
        RECT 95.350 194.090 95.630 194.370 ;
        RECT 103.630 194.610 103.910 194.890 ;
        RECT 104.150 194.610 104.430 194.890 ;
        RECT 103.630 194.090 103.910 194.370 ;
        RECT 104.150 194.090 104.430 194.370 ;
        RECT 120.030 194.610 120.310 194.890 ;
        RECT 120.550 194.610 120.830 194.890 ;
        RECT 120.030 194.090 120.310 194.370 ;
        RECT 120.550 194.090 120.830 194.370 ;
        RECT 15.270 191.010 15.550 191.290 ;
        RECT 15.790 191.010 16.070 191.290 ;
        RECT 15.270 190.490 15.550 190.770 ;
        RECT 15.790 190.490 16.070 190.770 ;
        RECT 31.990 191.010 32.270 191.290 ;
        RECT 32.510 191.010 32.790 191.290 ;
        RECT 31.990 190.490 32.270 190.770 ;
        RECT 32.510 190.490 32.790 190.770 ;
        RECT 40.470 191.010 40.750 191.290 ;
        RECT 40.990 191.010 41.270 191.290 ;
        RECT 40.470 190.490 40.750 190.770 ;
        RECT 40.990 190.490 41.270 190.770 ;
        RECT 57.190 191.010 57.470 191.290 ;
        RECT 57.710 191.010 57.990 191.290 ;
        RECT 57.190 190.490 57.470 190.770 ;
        RECT 57.710 190.490 57.990 190.770 ;
        RECT 65.670 191.010 65.950 191.290 ;
        RECT 66.190 191.010 66.470 191.290 ;
        RECT 65.670 190.490 65.950 190.770 ;
        RECT 66.190 190.490 66.470 190.770 ;
        RECT 82.390 191.010 82.670 191.290 ;
        RECT 82.910 191.010 83.190 191.290 ;
        RECT 82.390 190.490 82.670 190.770 ;
        RECT 82.910 190.490 83.190 190.770 ;
        RECT 90.870 191.010 91.150 191.290 ;
        RECT 91.390 191.010 91.670 191.290 ;
        RECT 90.870 190.490 91.150 190.770 ;
        RECT 91.390 190.490 91.670 190.770 ;
        RECT 107.590 191.010 107.870 191.290 ;
        RECT 108.110 191.010 108.390 191.290 ;
        RECT 107.590 190.490 107.870 190.770 ;
        RECT 108.110 190.490 108.390 190.770 ;
        RECT 116.070 191.010 116.350 191.290 ;
        RECT 116.590 191.010 116.870 191.290 ;
        RECT 116.070 190.490 116.350 190.770 ;
        RECT 116.590 190.490 116.870 190.770 ;
        RECT 15.270 187.170 15.550 187.450 ;
        RECT 15.790 187.170 16.070 187.450 ;
        RECT 19.230 187.170 19.510 187.450 ;
        RECT 19.750 187.170 20.030 187.450 ;
        RECT 28.030 187.170 28.310 187.450 ;
        RECT 28.550 187.170 28.830 187.450 ;
        RECT 31.990 187.170 32.270 187.450 ;
        RECT 32.510 187.170 32.790 187.450 ;
        RECT 40.470 187.170 40.750 187.450 ;
        RECT 40.990 187.170 41.270 187.450 ;
        RECT 44.430 187.170 44.710 187.450 ;
        RECT 44.950 187.170 45.230 187.450 ;
        RECT 53.230 187.170 53.510 187.450 ;
        RECT 53.750 187.170 54.030 187.450 ;
        RECT 57.190 187.170 57.470 187.450 ;
        RECT 57.710 187.170 57.990 187.450 ;
        RECT 65.670 187.170 65.950 187.450 ;
        RECT 66.190 187.170 66.470 187.450 ;
        RECT 69.630 187.170 69.910 187.450 ;
        RECT 70.150 187.170 70.430 187.450 ;
        RECT 78.430 187.170 78.710 187.450 ;
        RECT 78.950 187.170 79.230 187.450 ;
        RECT 82.390 187.170 82.670 187.450 ;
        RECT 82.910 187.170 83.190 187.450 ;
        RECT 90.870 187.170 91.150 187.450 ;
        RECT 91.390 187.170 91.670 187.450 ;
        RECT 94.830 187.170 95.110 187.450 ;
        RECT 95.350 187.170 95.630 187.450 ;
        RECT 103.630 187.170 103.910 187.450 ;
        RECT 104.150 187.170 104.430 187.450 ;
        RECT 107.590 187.170 107.870 187.450 ;
        RECT 108.110 187.170 108.390 187.450 ;
        RECT 15.270 186.290 15.550 186.570 ;
        RECT 15.790 186.290 16.070 186.570 ;
        RECT 19.230 186.290 19.510 186.570 ;
        RECT 19.750 186.290 20.030 186.570 ;
        RECT 28.030 186.290 28.310 186.570 ;
        RECT 28.550 186.290 28.830 186.570 ;
        RECT 31.990 186.290 32.270 186.570 ;
        RECT 32.510 186.290 32.790 186.570 ;
        RECT 40.470 186.290 40.750 186.570 ;
        RECT 40.990 186.290 41.270 186.570 ;
        RECT 44.430 186.290 44.710 186.570 ;
        RECT 44.950 186.290 45.230 186.570 ;
        RECT 53.230 186.290 53.510 186.570 ;
        RECT 53.750 186.290 54.030 186.570 ;
        RECT 57.190 186.290 57.470 186.570 ;
        RECT 57.710 186.290 57.990 186.570 ;
        RECT 65.670 186.290 65.950 186.570 ;
        RECT 66.190 186.290 66.470 186.570 ;
        RECT 69.630 186.290 69.910 186.570 ;
        RECT 70.150 186.290 70.430 186.570 ;
        RECT 78.430 186.290 78.710 186.570 ;
        RECT 78.950 186.290 79.230 186.570 ;
        RECT 82.390 186.290 82.670 186.570 ;
        RECT 82.910 186.290 83.190 186.570 ;
        RECT 90.870 186.290 91.150 186.570 ;
        RECT 91.390 186.290 91.670 186.570 ;
        RECT 94.830 186.290 95.110 186.570 ;
        RECT 95.350 186.290 95.630 186.570 ;
        RECT 103.630 186.290 103.910 186.570 ;
        RECT 104.150 186.290 104.430 186.570 ;
        RECT 107.590 186.290 107.870 186.570 ;
        RECT 108.110 186.290 108.390 186.570 ;
        RECT 19.230 185.580 19.510 185.860 ;
        RECT 19.750 185.580 20.030 185.860 ;
        RECT 44.430 185.580 44.710 185.860 ;
        RECT 44.950 185.580 45.230 185.860 ;
        RECT 69.630 185.580 69.910 185.860 ;
        RECT 70.150 185.580 70.430 185.860 ;
        RECT 94.830 185.580 95.110 185.860 ;
        RECT 95.350 185.580 95.630 185.860 ;
        RECT 103.470 185.410 103.750 185.690 ;
        RECT 103.990 185.410 104.270 185.690 ;
        RECT 15.270 184.530 15.550 184.810 ;
        RECT 15.790 184.530 16.070 184.810 ;
        RECT 19.230 184.530 19.510 184.810 ;
        RECT 19.750 184.530 20.030 184.810 ;
        RECT 28.030 184.530 28.310 184.810 ;
        RECT 28.550 184.530 28.830 184.810 ;
        RECT 15.270 183.650 15.550 183.930 ;
        RECT 15.790 183.650 16.070 183.930 ;
        RECT 31.990 184.530 32.270 184.810 ;
        RECT 32.510 184.530 32.790 184.810 ;
        RECT 40.470 184.530 40.750 184.810 ;
        RECT 40.990 184.530 41.270 184.810 ;
        RECT 44.430 184.530 44.710 184.810 ;
        RECT 44.950 184.530 45.230 184.810 ;
        RECT 53.230 184.530 53.510 184.810 ;
        RECT 53.750 184.530 54.030 184.810 ;
        RECT 31.990 183.650 32.270 183.930 ;
        RECT 32.510 183.650 32.790 183.930 ;
        RECT 40.470 183.650 40.750 183.930 ;
        RECT 40.990 183.650 41.270 183.930 ;
        RECT 33.990 183.210 34.270 183.490 ;
        RECT 34.510 183.210 34.790 183.490 ;
        RECT 57.190 184.530 57.470 184.810 ;
        RECT 57.710 184.530 57.990 184.810 ;
        RECT 65.670 184.530 65.950 184.810 ;
        RECT 66.190 184.530 66.470 184.810 ;
        RECT 69.630 184.530 69.910 184.810 ;
        RECT 70.150 184.530 70.430 184.810 ;
        RECT 78.430 184.530 78.710 184.810 ;
        RECT 78.950 184.530 79.230 184.810 ;
        RECT 57.190 183.650 57.470 183.930 ;
        RECT 57.710 183.650 57.990 183.930 ;
        RECT 65.670 183.650 65.950 183.930 ;
        RECT 66.190 183.650 66.470 183.930 ;
        RECT 59.190 183.210 59.470 183.490 ;
        RECT 59.710 183.210 59.990 183.490 ;
        RECT 82.390 184.530 82.670 184.810 ;
        RECT 82.910 184.530 83.190 184.810 ;
        RECT 90.870 184.530 91.150 184.810 ;
        RECT 91.390 184.530 91.670 184.810 ;
        RECT 94.830 184.530 95.110 184.810 ;
        RECT 95.350 184.530 95.630 184.810 ;
        RECT 103.630 184.530 103.910 184.810 ;
        RECT 104.150 184.530 104.430 184.810 ;
        RECT 107.590 184.530 107.870 184.810 ;
        RECT 108.110 184.530 108.390 184.810 ;
        RECT 82.390 183.650 82.670 183.930 ;
        RECT 82.910 183.650 83.190 183.930 ;
        RECT 90.870 183.650 91.150 183.930 ;
        RECT 91.390 183.650 91.670 183.930 ;
        RECT 107.590 183.650 107.870 183.930 ;
        RECT 108.110 183.650 108.390 183.930 ;
        RECT 84.390 183.210 84.670 183.490 ;
        RECT 84.910 183.210 85.190 183.490 ;
        RECT 109.590 183.210 109.870 183.490 ;
        RECT 110.110 183.210 110.390 183.490 ;
        RECT 116.070 182.770 116.350 183.050 ;
        RECT 116.590 182.770 116.870 183.050 ;
        RECT 120.030 182.770 120.310 183.050 ;
        RECT 120.550 182.770 120.830 183.050 ;
        RECT 15.270 181.890 15.550 182.170 ;
        RECT 15.790 181.890 16.070 182.170 ;
        RECT 19.230 181.890 19.510 182.170 ;
        RECT 19.750 181.890 20.030 182.170 ;
        RECT 28.030 181.890 28.310 182.170 ;
        RECT 28.550 181.890 28.830 182.170 ;
        RECT 31.990 181.890 32.270 182.170 ;
        RECT 32.510 181.890 32.790 182.170 ;
        RECT 40.470 181.890 40.750 182.170 ;
        RECT 40.990 181.890 41.270 182.170 ;
        RECT 44.430 181.890 44.710 182.170 ;
        RECT 44.950 181.890 45.230 182.170 ;
        RECT 53.230 181.890 53.510 182.170 ;
        RECT 53.750 181.890 54.030 182.170 ;
        RECT 57.190 181.890 57.470 182.170 ;
        RECT 57.710 181.890 57.990 182.170 ;
        RECT 65.670 181.890 65.950 182.170 ;
        RECT 66.190 181.890 66.470 182.170 ;
        RECT 69.630 181.890 69.910 182.170 ;
        RECT 70.150 181.890 70.430 182.170 ;
        RECT 78.430 181.890 78.710 182.170 ;
        RECT 78.950 181.890 79.230 182.170 ;
        RECT 82.390 181.890 82.670 182.170 ;
        RECT 82.910 181.890 83.190 182.170 ;
        RECT 90.870 181.890 91.150 182.170 ;
        RECT 91.390 181.890 91.670 182.170 ;
        RECT 94.830 181.890 95.110 182.170 ;
        RECT 95.350 181.890 95.630 182.170 ;
        RECT 103.630 181.890 103.910 182.170 ;
        RECT 104.150 181.890 104.430 182.170 ;
        RECT 107.590 181.890 107.870 182.170 ;
        RECT 108.110 181.890 108.390 182.170 ;
        RECT 116.070 181.890 116.350 182.170 ;
        RECT 116.590 181.890 116.870 182.170 ;
        RECT 120.030 181.890 120.310 182.170 ;
        RECT 120.550 181.890 120.830 182.170 ;
        RECT 113.910 180.740 114.190 181.020 ;
        RECT 114.430 180.740 114.710 181.020 ;
        RECT 15.270 180.130 15.550 180.410 ;
        RECT 15.790 180.130 16.070 180.410 ;
        RECT 19.230 180.130 19.510 180.410 ;
        RECT 19.750 180.130 20.030 180.410 ;
        RECT 28.030 180.130 28.310 180.410 ;
        RECT 28.550 180.130 28.830 180.410 ;
        RECT 31.990 180.130 32.270 180.410 ;
        RECT 32.510 180.130 32.790 180.410 ;
        RECT 40.470 180.130 40.750 180.410 ;
        RECT 40.990 180.130 41.270 180.410 ;
        RECT 44.430 180.130 44.710 180.410 ;
        RECT 44.950 180.130 45.230 180.410 ;
        RECT 53.230 180.130 53.510 180.410 ;
        RECT 53.750 180.130 54.030 180.410 ;
        RECT 57.190 180.130 57.470 180.410 ;
        RECT 57.710 180.130 57.990 180.410 ;
        RECT 65.670 180.130 65.950 180.410 ;
        RECT 66.190 180.130 66.470 180.410 ;
        RECT 69.630 180.130 69.910 180.410 ;
        RECT 70.150 180.130 70.430 180.410 ;
        RECT 78.430 180.130 78.710 180.410 ;
        RECT 78.950 180.130 79.230 180.410 ;
        RECT 82.390 180.130 82.670 180.410 ;
        RECT 82.910 180.130 83.190 180.410 ;
        RECT 90.870 180.130 91.150 180.410 ;
        RECT 91.390 180.130 91.670 180.410 ;
        RECT 94.830 180.130 95.110 180.410 ;
        RECT 95.350 180.130 95.630 180.410 ;
        RECT 103.630 180.130 103.910 180.410 ;
        RECT 104.150 180.130 104.430 180.410 ;
        RECT 107.590 180.130 107.870 180.410 ;
        RECT 108.110 180.130 108.390 180.410 ;
        RECT 116.070 180.130 116.350 180.410 ;
        RECT 116.590 180.130 116.870 180.410 ;
        RECT 120.030 180.130 120.310 180.410 ;
        RECT 120.550 180.130 120.830 180.410 ;
        RECT 19.230 179.250 19.510 179.530 ;
        RECT 19.750 179.250 20.030 179.530 ;
        RECT 28.030 179.250 28.310 179.530 ;
        RECT 28.550 179.250 28.830 179.530 ;
        RECT 44.430 179.250 44.710 179.530 ;
        RECT 44.950 179.250 45.230 179.530 ;
        RECT 53.230 179.250 53.510 179.530 ;
        RECT 53.750 179.250 54.030 179.530 ;
        RECT 69.630 179.250 69.910 179.530 ;
        RECT 70.150 179.250 70.430 179.530 ;
        RECT 78.430 179.250 78.710 179.530 ;
        RECT 78.950 179.250 79.230 179.530 ;
        RECT 94.830 179.250 95.110 179.530 ;
        RECT 95.350 179.250 95.630 179.530 ;
        RECT 103.630 179.250 103.910 179.530 ;
        RECT 104.150 179.250 104.430 179.530 ;
        RECT 116.070 179.250 116.350 179.530 ;
        RECT 116.590 179.250 116.870 179.530 ;
        RECT 15.270 177.490 15.550 177.770 ;
        RECT 15.790 177.490 16.070 177.770 ;
        RECT 19.230 177.490 19.510 177.770 ;
        RECT 19.750 177.490 20.030 177.770 ;
        RECT 28.030 177.490 28.310 177.770 ;
        RECT 28.550 177.490 28.830 177.770 ;
        RECT 31.990 177.490 32.270 177.770 ;
        RECT 32.510 177.490 32.790 177.770 ;
        RECT 15.270 176.610 15.550 176.890 ;
        RECT 15.790 176.610 16.070 176.890 ;
        RECT 31.830 176.610 32.110 176.890 ;
        RECT 32.350 176.610 32.630 176.890 ;
        RECT 15.270 175.730 15.550 176.010 ;
        RECT 15.790 175.730 16.070 176.010 ;
        RECT 19.230 175.730 19.510 176.010 ;
        RECT 19.750 175.730 20.030 176.010 ;
        RECT 28.030 175.730 28.310 176.010 ;
        RECT 28.550 175.730 28.830 176.010 ;
        RECT 31.990 175.730 32.270 176.010 ;
        RECT 32.510 175.730 32.790 176.010 ;
        RECT 15.270 173.970 15.550 174.250 ;
        RECT 15.790 173.970 16.070 174.250 ;
        RECT 19.230 173.970 19.510 174.250 ;
        RECT 19.750 173.970 20.030 174.250 ;
        RECT 15.270 171.330 15.550 171.610 ;
        RECT 15.790 171.330 16.070 171.610 ;
        RECT 19.230 171.330 19.510 171.610 ;
        RECT 19.750 171.330 20.030 171.610 ;
        RECT 13.110 170.890 13.390 171.170 ;
        RECT 13.630 170.890 13.910 171.170 ;
        RECT 15.270 169.570 15.550 169.850 ;
        RECT 15.790 169.570 16.070 169.850 ;
        RECT 15.270 168.690 15.550 168.970 ;
        RECT 15.790 168.690 16.070 168.970 ;
        RECT 19.230 168.690 19.510 168.970 ;
        RECT 19.750 168.690 20.030 168.970 ;
        RECT 15.270 166.930 15.550 167.210 ;
        RECT 15.790 166.930 16.070 167.210 ;
        RECT 19.230 166.930 19.510 167.210 ;
        RECT 19.750 166.930 20.030 167.210 ;
        RECT 18.190 166.310 18.470 166.590 ;
        RECT 18.190 165.790 18.470 166.070 ;
        RECT 15.270 165.170 15.550 165.450 ;
        RECT 15.790 165.170 16.070 165.450 ;
        RECT 19.230 165.170 19.510 165.450 ;
        RECT 19.750 165.170 20.030 165.450 ;
        RECT 15.270 164.290 15.550 164.570 ;
        RECT 15.790 164.290 16.070 164.570 ;
        RECT 19.230 164.290 19.510 164.570 ;
        RECT 19.750 164.290 20.030 164.570 ;
        RECT 15.270 162.530 15.550 162.810 ;
        RECT 15.790 162.530 16.070 162.810 ;
        RECT 19.230 162.530 19.510 162.810 ;
        RECT 19.750 162.530 20.030 162.810 ;
        RECT 17.405 161.910 17.685 162.190 ;
        RECT 17.405 161.390 17.685 161.670 ;
        RECT 13.270 156.810 13.550 157.090 ;
        RECT 13.790 156.810 14.070 157.090 ;
        RECT 13.110 150.650 13.390 150.930 ;
        RECT 13.630 150.650 13.910 150.930 ;
        RECT 13.110 148.890 13.390 149.170 ;
        RECT 13.630 148.890 13.910 149.170 ;
        RECT 15.270 160.770 15.550 161.050 ;
        RECT 15.790 160.770 16.070 161.050 ;
        RECT 19.230 160.770 19.510 161.050 ;
        RECT 19.750 160.770 20.030 161.050 ;
        RECT 15.270 159.890 15.550 160.170 ;
        RECT 15.790 159.890 16.070 160.170 ;
        RECT 19.230 159.890 19.510 160.170 ;
        RECT 19.750 159.890 20.030 160.170 ;
        RECT 15.270 158.130 15.550 158.410 ;
        RECT 15.790 158.130 16.070 158.410 ;
        RECT 19.230 158.130 19.510 158.410 ;
        RECT 19.750 158.130 20.030 158.410 ;
        RECT 16.690 157.510 16.970 157.790 ;
        RECT 16.690 156.990 16.970 157.270 ;
        RECT 15.270 156.370 15.550 156.650 ;
        RECT 15.790 156.370 16.070 156.650 ;
        RECT 19.230 156.370 19.510 156.650 ;
        RECT 19.750 156.370 20.030 156.650 ;
        RECT 15.270 155.490 15.550 155.770 ;
        RECT 15.790 155.490 16.070 155.770 ;
        RECT 19.230 155.490 19.510 155.770 ;
        RECT 19.750 155.490 20.030 155.770 ;
        RECT 15.270 153.730 15.550 154.010 ;
        RECT 15.790 153.730 16.070 154.010 ;
        RECT 19.230 153.730 19.510 154.010 ;
        RECT 19.750 153.730 20.030 154.010 ;
        RECT 15.270 151.970 15.550 152.250 ;
        RECT 15.790 151.970 16.070 152.250 ;
        RECT 19.230 151.970 19.510 152.250 ;
        RECT 19.750 151.970 20.030 152.250 ;
        RECT 21.390 150.650 21.670 150.930 ;
        RECT 21.910 150.650 22.190 150.930 ;
        RECT 15.270 148.450 15.550 148.730 ;
        RECT 15.790 148.450 16.070 148.730 ;
        RECT 19.230 148.450 19.510 148.730 ;
        RECT 19.750 148.450 20.030 148.730 ;
        RECT 13.270 145.370 13.550 145.650 ;
        RECT 13.790 145.370 14.070 145.650 ;
        RECT 15.270 144.930 15.550 145.210 ;
        RECT 15.790 144.930 16.070 145.210 ;
        RECT 19.230 144.930 19.510 145.210 ;
        RECT 19.750 144.930 20.030 145.210 ;
        RECT 15.270 143.170 15.550 143.450 ;
        RECT 15.790 143.170 16.070 143.450 ;
        RECT 19.230 143.170 19.510 143.450 ;
        RECT 19.750 143.170 20.030 143.450 ;
        RECT 19.230 142.290 19.510 142.570 ;
        RECT 19.750 142.290 20.030 142.570 ;
        RECT 15.270 141.410 15.550 141.690 ;
        RECT 15.790 141.410 16.070 141.690 ;
        RECT 15.270 140.530 15.550 140.810 ;
        RECT 15.790 140.530 16.070 140.810 ;
        RECT 15.270 137.890 15.550 138.170 ;
        RECT 15.790 137.890 16.070 138.170 ;
        RECT 19.390 137.890 19.670 138.170 ;
        RECT 19.910 137.890 20.190 138.170 ;
        RECT 28.030 173.970 28.310 174.250 ;
        RECT 28.550 173.970 28.830 174.250 ;
        RECT 31.990 173.970 32.270 174.250 ;
        RECT 32.510 173.970 32.790 174.250 ;
        RECT 40.470 177.490 40.750 177.770 ;
        RECT 40.990 177.490 41.270 177.770 ;
        RECT 44.430 177.490 44.710 177.770 ;
        RECT 44.950 177.490 45.230 177.770 ;
        RECT 53.230 177.490 53.510 177.770 ;
        RECT 53.750 177.490 54.030 177.770 ;
        RECT 57.190 177.490 57.470 177.770 ;
        RECT 57.710 177.490 57.990 177.770 ;
        RECT 40.470 176.610 40.750 176.890 ;
        RECT 40.990 176.610 41.270 176.890 ;
        RECT 57.030 176.610 57.310 176.890 ;
        RECT 57.550 176.610 57.830 176.890 ;
        RECT 40.470 175.730 40.750 176.010 ;
        RECT 40.990 175.730 41.270 176.010 ;
        RECT 44.430 175.730 44.710 176.010 ;
        RECT 44.950 175.730 45.230 176.010 ;
        RECT 53.230 175.730 53.510 176.010 ;
        RECT 53.750 175.730 54.030 176.010 ;
        RECT 57.190 175.730 57.470 176.010 ;
        RECT 57.710 175.730 57.990 176.010 ;
        RECT 40.470 173.970 40.750 174.250 ;
        RECT 40.990 173.970 41.270 174.250 ;
        RECT 44.430 173.970 44.710 174.250 ;
        RECT 44.950 173.970 45.230 174.250 ;
        RECT 28.030 171.330 28.310 171.610 ;
        RECT 28.550 171.330 28.830 171.610 ;
        RECT 31.990 171.330 32.270 171.610 ;
        RECT 32.510 171.330 32.790 171.610 ;
        RECT 40.470 171.330 40.750 171.610 ;
        RECT 40.990 171.330 41.270 171.610 ;
        RECT 44.430 171.330 44.710 171.610 ;
        RECT 44.950 171.330 45.230 171.610 ;
        RECT 33.990 170.890 34.270 171.170 ;
        RECT 34.510 170.890 34.790 171.170 ;
        RECT 38.310 170.890 38.590 171.170 ;
        RECT 38.830 170.890 39.110 171.170 ;
        RECT 31.990 169.570 32.270 169.850 ;
        RECT 32.510 169.570 32.790 169.850 ;
        RECT 40.470 169.570 40.750 169.850 ;
        RECT 40.990 169.570 41.270 169.850 ;
        RECT 28.030 168.690 28.310 168.970 ;
        RECT 28.550 168.690 28.830 168.970 ;
        RECT 31.990 168.690 32.270 168.970 ;
        RECT 32.510 168.690 32.790 168.970 ;
        RECT 40.470 168.690 40.750 168.970 ;
        RECT 40.990 168.690 41.270 168.970 ;
        RECT 44.430 168.690 44.710 168.970 ;
        RECT 44.950 168.690 45.230 168.970 ;
        RECT 28.030 166.930 28.310 167.210 ;
        RECT 28.550 166.930 28.830 167.210 ;
        RECT 31.990 166.930 32.270 167.210 ;
        RECT 32.510 166.930 32.790 167.210 ;
        RECT 40.470 166.930 40.750 167.210 ;
        RECT 40.990 166.930 41.270 167.210 ;
        RECT 44.430 166.930 44.710 167.210 ;
        RECT 44.950 166.930 45.230 167.210 ;
        RECT 29.590 166.310 29.870 166.590 ;
        RECT 29.590 165.790 29.870 166.070 ;
        RECT 43.390 166.310 43.670 166.590 ;
        RECT 43.390 165.790 43.670 166.070 ;
        RECT 28.030 165.170 28.310 165.450 ;
        RECT 28.550 165.170 28.830 165.450 ;
        RECT 31.990 165.170 32.270 165.450 ;
        RECT 32.510 165.170 32.790 165.450 ;
        RECT 40.470 165.170 40.750 165.450 ;
        RECT 40.990 165.170 41.270 165.450 ;
        RECT 44.430 165.170 44.710 165.450 ;
        RECT 44.950 165.170 45.230 165.450 ;
        RECT 28.030 164.290 28.310 164.570 ;
        RECT 28.550 164.290 28.830 164.570 ;
        RECT 31.990 164.290 32.270 164.570 ;
        RECT 32.510 164.290 32.790 164.570 ;
        RECT 40.470 164.290 40.750 164.570 ;
        RECT 40.990 164.290 41.270 164.570 ;
        RECT 44.430 164.290 44.710 164.570 ;
        RECT 44.950 164.290 45.230 164.570 ;
        RECT 28.030 162.530 28.310 162.810 ;
        RECT 28.550 162.530 28.830 162.810 ;
        RECT 31.990 162.530 32.270 162.810 ;
        RECT 32.510 162.530 32.790 162.810 ;
        RECT 40.470 162.530 40.750 162.810 ;
        RECT 40.990 162.530 41.270 162.810 ;
        RECT 44.430 162.530 44.710 162.810 ;
        RECT 44.950 162.530 45.230 162.810 ;
        RECT 30.375 161.910 30.655 162.190 ;
        RECT 30.375 161.390 30.655 161.670 ;
        RECT 42.605 161.910 42.885 162.190 ;
        RECT 42.605 161.390 42.885 161.670 ;
        RECT 28.030 160.770 28.310 161.050 ;
        RECT 28.550 160.770 28.830 161.050 ;
        RECT 31.990 160.770 32.270 161.050 ;
        RECT 32.510 160.770 32.790 161.050 ;
        RECT 28.030 159.890 28.310 160.170 ;
        RECT 28.550 159.890 28.830 160.170 ;
        RECT 31.990 159.890 32.270 160.170 ;
        RECT 32.510 159.890 32.790 160.170 ;
        RECT 28.030 158.130 28.310 158.410 ;
        RECT 28.550 158.130 28.830 158.410 ;
        RECT 31.990 158.130 32.270 158.410 ;
        RECT 32.510 158.130 32.790 158.410 ;
        RECT 31.090 157.510 31.370 157.790 ;
        RECT 31.090 156.990 31.370 157.270 ;
        RECT 28.030 156.370 28.310 156.650 ;
        RECT 28.550 156.370 28.830 156.650 ;
        RECT 31.990 156.370 32.270 156.650 ;
        RECT 32.510 156.370 32.790 156.650 ;
        RECT 28.030 155.490 28.310 155.770 ;
        RECT 28.550 155.490 28.830 155.770 ;
        RECT 31.990 155.490 32.270 155.770 ;
        RECT 32.510 155.490 32.790 155.770 ;
        RECT 28.030 153.730 28.310 154.010 ;
        RECT 28.550 153.730 28.830 154.010 ;
        RECT 31.990 153.730 32.270 154.010 ;
        RECT 32.510 153.730 32.790 154.010 ;
        RECT 28.030 151.970 28.310 152.250 ;
        RECT 28.550 151.970 28.830 152.250 ;
        RECT 31.990 151.970 32.270 152.250 ;
        RECT 32.510 151.970 32.790 152.250 ;
        RECT 25.710 150.650 25.990 150.930 ;
        RECT 26.230 150.650 26.510 150.930 ;
        RECT 28.030 148.450 28.310 148.730 ;
        RECT 28.550 148.450 28.830 148.730 ;
        RECT 31.990 148.450 32.270 148.730 ;
        RECT 32.510 148.450 32.790 148.730 ;
        RECT 33.990 156.810 34.270 157.090 ;
        RECT 34.510 156.810 34.790 157.090 ;
        RECT 38.470 156.810 38.750 157.090 ;
        RECT 38.990 156.810 39.270 157.090 ;
        RECT 33.990 148.890 34.270 149.170 ;
        RECT 34.510 148.890 34.790 149.170 ;
        RECT 33.990 145.370 34.270 145.650 ;
        RECT 34.510 145.370 34.790 145.650 ;
        RECT 28.030 144.930 28.310 145.210 ;
        RECT 28.550 144.930 28.830 145.210 ;
        RECT 31.990 144.930 32.270 145.210 ;
        RECT 32.510 144.930 32.790 145.210 ;
        RECT 28.030 143.170 28.310 143.450 ;
        RECT 28.550 143.170 28.830 143.450 ;
        RECT 31.990 143.170 32.270 143.450 ;
        RECT 32.510 143.170 32.790 143.450 ;
        RECT 28.030 142.290 28.310 142.570 ;
        RECT 28.550 142.290 28.830 142.570 ;
        RECT 31.990 141.410 32.270 141.690 ;
        RECT 32.510 141.410 32.790 141.690 ;
        RECT 31.990 140.530 32.270 140.810 ;
        RECT 32.510 140.530 32.790 140.810 ;
        RECT 27.870 137.890 28.150 138.170 ;
        RECT 28.390 137.890 28.670 138.170 ;
        RECT 31.990 137.890 32.270 138.170 ;
        RECT 32.510 137.890 32.790 138.170 ;
        RECT 19.230 137.010 19.510 137.290 ;
        RECT 19.750 137.010 20.030 137.290 ;
        RECT 28.030 137.010 28.310 137.290 ;
        RECT 28.550 137.010 28.830 137.290 ;
        RECT 13.270 136.570 13.550 136.850 ;
        RECT 13.790 136.570 14.070 136.850 ;
        RECT 33.990 136.570 34.270 136.850 ;
        RECT 34.510 136.570 34.790 136.850 ;
        RECT 38.310 148.890 38.590 149.170 ;
        RECT 38.830 148.890 39.110 149.170 ;
        RECT 40.470 160.770 40.750 161.050 ;
        RECT 40.990 160.770 41.270 161.050 ;
        RECT 44.430 160.770 44.710 161.050 ;
        RECT 44.950 160.770 45.230 161.050 ;
        RECT 40.470 159.890 40.750 160.170 ;
        RECT 40.990 159.890 41.270 160.170 ;
        RECT 44.430 159.890 44.710 160.170 ;
        RECT 44.950 159.890 45.230 160.170 ;
        RECT 40.470 158.130 40.750 158.410 ;
        RECT 40.990 158.130 41.270 158.410 ;
        RECT 44.430 158.130 44.710 158.410 ;
        RECT 44.950 158.130 45.230 158.410 ;
        RECT 41.890 157.510 42.170 157.790 ;
        RECT 41.890 156.990 42.170 157.270 ;
        RECT 40.470 156.370 40.750 156.650 ;
        RECT 40.990 156.370 41.270 156.650 ;
        RECT 44.430 156.370 44.710 156.650 ;
        RECT 44.950 156.370 45.230 156.650 ;
        RECT 40.470 155.490 40.750 155.770 ;
        RECT 40.990 155.490 41.270 155.770 ;
        RECT 44.430 155.490 44.710 155.770 ;
        RECT 44.950 155.490 45.230 155.770 ;
        RECT 40.470 153.730 40.750 154.010 ;
        RECT 40.990 153.730 41.270 154.010 ;
        RECT 44.430 153.730 44.710 154.010 ;
        RECT 44.950 153.730 45.230 154.010 ;
        RECT 40.470 151.970 40.750 152.250 ;
        RECT 40.990 151.970 41.270 152.250 ;
        RECT 44.430 151.970 44.710 152.250 ;
        RECT 44.950 151.970 45.230 152.250 ;
        RECT 46.590 150.650 46.870 150.930 ;
        RECT 47.110 150.650 47.390 150.930 ;
        RECT 40.470 148.450 40.750 148.730 ;
        RECT 40.990 148.450 41.270 148.730 ;
        RECT 44.430 148.450 44.710 148.730 ;
        RECT 44.950 148.450 45.230 148.730 ;
        RECT 38.470 145.370 38.750 145.650 ;
        RECT 38.990 145.370 39.270 145.650 ;
        RECT 40.470 144.930 40.750 145.210 ;
        RECT 40.990 144.930 41.270 145.210 ;
        RECT 44.430 144.930 44.710 145.210 ;
        RECT 44.950 144.930 45.230 145.210 ;
        RECT 40.470 143.170 40.750 143.450 ;
        RECT 40.990 143.170 41.270 143.450 ;
        RECT 44.430 143.170 44.710 143.450 ;
        RECT 44.950 143.170 45.230 143.450 ;
        RECT 44.430 142.290 44.710 142.570 ;
        RECT 44.950 142.290 45.230 142.570 ;
        RECT 40.470 141.410 40.750 141.690 ;
        RECT 40.990 141.410 41.270 141.690 ;
        RECT 40.470 140.530 40.750 140.810 ;
        RECT 40.990 140.530 41.270 140.810 ;
        RECT 40.470 137.890 40.750 138.170 ;
        RECT 40.990 137.890 41.270 138.170 ;
        RECT 44.590 137.890 44.870 138.170 ;
        RECT 45.110 137.890 45.390 138.170 ;
        RECT 53.230 173.970 53.510 174.250 ;
        RECT 53.750 173.970 54.030 174.250 ;
        RECT 57.190 173.970 57.470 174.250 ;
        RECT 57.710 173.970 57.990 174.250 ;
        RECT 65.670 177.490 65.950 177.770 ;
        RECT 66.190 177.490 66.470 177.770 ;
        RECT 69.630 177.490 69.910 177.770 ;
        RECT 70.150 177.490 70.430 177.770 ;
        RECT 78.430 177.490 78.710 177.770 ;
        RECT 78.950 177.490 79.230 177.770 ;
        RECT 82.390 177.490 82.670 177.770 ;
        RECT 82.910 177.490 83.190 177.770 ;
        RECT 65.670 176.610 65.950 176.890 ;
        RECT 66.190 176.610 66.470 176.890 ;
        RECT 82.230 176.610 82.510 176.890 ;
        RECT 82.750 176.610 83.030 176.890 ;
        RECT 65.670 175.730 65.950 176.010 ;
        RECT 66.190 175.730 66.470 176.010 ;
        RECT 69.630 175.730 69.910 176.010 ;
        RECT 70.150 175.730 70.430 176.010 ;
        RECT 78.430 175.730 78.710 176.010 ;
        RECT 78.950 175.730 79.230 176.010 ;
        RECT 82.390 175.730 82.670 176.010 ;
        RECT 82.910 175.730 83.190 176.010 ;
        RECT 65.670 173.970 65.950 174.250 ;
        RECT 66.190 173.970 66.470 174.250 ;
        RECT 69.630 173.970 69.910 174.250 ;
        RECT 70.150 173.970 70.430 174.250 ;
        RECT 53.230 171.330 53.510 171.610 ;
        RECT 53.750 171.330 54.030 171.610 ;
        RECT 57.190 171.330 57.470 171.610 ;
        RECT 57.710 171.330 57.990 171.610 ;
        RECT 65.670 171.330 65.950 171.610 ;
        RECT 66.190 171.330 66.470 171.610 ;
        RECT 69.630 171.330 69.910 171.610 ;
        RECT 70.150 171.330 70.430 171.610 ;
        RECT 59.190 170.890 59.470 171.170 ;
        RECT 59.710 170.890 59.990 171.170 ;
        RECT 63.510 170.890 63.790 171.170 ;
        RECT 64.030 170.890 64.310 171.170 ;
        RECT 57.190 169.570 57.470 169.850 ;
        RECT 57.710 169.570 57.990 169.850 ;
        RECT 65.670 169.570 65.950 169.850 ;
        RECT 66.190 169.570 66.470 169.850 ;
        RECT 53.230 168.690 53.510 168.970 ;
        RECT 53.750 168.690 54.030 168.970 ;
        RECT 57.190 168.690 57.470 168.970 ;
        RECT 57.710 168.690 57.990 168.970 ;
        RECT 65.670 168.690 65.950 168.970 ;
        RECT 66.190 168.690 66.470 168.970 ;
        RECT 69.630 168.690 69.910 168.970 ;
        RECT 70.150 168.690 70.430 168.970 ;
        RECT 53.230 166.930 53.510 167.210 ;
        RECT 53.750 166.930 54.030 167.210 ;
        RECT 57.190 166.930 57.470 167.210 ;
        RECT 57.710 166.930 57.990 167.210 ;
        RECT 65.670 166.930 65.950 167.210 ;
        RECT 66.190 166.930 66.470 167.210 ;
        RECT 69.630 166.930 69.910 167.210 ;
        RECT 70.150 166.930 70.430 167.210 ;
        RECT 54.790 166.310 55.070 166.590 ;
        RECT 54.790 165.790 55.070 166.070 ;
        RECT 68.590 166.310 68.870 166.590 ;
        RECT 68.590 165.790 68.870 166.070 ;
        RECT 53.230 165.170 53.510 165.450 ;
        RECT 53.750 165.170 54.030 165.450 ;
        RECT 57.190 165.170 57.470 165.450 ;
        RECT 57.710 165.170 57.990 165.450 ;
        RECT 65.670 165.170 65.950 165.450 ;
        RECT 66.190 165.170 66.470 165.450 ;
        RECT 69.630 165.170 69.910 165.450 ;
        RECT 70.150 165.170 70.430 165.450 ;
        RECT 53.230 164.290 53.510 164.570 ;
        RECT 53.750 164.290 54.030 164.570 ;
        RECT 57.190 164.290 57.470 164.570 ;
        RECT 57.710 164.290 57.990 164.570 ;
        RECT 65.670 164.290 65.950 164.570 ;
        RECT 66.190 164.290 66.470 164.570 ;
        RECT 69.630 164.290 69.910 164.570 ;
        RECT 70.150 164.290 70.430 164.570 ;
        RECT 53.230 162.530 53.510 162.810 ;
        RECT 53.750 162.530 54.030 162.810 ;
        RECT 57.190 162.530 57.470 162.810 ;
        RECT 57.710 162.530 57.990 162.810 ;
        RECT 65.670 162.530 65.950 162.810 ;
        RECT 66.190 162.530 66.470 162.810 ;
        RECT 69.630 162.530 69.910 162.810 ;
        RECT 70.150 162.530 70.430 162.810 ;
        RECT 55.575 161.910 55.855 162.190 ;
        RECT 55.575 161.390 55.855 161.670 ;
        RECT 67.805 161.910 68.085 162.190 ;
        RECT 67.805 161.390 68.085 161.670 ;
        RECT 53.230 160.770 53.510 161.050 ;
        RECT 53.750 160.770 54.030 161.050 ;
        RECT 57.190 160.770 57.470 161.050 ;
        RECT 57.710 160.770 57.990 161.050 ;
        RECT 53.230 159.890 53.510 160.170 ;
        RECT 53.750 159.890 54.030 160.170 ;
        RECT 57.190 159.890 57.470 160.170 ;
        RECT 57.710 159.890 57.990 160.170 ;
        RECT 53.230 158.130 53.510 158.410 ;
        RECT 53.750 158.130 54.030 158.410 ;
        RECT 57.190 158.130 57.470 158.410 ;
        RECT 57.710 158.130 57.990 158.410 ;
        RECT 56.290 157.510 56.570 157.790 ;
        RECT 56.290 156.990 56.570 157.270 ;
        RECT 53.230 156.370 53.510 156.650 ;
        RECT 53.750 156.370 54.030 156.650 ;
        RECT 57.190 156.370 57.470 156.650 ;
        RECT 57.710 156.370 57.990 156.650 ;
        RECT 53.230 155.490 53.510 155.770 ;
        RECT 53.750 155.490 54.030 155.770 ;
        RECT 57.190 155.490 57.470 155.770 ;
        RECT 57.710 155.490 57.990 155.770 ;
        RECT 53.230 153.730 53.510 154.010 ;
        RECT 53.750 153.730 54.030 154.010 ;
        RECT 57.190 153.730 57.470 154.010 ;
        RECT 57.710 153.730 57.990 154.010 ;
        RECT 53.230 151.970 53.510 152.250 ;
        RECT 53.750 151.970 54.030 152.250 ;
        RECT 57.190 151.970 57.470 152.250 ;
        RECT 57.710 151.970 57.990 152.250 ;
        RECT 50.910 150.650 51.190 150.930 ;
        RECT 51.430 150.650 51.710 150.930 ;
        RECT 53.230 148.450 53.510 148.730 ;
        RECT 53.750 148.450 54.030 148.730 ;
        RECT 57.190 148.450 57.470 148.730 ;
        RECT 57.710 148.450 57.990 148.730 ;
        RECT 59.190 156.810 59.470 157.090 ;
        RECT 59.710 156.810 59.990 157.090 ;
        RECT 63.670 156.810 63.950 157.090 ;
        RECT 64.190 156.810 64.470 157.090 ;
        RECT 59.190 148.890 59.470 149.170 ;
        RECT 59.710 148.890 59.990 149.170 ;
        RECT 59.190 145.370 59.470 145.650 ;
        RECT 59.710 145.370 59.990 145.650 ;
        RECT 53.230 144.930 53.510 145.210 ;
        RECT 53.750 144.930 54.030 145.210 ;
        RECT 57.190 144.930 57.470 145.210 ;
        RECT 57.710 144.930 57.990 145.210 ;
        RECT 53.230 143.170 53.510 143.450 ;
        RECT 53.750 143.170 54.030 143.450 ;
        RECT 57.190 143.170 57.470 143.450 ;
        RECT 57.710 143.170 57.990 143.450 ;
        RECT 53.230 142.290 53.510 142.570 ;
        RECT 53.750 142.290 54.030 142.570 ;
        RECT 57.190 141.410 57.470 141.690 ;
        RECT 57.710 141.410 57.990 141.690 ;
        RECT 57.190 140.530 57.470 140.810 ;
        RECT 57.710 140.530 57.990 140.810 ;
        RECT 53.070 137.890 53.350 138.170 ;
        RECT 53.590 137.890 53.870 138.170 ;
        RECT 57.190 137.890 57.470 138.170 ;
        RECT 57.710 137.890 57.990 138.170 ;
        RECT 44.430 137.010 44.710 137.290 ;
        RECT 44.950 137.010 45.230 137.290 ;
        RECT 53.230 137.010 53.510 137.290 ;
        RECT 53.750 137.010 54.030 137.290 ;
        RECT 38.470 136.570 38.750 136.850 ;
        RECT 38.990 136.570 39.270 136.850 ;
        RECT 59.190 136.570 59.470 136.850 ;
        RECT 59.710 136.570 59.990 136.850 ;
        RECT 63.510 148.890 63.790 149.170 ;
        RECT 64.030 148.890 64.310 149.170 ;
        RECT 65.670 160.770 65.950 161.050 ;
        RECT 66.190 160.770 66.470 161.050 ;
        RECT 69.630 160.770 69.910 161.050 ;
        RECT 70.150 160.770 70.430 161.050 ;
        RECT 65.670 159.890 65.950 160.170 ;
        RECT 66.190 159.890 66.470 160.170 ;
        RECT 69.630 159.890 69.910 160.170 ;
        RECT 70.150 159.890 70.430 160.170 ;
        RECT 65.670 158.130 65.950 158.410 ;
        RECT 66.190 158.130 66.470 158.410 ;
        RECT 69.630 158.130 69.910 158.410 ;
        RECT 70.150 158.130 70.430 158.410 ;
        RECT 67.090 157.510 67.370 157.790 ;
        RECT 67.090 156.990 67.370 157.270 ;
        RECT 65.670 156.370 65.950 156.650 ;
        RECT 66.190 156.370 66.470 156.650 ;
        RECT 69.630 156.370 69.910 156.650 ;
        RECT 70.150 156.370 70.430 156.650 ;
        RECT 65.670 155.490 65.950 155.770 ;
        RECT 66.190 155.490 66.470 155.770 ;
        RECT 69.630 155.490 69.910 155.770 ;
        RECT 70.150 155.490 70.430 155.770 ;
        RECT 65.670 153.730 65.950 154.010 ;
        RECT 66.190 153.730 66.470 154.010 ;
        RECT 69.630 153.730 69.910 154.010 ;
        RECT 70.150 153.730 70.430 154.010 ;
        RECT 65.670 151.970 65.950 152.250 ;
        RECT 66.190 151.970 66.470 152.250 ;
        RECT 69.630 151.970 69.910 152.250 ;
        RECT 70.150 151.970 70.430 152.250 ;
        RECT 71.790 150.650 72.070 150.930 ;
        RECT 72.310 150.650 72.590 150.930 ;
        RECT 65.670 148.450 65.950 148.730 ;
        RECT 66.190 148.450 66.470 148.730 ;
        RECT 69.630 148.450 69.910 148.730 ;
        RECT 70.150 148.450 70.430 148.730 ;
        RECT 63.670 145.370 63.950 145.650 ;
        RECT 64.190 145.370 64.470 145.650 ;
        RECT 65.670 144.930 65.950 145.210 ;
        RECT 66.190 144.930 66.470 145.210 ;
        RECT 69.630 144.930 69.910 145.210 ;
        RECT 70.150 144.930 70.430 145.210 ;
        RECT 65.670 143.170 65.950 143.450 ;
        RECT 66.190 143.170 66.470 143.450 ;
        RECT 69.630 143.170 69.910 143.450 ;
        RECT 70.150 143.170 70.430 143.450 ;
        RECT 69.630 142.290 69.910 142.570 ;
        RECT 70.150 142.290 70.430 142.570 ;
        RECT 65.670 141.410 65.950 141.690 ;
        RECT 66.190 141.410 66.470 141.690 ;
        RECT 65.670 140.530 65.950 140.810 ;
        RECT 66.190 140.530 66.470 140.810 ;
        RECT 65.670 137.890 65.950 138.170 ;
        RECT 66.190 137.890 66.470 138.170 ;
        RECT 69.790 137.890 70.070 138.170 ;
        RECT 70.310 137.890 70.590 138.170 ;
        RECT 78.430 173.970 78.710 174.250 ;
        RECT 78.950 173.970 79.230 174.250 ;
        RECT 82.390 173.970 82.670 174.250 ;
        RECT 82.910 173.970 83.190 174.250 ;
        RECT 113.910 178.810 114.190 179.090 ;
        RECT 114.430 178.810 114.710 179.090 ;
        RECT 90.870 177.490 91.150 177.770 ;
        RECT 91.390 177.490 91.670 177.770 ;
        RECT 94.830 177.490 95.110 177.770 ;
        RECT 95.350 177.490 95.630 177.770 ;
        RECT 103.630 177.490 103.910 177.770 ;
        RECT 104.150 177.490 104.430 177.770 ;
        RECT 107.590 177.490 107.870 177.770 ;
        RECT 108.110 177.490 108.390 177.770 ;
        RECT 90.870 176.610 91.150 176.890 ;
        RECT 91.390 176.610 91.670 176.890 ;
        RECT 107.430 176.610 107.710 176.890 ;
        RECT 107.950 176.610 108.230 176.890 ;
        RECT 90.870 175.730 91.150 176.010 ;
        RECT 91.390 175.730 91.670 176.010 ;
        RECT 94.830 175.730 95.110 176.010 ;
        RECT 95.350 175.730 95.630 176.010 ;
        RECT 103.630 175.730 103.910 176.010 ;
        RECT 104.150 175.730 104.430 176.010 ;
        RECT 107.590 175.730 107.870 176.010 ;
        RECT 108.110 175.730 108.390 176.010 ;
        RECT 90.870 173.970 91.150 174.250 ;
        RECT 91.390 173.970 91.670 174.250 ;
        RECT 94.830 173.970 95.110 174.250 ;
        RECT 95.350 173.970 95.630 174.250 ;
        RECT 78.430 171.330 78.710 171.610 ;
        RECT 78.950 171.330 79.230 171.610 ;
        RECT 82.390 171.330 82.670 171.610 ;
        RECT 82.910 171.330 83.190 171.610 ;
        RECT 90.870 171.330 91.150 171.610 ;
        RECT 91.390 171.330 91.670 171.610 ;
        RECT 94.830 171.330 95.110 171.610 ;
        RECT 95.350 171.330 95.630 171.610 ;
        RECT 84.390 170.890 84.670 171.170 ;
        RECT 84.910 170.890 85.190 171.170 ;
        RECT 88.710 170.890 88.990 171.170 ;
        RECT 89.230 170.890 89.510 171.170 ;
        RECT 82.390 169.570 82.670 169.850 ;
        RECT 82.910 169.570 83.190 169.850 ;
        RECT 90.870 169.570 91.150 169.850 ;
        RECT 91.390 169.570 91.670 169.850 ;
        RECT 78.430 168.690 78.710 168.970 ;
        RECT 78.950 168.690 79.230 168.970 ;
        RECT 82.390 168.690 82.670 168.970 ;
        RECT 82.910 168.690 83.190 168.970 ;
        RECT 90.870 168.690 91.150 168.970 ;
        RECT 91.390 168.690 91.670 168.970 ;
        RECT 94.830 168.690 95.110 168.970 ;
        RECT 95.350 168.690 95.630 168.970 ;
        RECT 78.430 166.930 78.710 167.210 ;
        RECT 78.950 166.930 79.230 167.210 ;
        RECT 82.390 166.930 82.670 167.210 ;
        RECT 82.910 166.930 83.190 167.210 ;
        RECT 90.870 166.930 91.150 167.210 ;
        RECT 91.390 166.930 91.670 167.210 ;
        RECT 94.830 166.930 95.110 167.210 ;
        RECT 95.350 166.930 95.630 167.210 ;
        RECT 79.990 166.310 80.270 166.590 ;
        RECT 79.990 165.790 80.270 166.070 ;
        RECT 93.790 166.310 94.070 166.590 ;
        RECT 93.790 165.790 94.070 166.070 ;
        RECT 78.430 165.170 78.710 165.450 ;
        RECT 78.950 165.170 79.230 165.450 ;
        RECT 82.390 165.170 82.670 165.450 ;
        RECT 82.910 165.170 83.190 165.450 ;
        RECT 90.870 165.170 91.150 165.450 ;
        RECT 91.390 165.170 91.670 165.450 ;
        RECT 94.830 165.170 95.110 165.450 ;
        RECT 95.350 165.170 95.630 165.450 ;
        RECT 78.430 164.290 78.710 164.570 ;
        RECT 78.950 164.290 79.230 164.570 ;
        RECT 82.390 164.290 82.670 164.570 ;
        RECT 82.910 164.290 83.190 164.570 ;
        RECT 90.870 164.290 91.150 164.570 ;
        RECT 91.390 164.290 91.670 164.570 ;
        RECT 94.830 164.290 95.110 164.570 ;
        RECT 95.350 164.290 95.630 164.570 ;
        RECT 78.430 162.530 78.710 162.810 ;
        RECT 78.950 162.530 79.230 162.810 ;
        RECT 82.390 162.530 82.670 162.810 ;
        RECT 82.910 162.530 83.190 162.810 ;
        RECT 90.870 162.530 91.150 162.810 ;
        RECT 91.390 162.530 91.670 162.810 ;
        RECT 94.830 162.530 95.110 162.810 ;
        RECT 95.350 162.530 95.630 162.810 ;
        RECT 80.775 161.910 81.055 162.190 ;
        RECT 80.775 161.390 81.055 161.670 ;
        RECT 93.005 161.910 93.285 162.190 ;
        RECT 93.005 161.390 93.285 161.670 ;
        RECT 78.430 160.770 78.710 161.050 ;
        RECT 78.950 160.770 79.230 161.050 ;
        RECT 82.390 160.770 82.670 161.050 ;
        RECT 82.910 160.770 83.190 161.050 ;
        RECT 78.430 159.890 78.710 160.170 ;
        RECT 78.950 159.890 79.230 160.170 ;
        RECT 82.390 159.890 82.670 160.170 ;
        RECT 82.910 159.890 83.190 160.170 ;
        RECT 78.430 158.130 78.710 158.410 ;
        RECT 78.950 158.130 79.230 158.410 ;
        RECT 82.390 158.130 82.670 158.410 ;
        RECT 82.910 158.130 83.190 158.410 ;
        RECT 81.490 157.510 81.770 157.790 ;
        RECT 81.490 156.990 81.770 157.270 ;
        RECT 78.430 156.370 78.710 156.650 ;
        RECT 78.950 156.370 79.230 156.650 ;
        RECT 82.390 156.370 82.670 156.650 ;
        RECT 82.910 156.370 83.190 156.650 ;
        RECT 78.430 155.490 78.710 155.770 ;
        RECT 78.950 155.490 79.230 155.770 ;
        RECT 82.390 155.490 82.670 155.770 ;
        RECT 82.910 155.490 83.190 155.770 ;
        RECT 78.430 153.730 78.710 154.010 ;
        RECT 78.950 153.730 79.230 154.010 ;
        RECT 82.390 153.730 82.670 154.010 ;
        RECT 82.910 153.730 83.190 154.010 ;
        RECT 78.430 151.970 78.710 152.250 ;
        RECT 78.950 151.970 79.230 152.250 ;
        RECT 82.390 151.970 82.670 152.250 ;
        RECT 82.910 151.970 83.190 152.250 ;
        RECT 76.110 150.650 76.390 150.930 ;
        RECT 76.630 150.650 76.910 150.930 ;
        RECT 78.430 148.450 78.710 148.730 ;
        RECT 78.950 148.450 79.230 148.730 ;
        RECT 82.390 148.450 82.670 148.730 ;
        RECT 82.910 148.450 83.190 148.730 ;
        RECT 84.390 156.810 84.670 157.090 ;
        RECT 84.910 156.810 85.190 157.090 ;
        RECT 88.870 156.810 89.150 157.090 ;
        RECT 89.390 156.810 89.670 157.090 ;
        RECT 84.390 148.890 84.670 149.170 ;
        RECT 84.910 148.890 85.190 149.170 ;
        RECT 84.390 145.370 84.670 145.650 ;
        RECT 84.910 145.370 85.190 145.650 ;
        RECT 78.430 144.930 78.710 145.210 ;
        RECT 78.950 144.930 79.230 145.210 ;
        RECT 82.390 144.930 82.670 145.210 ;
        RECT 82.910 144.930 83.190 145.210 ;
        RECT 78.430 143.170 78.710 143.450 ;
        RECT 78.950 143.170 79.230 143.450 ;
        RECT 82.390 143.170 82.670 143.450 ;
        RECT 82.910 143.170 83.190 143.450 ;
        RECT 78.430 142.290 78.710 142.570 ;
        RECT 78.950 142.290 79.230 142.570 ;
        RECT 82.390 141.410 82.670 141.690 ;
        RECT 82.910 141.410 83.190 141.690 ;
        RECT 82.390 140.530 82.670 140.810 ;
        RECT 82.910 140.530 83.190 140.810 ;
        RECT 78.270 137.890 78.550 138.170 ;
        RECT 78.790 137.890 79.070 138.170 ;
        RECT 82.390 137.890 82.670 138.170 ;
        RECT 82.910 137.890 83.190 138.170 ;
        RECT 69.630 137.010 69.910 137.290 ;
        RECT 70.150 137.010 70.430 137.290 ;
        RECT 78.430 137.010 78.710 137.290 ;
        RECT 78.950 137.010 79.230 137.290 ;
        RECT 63.670 136.570 63.950 136.850 ;
        RECT 64.190 136.570 64.470 136.850 ;
        RECT 84.390 136.570 84.670 136.850 ;
        RECT 84.910 136.570 85.190 136.850 ;
        RECT 88.710 148.890 88.990 149.170 ;
        RECT 89.230 148.890 89.510 149.170 ;
        RECT 90.870 160.770 91.150 161.050 ;
        RECT 91.390 160.770 91.670 161.050 ;
        RECT 94.830 160.770 95.110 161.050 ;
        RECT 95.350 160.770 95.630 161.050 ;
        RECT 90.870 159.890 91.150 160.170 ;
        RECT 91.390 159.890 91.670 160.170 ;
        RECT 94.830 159.890 95.110 160.170 ;
        RECT 95.350 159.890 95.630 160.170 ;
        RECT 90.870 158.130 91.150 158.410 ;
        RECT 91.390 158.130 91.670 158.410 ;
        RECT 94.830 158.130 95.110 158.410 ;
        RECT 95.350 158.130 95.630 158.410 ;
        RECT 92.290 157.510 92.570 157.790 ;
        RECT 92.290 156.990 92.570 157.270 ;
        RECT 90.870 156.370 91.150 156.650 ;
        RECT 91.390 156.370 91.670 156.650 ;
        RECT 94.830 156.370 95.110 156.650 ;
        RECT 95.350 156.370 95.630 156.650 ;
        RECT 90.870 155.490 91.150 155.770 ;
        RECT 91.390 155.490 91.670 155.770 ;
        RECT 94.830 155.490 95.110 155.770 ;
        RECT 95.350 155.490 95.630 155.770 ;
        RECT 90.870 153.730 91.150 154.010 ;
        RECT 91.390 153.730 91.670 154.010 ;
        RECT 94.830 153.730 95.110 154.010 ;
        RECT 95.350 153.730 95.630 154.010 ;
        RECT 90.870 151.970 91.150 152.250 ;
        RECT 91.390 151.970 91.670 152.250 ;
        RECT 94.830 151.970 95.110 152.250 ;
        RECT 95.350 151.970 95.630 152.250 ;
        RECT 96.990 150.650 97.270 150.930 ;
        RECT 97.510 150.650 97.790 150.930 ;
        RECT 90.870 148.450 91.150 148.730 ;
        RECT 91.390 148.450 91.670 148.730 ;
        RECT 94.830 148.450 95.110 148.730 ;
        RECT 95.350 148.450 95.630 148.730 ;
        RECT 88.870 145.370 89.150 145.650 ;
        RECT 89.390 145.370 89.670 145.650 ;
        RECT 90.870 144.930 91.150 145.210 ;
        RECT 91.390 144.930 91.670 145.210 ;
        RECT 94.830 144.930 95.110 145.210 ;
        RECT 95.350 144.930 95.630 145.210 ;
        RECT 90.870 143.170 91.150 143.450 ;
        RECT 91.390 143.170 91.670 143.450 ;
        RECT 94.830 143.170 95.110 143.450 ;
        RECT 95.350 143.170 95.630 143.450 ;
        RECT 94.830 142.290 95.110 142.570 ;
        RECT 95.350 142.290 95.630 142.570 ;
        RECT 90.870 141.410 91.150 141.690 ;
        RECT 91.390 141.410 91.670 141.690 ;
        RECT 90.870 140.530 91.150 140.810 ;
        RECT 91.390 140.530 91.670 140.810 ;
        RECT 90.870 137.890 91.150 138.170 ;
        RECT 91.390 137.890 91.670 138.170 ;
        RECT 94.990 137.890 95.270 138.170 ;
        RECT 95.510 137.890 95.790 138.170 ;
        RECT 103.630 173.970 103.910 174.250 ;
        RECT 104.150 173.970 104.430 174.250 ;
        RECT 107.590 173.970 107.870 174.250 ;
        RECT 108.110 173.970 108.390 174.250 ;
        RECT 122.190 177.930 122.470 178.210 ;
        RECT 122.710 177.930 122.990 178.210 ;
        RECT 116.070 177.490 116.350 177.770 ;
        RECT 116.590 177.490 116.870 177.770 ;
        RECT 120.030 177.490 120.310 177.770 ;
        RECT 120.550 177.490 120.830 177.770 ;
        RECT 120.030 176.610 120.310 176.890 ;
        RECT 120.550 176.610 120.830 176.890 ;
        RECT 116.070 174.850 116.350 175.130 ;
        RECT 116.590 174.850 116.870 175.130 ;
        RECT 120.030 174.850 120.310 175.130 ;
        RECT 120.550 174.850 120.830 175.130 ;
        RECT 109.590 172.650 109.870 172.930 ;
        RECT 110.110 172.650 110.390 172.930 ;
        RECT 103.630 171.330 103.910 171.610 ;
        RECT 104.150 171.330 104.430 171.610 ;
        RECT 107.590 171.330 107.870 171.610 ;
        RECT 108.110 171.330 108.390 171.610 ;
        RECT 109.590 170.890 109.870 171.170 ;
        RECT 110.110 170.890 110.390 171.170 ;
        RECT 107.590 169.570 107.870 169.850 ;
        RECT 108.110 169.570 108.390 169.850 ;
        RECT 103.630 168.690 103.910 168.970 ;
        RECT 104.150 168.690 104.430 168.970 ;
        RECT 107.590 168.690 107.870 168.970 ;
        RECT 108.110 168.690 108.390 168.970 ;
        RECT 103.630 166.930 103.910 167.210 ;
        RECT 104.150 166.930 104.430 167.210 ;
        RECT 107.590 166.930 107.870 167.210 ;
        RECT 108.110 166.930 108.390 167.210 ;
        RECT 116.070 173.090 116.350 173.370 ;
        RECT 116.590 173.090 116.870 173.370 ;
        RECT 120.030 173.090 120.310 173.370 ;
        RECT 120.550 173.090 120.830 173.370 ;
        RECT 140.095 206.345 140.375 206.625 ;
        RECT 140.615 206.345 140.895 206.625 ;
        RECT 144.055 206.345 144.335 206.625 ;
        RECT 144.575 206.345 144.855 206.625 ;
        RECT 140.095 205.465 140.375 205.745 ;
        RECT 140.615 205.465 140.895 205.745 ;
        RECT 144.055 205.465 144.335 205.745 ;
        RECT 144.575 205.465 144.855 205.745 ;
        RECT 140.095 203.705 140.375 203.985 ;
        RECT 140.615 203.705 140.895 203.985 ;
        RECT 144.055 203.705 144.335 203.985 ;
        RECT 144.575 203.705 144.855 203.985 ;
        RECT 140.095 201.945 140.375 202.225 ;
        RECT 140.615 201.945 140.895 202.225 ;
        RECT 144.055 201.945 144.335 202.225 ;
        RECT 144.575 201.945 144.855 202.225 ;
        RECT 140.095 201.065 140.375 201.345 ;
        RECT 140.615 201.065 140.895 201.345 ;
        RECT 144.055 201.065 144.335 201.345 ;
        RECT 144.575 201.065 144.855 201.345 ;
        RECT 126.710 170.220 127.050 170.560 ;
        RECT 105.190 166.310 105.470 166.590 ;
        RECT 105.190 165.790 105.470 166.070 ;
        RECT 103.630 165.170 103.910 165.450 ;
        RECT 104.150 165.170 104.430 165.450 ;
        RECT 107.590 165.170 107.870 165.450 ;
        RECT 108.110 165.170 108.390 165.450 ;
        RECT 103.630 164.290 103.910 164.570 ;
        RECT 104.150 164.290 104.430 164.570 ;
        RECT 107.590 164.290 107.870 164.570 ;
        RECT 108.110 164.290 108.390 164.570 ;
        RECT 103.630 162.530 103.910 162.810 ;
        RECT 104.150 162.530 104.430 162.810 ;
        RECT 107.590 162.530 107.870 162.810 ;
        RECT 108.110 162.530 108.390 162.810 ;
        RECT 105.975 161.910 106.255 162.190 ;
        RECT 105.975 161.390 106.255 161.670 ;
        RECT 103.630 160.770 103.910 161.050 ;
        RECT 104.150 160.770 104.430 161.050 ;
        RECT 107.590 160.770 107.870 161.050 ;
        RECT 108.110 160.770 108.390 161.050 ;
        RECT 103.630 159.890 103.910 160.170 ;
        RECT 104.150 159.890 104.430 160.170 ;
        RECT 107.590 159.890 107.870 160.170 ;
        RECT 108.110 159.890 108.390 160.170 ;
        RECT 103.630 158.130 103.910 158.410 ;
        RECT 104.150 158.130 104.430 158.410 ;
        RECT 107.590 158.130 107.870 158.410 ;
        RECT 108.110 158.130 108.390 158.410 ;
        RECT 106.690 157.510 106.970 157.790 ;
        RECT 106.690 156.990 106.970 157.270 ;
        RECT 103.630 156.370 103.910 156.650 ;
        RECT 104.150 156.370 104.430 156.650 ;
        RECT 107.590 156.370 107.870 156.650 ;
        RECT 108.110 156.370 108.390 156.650 ;
        RECT 103.630 155.490 103.910 155.770 ;
        RECT 104.150 155.490 104.430 155.770 ;
        RECT 107.590 155.490 107.870 155.770 ;
        RECT 108.110 155.490 108.390 155.770 ;
        RECT 103.630 153.730 103.910 154.010 ;
        RECT 104.150 153.730 104.430 154.010 ;
        RECT 107.590 153.730 107.870 154.010 ;
        RECT 108.110 153.730 108.390 154.010 ;
        RECT 103.630 151.970 103.910 152.250 ;
        RECT 104.150 151.970 104.430 152.250 ;
        RECT 107.590 151.970 107.870 152.250 ;
        RECT 108.110 151.970 108.390 152.250 ;
        RECT 101.310 150.650 101.590 150.930 ;
        RECT 101.830 150.650 102.110 150.930 ;
        RECT 103.630 148.450 103.910 148.730 ;
        RECT 104.150 148.450 104.430 148.730 ;
        RECT 107.590 148.450 107.870 148.730 ;
        RECT 108.110 148.450 108.390 148.730 ;
        RECT 109.590 156.810 109.870 157.090 ;
        RECT 110.110 156.810 110.390 157.090 ;
        RECT 109.590 148.890 109.870 149.170 ;
        RECT 110.110 148.890 110.390 149.170 ;
        RECT 109.590 145.370 109.870 145.650 ;
        RECT 110.110 145.370 110.390 145.650 ;
        RECT 103.630 144.930 103.910 145.210 ;
        RECT 104.150 144.930 104.430 145.210 ;
        RECT 107.590 144.930 107.870 145.210 ;
        RECT 108.110 144.930 108.390 145.210 ;
        RECT 103.630 143.170 103.910 143.450 ;
        RECT 104.150 143.170 104.430 143.450 ;
        RECT 107.590 143.170 107.870 143.450 ;
        RECT 108.110 143.170 108.390 143.450 ;
        RECT 103.630 142.290 103.910 142.570 ;
        RECT 104.150 142.290 104.430 142.570 ;
        RECT 107.590 141.410 107.870 141.690 ;
        RECT 108.110 141.410 108.390 141.690 ;
        RECT 107.590 140.530 107.870 140.810 ;
        RECT 108.110 140.530 108.390 140.810 ;
        RECT 103.470 137.890 103.750 138.170 ;
        RECT 103.990 137.890 104.270 138.170 ;
        RECT 107.590 137.890 107.870 138.170 ;
        RECT 108.110 137.890 108.390 138.170 ;
        RECT 94.830 137.010 95.110 137.290 ;
        RECT 95.350 137.010 95.630 137.290 ;
        RECT 103.630 137.010 103.910 137.290 ;
        RECT 104.150 137.010 104.430 137.290 ;
        RECT 88.870 136.570 89.150 136.850 ;
        RECT 89.390 136.570 89.670 136.850 ;
        RECT 109.590 136.570 109.870 136.850 ;
        RECT 110.110 136.570 110.390 136.850 ;
        RECT 120.030 166.930 120.310 167.210 ;
        RECT 120.550 166.930 120.830 167.210 ;
        RECT 116.070 166.050 116.350 166.330 ;
        RECT 116.590 166.050 116.870 166.330 ;
        RECT 120.030 165.170 120.310 165.450 ;
        RECT 120.550 165.170 120.830 165.450 ;
        RECT 113.910 163.850 114.190 164.130 ;
        RECT 114.430 163.850 114.710 164.130 ;
        RECT 120.030 163.410 120.310 163.690 ;
        RECT 120.550 163.410 120.830 163.690 ;
        RECT 120.030 161.650 120.310 161.930 ;
        RECT 120.550 161.650 120.830 161.930 ;
        RECT 120.030 159.890 120.310 160.170 ;
        RECT 120.550 159.890 120.830 160.170 ;
        RECT 116.070 159.010 116.350 159.290 ;
        RECT 116.590 159.010 116.870 159.290 ;
        RECT 116.070 158.130 116.350 158.410 ;
        RECT 116.590 158.130 116.870 158.410 ;
        RECT 120.030 158.130 120.310 158.410 ;
        RECT 120.550 158.130 120.830 158.410 ;
        RECT 116.070 156.370 116.350 156.650 ;
        RECT 116.590 156.370 116.870 156.650 ;
        RECT 120.030 156.370 120.310 156.650 ;
        RECT 120.550 156.370 120.830 156.650 ;
        RECT 120.030 155.490 120.310 155.770 ;
        RECT 120.550 155.490 120.830 155.770 ;
        RECT 116.070 154.610 116.350 154.890 ;
        RECT 116.590 154.610 116.870 154.890 ;
        RECT 120.030 154.610 120.310 154.890 ;
        RECT 120.550 154.610 120.830 154.890 ;
        RECT 116.070 153.730 116.350 154.010 ;
        RECT 116.590 153.730 116.870 154.010 ;
        RECT 120.030 153.730 120.310 154.010 ;
        RECT 120.550 153.730 120.830 154.010 ;
        RECT 116.070 151.970 116.350 152.250 ;
        RECT 116.590 151.970 116.870 152.250 ;
        RECT 120.030 151.970 120.310 152.250 ;
        RECT 120.550 151.970 120.830 152.250 ;
        RECT 116.230 151.260 116.510 151.540 ;
        RECT 116.750 151.260 117.030 151.540 ;
        RECT 122.190 161.210 122.470 161.490 ;
        RECT 122.710 161.210 122.990 161.490 ;
        RECT 116.070 150.210 116.350 150.490 ;
        RECT 116.590 150.210 116.870 150.490 ;
        RECT 120.030 150.210 120.310 150.490 ;
        RECT 120.550 150.210 120.830 150.490 ;
        RECT 120.030 149.330 120.310 149.610 ;
        RECT 120.550 149.330 120.830 149.610 ;
        RECT 120.030 147.570 120.310 147.850 ;
        RECT 120.550 147.570 120.830 147.850 ;
        RECT 120.030 145.810 120.310 146.090 ;
        RECT 120.550 145.810 120.830 146.090 ;
        RECT 122.190 145.370 122.470 145.650 ;
        RECT 122.710 145.370 122.990 145.650 ;
        RECT 120.030 144.050 120.310 144.330 ;
        RECT 120.550 144.050 120.830 144.330 ;
        RECT 116.070 143.170 116.350 143.450 ;
        RECT 116.590 143.170 116.870 143.450 ;
        RECT 113.910 140.970 114.190 141.250 ;
        RECT 114.430 140.970 114.710 141.250 ;
        RECT 120.030 137.010 120.310 137.290 ;
        RECT 120.550 137.010 120.830 137.290 ;
        RECT 116.070 136.130 116.350 136.410 ;
        RECT 116.590 136.130 116.870 136.410 ;
        RECT 15.270 135.250 15.550 135.530 ;
        RECT 15.790 135.250 16.070 135.530 ;
        RECT 19.230 135.250 19.510 135.530 ;
        RECT 19.750 135.250 20.030 135.530 ;
        RECT 28.030 135.250 28.310 135.530 ;
        RECT 28.550 135.250 28.830 135.530 ;
        RECT 31.990 135.250 32.270 135.530 ;
        RECT 32.510 135.250 32.790 135.530 ;
        RECT 40.470 135.250 40.750 135.530 ;
        RECT 40.990 135.250 41.270 135.530 ;
        RECT 44.430 135.250 44.710 135.530 ;
        RECT 44.950 135.250 45.230 135.530 ;
        RECT 53.230 135.250 53.510 135.530 ;
        RECT 53.750 135.250 54.030 135.530 ;
        RECT 57.190 135.250 57.470 135.530 ;
        RECT 57.710 135.250 57.990 135.530 ;
        RECT 65.670 135.250 65.950 135.530 ;
        RECT 66.190 135.250 66.470 135.530 ;
        RECT 69.630 135.250 69.910 135.530 ;
        RECT 70.150 135.250 70.430 135.530 ;
        RECT 78.430 135.250 78.710 135.530 ;
        RECT 78.950 135.250 79.230 135.530 ;
        RECT 82.390 135.250 82.670 135.530 ;
        RECT 82.910 135.250 83.190 135.530 ;
        RECT 90.870 135.250 91.150 135.530 ;
        RECT 91.390 135.250 91.670 135.530 ;
        RECT 94.830 135.250 95.110 135.530 ;
        RECT 95.350 135.250 95.630 135.530 ;
        RECT 103.630 135.250 103.910 135.530 ;
        RECT 104.150 135.250 104.430 135.530 ;
        RECT 107.590 135.250 107.870 135.530 ;
        RECT 108.110 135.250 108.390 135.530 ;
        RECT 116.070 135.250 116.350 135.530 ;
        RECT 116.590 135.250 116.870 135.530 ;
        RECT 120.030 135.250 120.310 135.530 ;
        RECT 120.550 135.250 120.830 135.530 ;
        RECT 15.270 134.370 15.550 134.650 ;
        RECT 15.790 134.370 16.070 134.650 ;
        RECT 19.230 134.370 19.510 134.650 ;
        RECT 19.750 134.370 20.030 134.650 ;
        RECT 28.030 134.370 28.310 134.650 ;
        RECT 28.550 134.370 28.830 134.650 ;
        RECT 31.990 134.370 32.270 134.650 ;
        RECT 32.510 134.370 32.790 134.650 ;
        RECT 40.470 134.370 40.750 134.650 ;
        RECT 40.990 134.370 41.270 134.650 ;
        RECT 44.430 134.370 44.710 134.650 ;
        RECT 44.950 134.370 45.230 134.650 ;
        RECT 53.230 134.370 53.510 134.650 ;
        RECT 53.750 134.370 54.030 134.650 ;
        RECT 57.190 134.370 57.470 134.650 ;
        RECT 57.710 134.370 57.990 134.650 ;
        RECT 65.670 134.370 65.950 134.650 ;
        RECT 66.190 134.370 66.470 134.650 ;
        RECT 69.630 134.370 69.910 134.650 ;
        RECT 70.150 134.370 70.430 134.650 ;
        RECT 78.430 134.370 78.710 134.650 ;
        RECT 78.950 134.370 79.230 134.650 ;
        RECT 82.390 134.370 82.670 134.650 ;
        RECT 82.910 134.370 83.190 134.650 ;
        RECT 90.870 134.370 91.150 134.650 ;
        RECT 91.390 134.370 91.670 134.650 ;
        RECT 94.830 134.370 95.110 134.650 ;
        RECT 95.350 134.370 95.630 134.650 ;
        RECT 103.630 134.370 103.910 134.650 ;
        RECT 104.150 134.370 104.430 134.650 ;
        RECT 107.590 134.370 107.870 134.650 ;
        RECT 108.110 134.370 108.390 134.650 ;
        RECT 116.070 134.370 116.350 134.650 ;
        RECT 116.590 134.370 116.870 134.650 ;
        RECT 120.030 134.370 120.310 134.650 ;
        RECT 120.550 134.370 120.830 134.650 ;
        RECT 69.590 130.640 69.870 130.920 ;
        RECT 69.590 130.120 69.870 130.400 ;
        RECT 62.630 124.130 62.910 124.410 ;
        RECT 62.630 123.610 62.910 123.890 ;
        RECT 60.750 123.200 61.030 123.480 ;
        RECT 60.750 122.680 61.030 122.960 ;
        RECT 58.870 122.270 59.150 122.550 ;
        RECT 58.870 121.750 59.150 122.030 ;
        RECT 57.930 115.760 58.210 116.040 ;
        RECT 57.930 115.240 58.210 115.520 ;
        RECT 12.270 97.500 12.550 97.780 ;
        RECT 12.270 96.980 12.550 97.260 ;
        RECT 13.590 93.430 13.870 93.710 ;
        RECT 13.590 92.910 13.870 93.190 ;
        RECT 14.910 93.430 15.190 93.710 ;
        RECT 14.910 92.910 15.190 93.190 ;
        RECT 16.230 93.430 16.510 93.710 ;
        RECT 16.230 92.910 16.510 93.190 ;
        RECT 17.550 93.430 17.830 93.710 ;
        RECT 17.550 92.910 17.830 93.190 ;
        RECT 18.870 99.470 19.150 99.750 ;
        RECT 18.870 98.950 19.150 99.230 ;
        RECT 20.190 99.470 20.470 99.750 ;
        RECT 20.190 98.950 20.470 99.230 ;
        RECT 21.510 102.490 21.790 102.770 ;
        RECT 21.510 101.970 21.790 102.250 ;
        RECT 22.830 105.510 23.110 105.790 ;
        RECT 22.830 104.990 23.110 105.270 ;
        RECT 24.150 96.450 24.430 96.730 ;
        RECT 24.150 95.930 24.430 96.210 ;
        RECT 25.470 102.490 25.750 102.770 ;
        RECT 25.470 101.970 25.750 102.250 ;
        RECT 26.790 99.470 27.070 99.750 ;
        RECT 26.790 98.950 27.070 99.230 ;
        RECT 28.110 99.470 28.390 99.750 ;
        RECT 28.110 98.950 28.390 99.230 ;
        RECT 29.430 93.430 29.710 93.710 ;
        RECT 29.430 92.910 29.710 93.190 ;
        RECT 30.750 93.430 31.030 93.710 ;
        RECT 30.750 92.910 31.030 93.190 ;
        RECT 32.070 93.430 32.350 93.710 ;
        RECT 32.070 92.910 32.350 93.190 ;
        RECT 33.390 93.430 33.670 93.710 ;
        RECT 33.390 92.910 33.670 93.190 ;
        RECT 34.710 93.430 34.990 93.710 ;
        RECT 34.710 92.910 34.990 93.190 ;
        RECT 36.030 93.430 36.310 93.710 ;
        RECT 36.030 92.910 36.310 93.190 ;
        RECT 37.350 93.430 37.630 93.710 ;
        RECT 37.350 92.910 37.630 93.190 ;
        RECT 38.670 93.430 38.950 93.710 ;
        RECT 38.670 92.910 38.950 93.190 ;
        RECT 39.990 99.470 40.270 99.750 ;
        RECT 39.990 98.950 40.270 99.230 ;
        RECT 41.310 99.470 41.590 99.750 ;
        RECT 41.310 98.950 41.590 99.230 ;
        RECT 42.630 102.490 42.910 102.770 ;
        RECT 42.630 101.970 42.910 102.250 ;
        RECT 43.950 96.450 44.230 96.730 ;
        RECT 43.950 95.930 44.230 96.210 ;
        RECT 45.270 90.410 45.550 90.690 ;
        RECT 45.270 89.890 45.550 90.170 ;
        RECT 46.590 102.490 46.870 102.770 ;
        RECT 46.590 101.970 46.870 102.250 ;
        RECT 47.910 99.470 48.190 99.750 ;
        RECT 47.910 98.950 48.190 99.230 ;
        RECT 49.230 99.470 49.510 99.750 ;
        RECT 49.230 98.950 49.510 99.230 ;
        RECT 50.550 93.430 50.830 93.710 ;
        RECT 50.550 92.910 50.830 93.190 ;
        RECT 51.870 93.430 52.150 93.710 ;
        RECT 51.870 92.910 52.150 93.190 ;
        RECT 53.190 93.430 53.470 93.710 ;
        RECT 53.190 92.910 53.470 93.190 ;
        RECT 54.510 93.430 54.790 93.710 ;
        RECT 54.510 92.910 54.790 93.190 ;
        RECT 56.180 105.250 56.460 105.530 ;
        RECT 56.700 105.250 56.980 105.530 ;
        RECT 57.930 105.510 58.210 105.790 ;
        RECT 57.930 104.990 58.210 105.270 ;
        RECT 56.180 102.230 56.460 102.510 ;
        RECT 56.700 102.230 56.980 102.510 ;
        RECT 57.930 102.490 58.210 102.770 ;
        RECT 57.930 101.970 58.210 102.250 ;
        RECT 56.180 99.210 56.460 99.490 ;
        RECT 56.700 99.210 56.980 99.490 ;
        RECT 57.930 99.470 58.210 99.750 ;
        RECT 57.930 98.950 58.210 99.230 ;
        RECT 56.180 96.190 56.460 96.470 ;
        RECT 56.700 96.190 56.980 96.470 ;
        RECT 57.930 96.450 58.210 96.730 ;
        RECT 57.930 95.930 58.210 96.210 ;
        RECT 56.180 93.170 56.460 93.450 ;
        RECT 56.700 93.170 56.980 93.450 ;
        RECT 57.930 93.430 58.210 93.710 ;
        RECT 57.930 92.910 58.210 93.190 ;
        RECT 56.180 90.150 56.460 90.430 ;
        RECT 56.700 90.150 56.980 90.430 ;
        RECT 57.930 90.410 58.210 90.690 ;
        RECT 57.930 89.890 58.210 90.170 ;
        RECT 12.270 80.500 12.550 80.780 ;
        RECT 12.270 79.980 12.550 80.260 ;
        RECT 13.590 76.430 13.870 76.710 ;
        RECT 13.590 75.910 13.870 76.190 ;
        RECT 14.910 76.430 15.190 76.710 ;
        RECT 14.910 75.910 15.190 76.190 ;
        RECT 16.230 76.430 16.510 76.710 ;
        RECT 16.230 75.910 16.510 76.190 ;
        RECT 17.550 76.430 17.830 76.710 ;
        RECT 17.550 75.910 17.830 76.190 ;
        RECT 18.870 82.470 19.150 82.750 ;
        RECT 18.870 81.950 19.150 82.230 ;
        RECT 20.190 82.470 20.470 82.750 ;
        RECT 20.190 81.950 20.470 82.230 ;
        RECT 21.510 85.490 21.790 85.770 ;
        RECT 21.510 84.970 21.790 85.250 ;
        RECT 22.830 88.510 23.110 88.790 ;
        RECT 22.830 87.990 23.110 88.270 ;
        RECT 24.150 79.450 24.430 79.730 ;
        RECT 24.150 78.930 24.430 79.210 ;
        RECT 25.470 85.490 25.750 85.770 ;
        RECT 25.470 84.970 25.750 85.250 ;
        RECT 26.790 82.470 27.070 82.750 ;
        RECT 26.790 81.950 27.070 82.230 ;
        RECT 28.110 82.470 28.390 82.750 ;
        RECT 28.110 81.950 28.390 82.230 ;
        RECT 29.430 76.430 29.710 76.710 ;
        RECT 29.430 75.910 29.710 76.190 ;
        RECT 30.750 76.430 31.030 76.710 ;
        RECT 30.750 75.910 31.030 76.190 ;
        RECT 32.070 76.430 32.350 76.710 ;
        RECT 32.070 75.910 32.350 76.190 ;
        RECT 33.390 76.430 33.670 76.710 ;
        RECT 33.390 75.910 33.670 76.190 ;
        RECT 34.710 76.430 34.990 76.710 ;
        RECT 34.710 75.910 34.990 76.190 ;
        RECT 36.030 76.430 36.310 76.710 ;
        RECT 36.030 75.910 36.310 76.190 ;
        RECT 37.350 76.430 37.630 76.710 ;
        RECT 37.350 75.910 37.630 76.190 ;
        RECT 38.670 76.430 38.950 76.710 ;
        RECT 38.670 75.910 38.950 76.190 ;
        RECT 39.990 82.470 40.270 82.750 ;
        RECT 39.990 81.950 40.270 82.230 ;
        RECT 41.310 82.470 41.590 82.750 ;
        RECT 41.310 81.950 41.590 82.230 ;
        RECT 42.630 85.490 42.910 85.770 ;
        RECT 42.630 84.970 42.910 85.250 ;
        RECT 43.950 79.450 44.230 79.730 ;
        RECT 43.950 78.930 44.230 79.210 ;
        RECT 45.270 73.410 45.550 73.690 ;
        RECT 45.270 72.890 45.550 73.170 ;
        RECT 46.590 85.490 46.870 85.770 ;
        RECT 46.590 84.970 46.870 85.250 ;
        RECT 47.910 82.470 48.190 82.750 ;
        RECT 47.910 81.950 48.190 82.230 ;
        RECT 49.230 82.470 49.510 82.750 ;
        RECT 49.230 81.950 49.510 82.230 ;
        RECT 50.550 76.430 50.830 76.710 ;
        RECT 50.550 75.910 50.830 76.190 ;
        RECT 51.870 76.430 52.150 76.710 ;
        RECT 51.870 75.910 52.150 76.190 ;
        RECT 53.190 76.430 53.470 76.710 ;
        RECT 53.190 75.910 53.470 76.190 ;
        RECT 54.510 76.430 54.790 76.710 ;
        RECT 54.510 75.910 54.790 76.190 ;
        RECT 56.180 88.250 56.460 88.530 ;
        RECT 56.700 88.250 56.980 88.530 ;
        RECT 56.180 85.230 56.460 85.510 ;
        RECT 56.700 85.230 56.980 85.510 ;
        RECT 56.180 82.210 56.460 82.490 ;
        RECT 56.700 82.210 56.980 82.490 ;
        RECT 56.180 79.190 56.460 79.470 ;
        RECT 56.700 79.190 56.980 79.470 ;
        RECT 56.180 76.170 56.460 76.450 ;
        RECT 56.700 76.170 56.980 76.450 ;
        RECT 56.180 73.150 56.460 73.430 ;
        RECT 56.700 73.150 56.980 73.430 ;
        RECT 12.270 63.500 12.550 63.780 ;
        RECT 12.270 62.980 12.550 63.260 ;
        RECT 13.590 59.430 13.870 59.710 ;
        RECT 13.590 58.910 13.870 59.190 ;
        RECT 14.910 59.430 15.190 59.710 ;
        RECT 14.910 58.910 15.190 59.190 ;
        RECT 16.230 59.430 16.510 59.710 ;
        RECT 16.230 58.910 16.510 59.190 ;
        RECT 17.550 59.430 17.830 59.710 ;
        RECT 17.550 58.910 17.830 59.190 ;
        RECT 18.870 65.470 19.150 65.750 ;
        RECT 18.870 64.950 19.150 65.230 ;
        RECT 20.190 65.470 20.470 65.750 ;
        RECT 20.190 64.950 20.470 65.230 ;
        RECT 21.510 68.490 21.790 68.770 ;
        RECT 21.510 67.970 21.790 68.250 ;
        RECT 22.830 71.510 23.110 71.790 ;
        RECT 22.830 70.990 23.110 71.270 ;
        RECT 24.150 62.450 24.430 62.730 ;
        RECT 24.150 61.930 24.430 62.210 ;
        RECT 25.470 68.490 25.750 68.770 ;
        RECT 25.470 67.970 25.750 68.250 ;
        RECT 26.790 65.470 27.070 65.750 ;
        RECT 26.790 64.950 27.070 65.230 ;
        RECT 28.110 65.470 28.390 65.750 ;
        RECT 28.110 64.950 28.390 65.230 ;
        RECT 29.430 59.430 29.710 59.710 ;
        RECT 29.430 58.910 29.710 59.190 ;
        RECT 30.750 59.430 31.030 59.710 ;
        RECT 30.750 58.910 31.030 59.190 ;
        RECT 32.070 59.430 32.350 59.710 ;
        RECT 32.070 58.910 32.350 59.190 ;
        RECT 33.390 59.430 33.670 59.710 ;
        RECT 33.390 58.910 33.670 59.190 ;
        RECT 34.710 59.430 34.990 59.710 ;
        RECT 34.710 58.910 34.990 59.190 ;
        RECT 36.030 59.430 36.310 59.710 ;
        RECT 36.030 58.910 36.310 59.190 ;
        RECT 37.350 59.430 37.630 59.710 ;
        RECT 37.350 58.910 37.630 59.190 ;
        RECT 38.670 59.430 38.950 59.710 ;
        RECT 38.670 58.910 38.950 59.190 ;
        RECT 39.990 65.470 40.270 65.750 ;
        RECT 39.990 64.950 40.270 65.230 ;
        RECT 41.310 65.470 41.590 65.750 ;
        RECT 41.310 64.950 41.590 65.230 ;
        RECT 42.630 68.490 42.910 68.770 ;
        RECT 42.630 67.970 42.910 68.250 ;
        RECT 43.950 62.450 44.230 62.730 ;
        RECT 43.950 61.930 44.230 62.210 ;
        RECT 45.270 56.410 45.550 56.690 ;
        RECT 45.270 55.890 45.550 56.170 ;
        RECT 46.590 68.490 46.870 68.770 ;
        RECT 46.590 67.970 46.870 68.250 ;
        RECT 47.910 65.470 48.190 65.750 ;
        RECT 47.910 64.950 48.190 65.230 ;
        RECT 49.230 65.470 49.510 65.750 ;
        RECT 49.230 64.950 49.510 65.230 ;
        RECT 50.550 59.430 50.830 59.710 ;
        RECT 50.550 58.910 50.830 59.190 ;
        RECT 51.870 59.430 52.150 59.710 ;
        RECT 51.870 58.910 52.150 59.190 ;
        RECT 53.190 59.430 53.470 59.710 ;
        RECT 53.190 58.910 53.470 59.190 ;
        RECT 54.510 59.430 54.790 59.710 ;
        RECT 54.510 58.910 54.790 59.190 ;
        RECT 56.180 71.250 56.460 71.530 ;
        RECT 56.700 71.250 56.980 71.530 ;
        RECT 56.180 68.230 56.460 68.510 ;
        RECT 56.700 68.230 56.980 68.510 ;
        RECT 56.180 65.210 56.460 65.490 ;
        RECT 56.700 65.210 56.980 65.490 ;
        RECT 56.180 62.190 56.460 62.470 ;
        RECT 56.700 62.190 56.980 62.470 ;
        RECT 56.180 59.170 56.460 59.450 ;
        RECT 56.700 59.170 56.980 59.450 ;
        RECT 12.270 46.500 12.550 46.780 ;
        RECT 12.270 45.980 12.550 46.260 ;
        RECT 13.590 42.430 13.870 42.710 ;
        RECT 13.590 41.910 13.870 42.190 ;
        RECT 14.910 42.430 15.190 42.710 ;
        RECT 14.910 41.910 15.190 42.190 ;
        RECT 16.230 42.430 16.510 42.710 ;
        RECT 16.230 41.910 16.510 42.190 ;
        RECT 17.550 42.430 17.830 42.710 ;
        RECT 17.550 41.910 17.830 42.190 ;
        RECT 18.870 48.470 19.150 48.750 ;
        RECT 18.870 47.950 19.150 48.230 ;
        RECT 20.190 48.470 20.470 48.750 ;
        RECT 20.190 47.950 20.470 48.230 ;
        RECT 21.510 51.490 21.790 51.770 ;
        RECT 21.510 50.970 21.790 51.250 ;
        RECT 22.830 54.510 23.110 54.790 ;
        RECT 22.830 53.990 23.110 54.270 ;
        RECT 24.150 45.450 24.430 45.730 ;
        RECT 24.150 44.930 24.430 45.210 ;
        RECT 25.470 51.490 25.750 51.770 ;
        RECT 25.470 50.970 25.750 51.250 ;
        RECT 26.790 48.470 27.070 48.750 ;
        RECT 26.790 47.950 27.070 48.230 ;
        RECT 28.110 48.470 28.390 48.750 ;
        RECT 28.110 47.950 28.390 48.230 ;
        RECT 29.430 42.430 29.710 42.710 ;
        RECT 29.430 41.910 29.710 42.190 ;
        RECT 30.750 42.430 31.030 42.710 ;
        RECT 30.750 41.910 31.030 42.190 ;
        RECT 32.070 42.430 32.350 42.710 ;
        RECT 32.070 41.910 32.350 42.190 ;
        RECT 33.390 42.430 33.670 42.710 ;
        RECT 33.390 41.910 33.670 42.190 ;
        RECT 34.710 42.430 34.990 42.710 ;
        RECT 34.710 41.910 34.990 42.190 ;
        RECT 36.030 42.430 36.310 42.710 ;
        RECT 36.030 41.910 36.310 42.190 ;
        RECT 37.350 42.430 37.630 42.710 ;
        RECT 37.350 41.910 37.630 42.190 ;
        RECT 38.670 42.430 38.950 42.710 ;
        RECT 38.670 41.910 38.950 42.190 ;
        RECT 39.990 48.470 40.270 48.750 ;
        RECT 39.990 47.950 40.270 48.230 ;
        RECT 41.310 48.470 41.590 48.750 ;
        RECT 41.310 47.950 41.590 48.230 ;
        RECT 42.630 51.490 42.910 51.770 ;
        RECT 42.630 50.970 42.910 51.250 ;
        RECT 43.950 45.450 44.230 45.730 ;
        RECT 43.950 44.930 44.230 45.210 ;
        RECT 45.270 39.410 45.550 39.690 ;
        RECT 45.270 38.890 45.550 39.170 ;
        RECT 46.590 51.490 46.870 51.770 ;
        RECT 46.590 50.970 46.870 51.250 ;
        RECT 47.910 48.470 48.190 48.750 ;
        RECT 47.910 47.950 48.190 48.230 ;
        RECT 49.230 48.470 49.510 48.750 ;
        RECT 49.230 47.950 49.510 48.230 ;
        RECT 50.550 42.430 50.830 42.710 ;
        RECT 50.550 41.910 50.830 42.190 ;
        RECT 51.870 42.430 52.150 42.710 ;
        RECT 51.870 41.910 52.150 42.190 ;
        RECT 53.190 42.430 53.470 42.710 ;
        RECT 53.190 41.910 53.470 42.190 ;
        RECT 54.510 42.430 54.790 42.710 ;
        RECT 54.510 41.910 54.790 42.190 ;
        RECT 59.810 116.690 60.090 116.970 ;
        RECT 59.810 116.170 60.090 116.450 ;
        RECT 60.750 76.430 61.030 76.710 ;
        RECT 60.750 75.910 61.030 76.190 ;
        RECT 61.690 117.620 61.970 117.900 ;
        RECT 61.690 117.100 61.970 117.380 ;
        RECT 61.690 88.510 61.970 88.790 ;
        RECT 61.690 87.990 61.970 88.270 ;
        RECT 61.690 85.490 61.970 85.770 ;
        RECT 61.690 84.970 61.970 85.250 ;
        RECT 66.390 121.340 66.670 121.620 ;
        RECT 66.390 120.820 66.670 121.100 ;
        RECT 65.450 120.410 65.730 120.690 ;
        RECT 65.450 119.890 65.730 120.170 ;
        RECT 64.510 119.480 64.790 119.760 ;
        RECT 64.510 118.960 64.790 119.240 ;
        RECT 62.630 82.470 62.910 82.750 ;
        RECT 62.630 81.950 62.910 82.230 ;
        RECT 63.570 118.550 63.850 118.830 ;
        RECT 63.570 118.030 63.850 118.310 ;
        RECT 61.690 79.450 61.970 79.730 ;
        RECT 61.690 78.930 61.970 79.210 ;
        RECT 61.690 73.410 61.970 73.690 ;
        RECT 61.690 72.890 61.970 73.170 ;
        RECT 64.510 68.490 64.790 68.770 ;
        RECT 64.510 67.970 64.790 68.250 ;
        RECT 63.570 65.470 63.850 65.750 ;
        RECT 63.570 64.950 63.850 65.230 ;
        RECT 66.390 71.510 66.670 71.790 ;
        RECT 66.390 70.990 66.670 71.270 ;
        RECT 69.590 71.510 69.870 71.790 ;
        RECT 69.590 70.990 69.870 71.270 ;
        RECT 70.530 129.710 70.810 129.990 ;
        RECT 70.530 129.190 70.810 129.470 ;
        RECT 65.450 62.450 65.730 62.730 ;
        RECT 65.450 61.930 65.730 62.210 ;
        RECT 71.470 128.780 71.750 129.060 ;
        RECT 71.470 128.260 71.750 128.540 ;
        RECT 71.470 68.490 71.750 68.770 ;
        RECT 71.470 67.970 71.750 68.250 ;
        RECT 72.410 127.850 72.690 128.130 ;
        RECT 72.410 127.330 72.690 127.610 ;
        RECT 73.350 126.920 73.630 127.200 ;
        RECT 73.350 126.400 73.630 126.680 ;
        RECT 75.230 125.990 75.510 126.270 ;
        RECT 75.230 125.470 75.510 125.750 ;
        RECT 73.350 82.470 73.630 82.750 ;
        RECT 73.350 81.950 73.630 82.230 ;
        RECT 74.290 114.830 74.570 115.110 ;
        RECT 74.290 114.310 74.570 114.590 ;
        RECT 74.290 88.510 74.570 88.790 ;
        RECT 74.290 87.990 74.570 88.270 ;
        RECT 74.290 85.490 74.570 85.770 ;
        RECT 74.290 84.970 74.570 85.250 ;
        RECT 74.290 79.450 74.570 79.730 ;
        RECT 74.290 78.930 74.570 79.210 ;
        RECT 77.110 125.060 77.390 125.340 ;
        RECT 77.110 124.540 77.390 124.820 ;
        RECT 75.230 76.430 75.510 76.710 ;
        RECT 75.230 75.910 75.510 76.190 ;
        RECT 76.170 113.900 76.450 114.180 ;
        RECT 76.170 113.380 76.450 113.660 ;
        RECT 74.290 73.410 74.570 73.690 ;
        RECT 74.290 72.890 74.570 73.170 ;
        RECT 72.410 65.470 72.690 65.750 ;
        RECT 72.410 64.950 72.690 65.230 ;
        RECT 70.530 62.450 70.810 62.730 ;
        RECT 70.530 61.930 70.810 62.210 ;
        RECT 59.810 59.430 60.090 59.710 ;
        RECT 59.810 58.910 60.090 59.190 ;
        RECT 76.170 59.430 76.450 59.710 ;
        RECT 76.170 58.910 76.450 59.190 ;
        RECT 56.180 54.250 56.460 54.530 ;
        RECT 56.700 54.250 56.980 54.530 ;
        RECT 58.870 54.510 59.150 54.790 ;
        RECT 58.870 53.990 59.150 54.270 ;
        RECT 56.180 51.230 56.460 51.510 ;
        RECT 56.700 51.230 56.980 51.510 ;
        RECT 58.870 51.490 59.150 51.770 ;
        RECT 58.870 50.970 59.150 51.250 ;
        RECT 56.180 48.210 56.460 48.490 ;
        RECT 56.700 48.210 56.980 48.490 ;
        RECT 58.870 48.470 59.150 48.750 ;
        RECT 58.870 47.950 59.150 48.230 ;
        RECT 56.180 45.190 56.460 45.470 ;
        RECT 56.700 45.190 56.980 45.470 ;
        RECT 58.870 45.450 59.150 45.730 ;
        RECT 58.870 44.930 59.150 45.210 ;
        RECT 56.180 42.170 56.460 42.450 ;
        RECT 56.700 42.170 56.980 42.450 ;
        RECT 58.870 42.430 59.150 42.710 ;
        RECT 58.870 41.910 59.150 42.190 ;
        RECT 56.180 39.150 56.460 39.430 ;
        RECT 56.700 39.150 56.980 39.430 ;
        RECT 58.870 39.410 59.150 39.690 ;
        RECT 58.870 38.890 59.150 39.170 ;
        RECT 78.050 112.970 78.330 113.250 ;
        RECT 78.050 112.450 78.330 112.730 ;
        RECT 78.050 105.510 78.330 105.790 ;
        RECT 78.050 104.990 78.330 105.270 ;
        RECT 79.280 105.250 79.560 105.530 ;
        RECT 79.800 105.250 80.080 105.530 ;
        RECT 78.050 102.490 78.330 102.770 ;
        RECT 78.050 101.970 78.330 102.250 ;
        RECT 79.280 102.230 79.560 102.510 ;
        RECT 79.800 102.230 80.080 102.510 ;
        RECT 78.050 99.470 78.330 99.750 ;
        RECT 78.050 98.950 78.330 99.230 ;
        RECT 79.280 99.210 79.560 99.490 ;
        RECT 79.800 99.210 80.080 99.490 ;
        RECT 78.050 96.450 78.330 96.730 ;
        RECT 78.050 95.930 78.330 96.210 ;
        RECT 79.280 96.190 79.560 96.470 ;
        RECT 79.800 96.190 80.080 96.470 ;
        RECT 78.050 93.430 78.330 93.710 ;
        RECT 78.050 92.910 78.330 93.190 ;
        RECT 79.280 93.170 79.560 93.450 ;
        RECT 79.800 93.170 80.080 93.450 ;
        RECT 78.050 90.410 78.330 90.690 ;
        RECT 78.050 89.890 78.330 90.170 ;
        RECT 79.280 90.150 79.560 90.430 ;
        RECT 79.800 90.150 80.080 90.430 ;
        RECT 81.470 93.430 81.750 93.710 ;
        RECT 81.470 92.910 81.750 93.190 ;
        RECT 82.790 93.430 83.070 93.710 ;
        RECT 82.790 92.910 83.070 93.190 ;
        RECT 84.110 93.430 84.390 93.710 ;
        RECT 84.110 92.910 84.390 93.190 ;
        RECT 85.430 93.430 85.710 93.710 ;
        RECT 85.430 92.910 85.710 93.190 ;
        RECT 86.750 99.470 87.030 99.750 ;
        RECT 86.750 98.950 87.030 99.230 ;
        RECT 88.070 99.470 88.350 99.750 ;
        RECT 88.070 98.950 88.350 99.230 ;
        RECT 89.390 102.490 89.670 102.770 ;
        RECT 89.390 101.970 89.670 102.250 ;
        RECT 90.710 90.410 90.990 90.690 ;
        RECT 90.710 89.890 90.990 90.170 ;
        RECT 92.030 96.450 92.310 96.730 ;
        RECT 92.030 95.930 92.310 96.210 ;
        RECT 93.350 102.490 93.630 102.770 ;
        RECT 93.350 101.970 93.630 102.250 ;
        RECT 94.670 99.470 94.950 99.750 ;
        RECT 94.670 98.950 94.950 99.230 ;
        RECT 95.990 99.470 96.270 99.750 ;
        RECT 95.990 98.950 96.270 99.230 ;
        RECT 97.310 93.430 97.590 93.710 ;
        RECT 97.310 92.910 97.590 93.190 ;
        RECT 98.630 93.430 98.910 93.710 ;
        RECT 98.630 92.910 98.910 93.190 ;
        RECT 99.950 93.430 100.230 93.710 ;
        RECT 99.950 92.910 100.230 93.190 ;
        RECT 101.270 93.430 101.550 93.710 ;
        RECT 101.270 92.910 101.550 93.190 ;
        RECT 102.590 93.430 102.870 93.710 ;
        RECT 102.590 92.910 102.870 93.190 ;
        RECT 103.910 93.430 104.190 93.710 ;
        RECT 103.910 92.910 104.190 93.190 ;
        RECT 105.230 93.430 105.510 93.710 ;
        RECT 105.230 92.910 105.510 93.190 ;
        RECT 106.550 93.430 106.830 93.710 ;
        RECT 106.550 92.910 106.830 93.190 ;
        RECT 107.870 99.470 108.150 99.750 ;
        RECT 107.870 98.950 108.150 99.230 ;
        RECT 109.190 99.470 109.470 99.750 ;
        RECT 109.190 98.950 109.470 99.230 ;
        RECT 110.510 102.490 110.790 102.770 ;
        RECT 110.510 101.970 110.790 102.250 ;
        RECT 111.830 96.450 112.110 96.730 ;
        RECT 111.830 95.930 112.110 96.210 ;
        RECT 113.150 105.510 113.430 105.790 ;
        RECT 113.150 104.990 113.430 105.270 ;
        RECT 114.470 102.490 114.750 102.770 ;
        RECT 114.470 101.970 114.750 102.250 ;
        RECT 115.790 99.470 116.070 99.750 ;
        RECT 115.790 98.950 116.070 99.230 ;
        RECT 117.110 99.470 117.390 99.750 ;
        RECT 117.110 98.950 117.390 99.230 ;
        RECT 118.430 93.430 118.710 93.710 ;
        RECT 118.430 92.910 118.710 93.190 ;
        RECT 119.750 93.430 120.030 93.710 ;
        RECT 119.750 92.910 120.030 93.190 ;
        RECT 121.070 93.430 121.350 93.710 ;
        RECT 121.070 92.910 121.350 93.190 ;
        RECT 122.390 93.430 122.670 93.710 ;
        RECT 122.390 92.910 122.670 93.190 ;
        RECT 123.710 97.500 123.990 97.780 ;
        RECT 123.710 96.980 123.990 97.260 ;
        RECT 79.280 88.250 79.560 88.530 ;
        RECT 79.800 88.250 80.080 88.530 ;
        RECT 79.280 85.230 79.560 85.510 ;
        RECT 79.800 85.230 80.080 85.510 ;
        RECT 79.280 82.210 79.560 82.490 ;
        RECT 79.800 82.210 80.080 82.490 ;
        RECT 79.280 79.190 79.560 79.470 ;
        RECT 79.800 79.190 80.080 79.470 ;
        RECT 79.280 76.170 79.560 76.450 ;
        RECT 79.800 76.170 80.080 76.450 ;
        RECT 79.280 73.150 79.560 73.430 ;
        RECT 79.800 73.150 80.080 73.430 ;
        RECT 81.470 76.430 81.750 76.710 ;
        RECT 81.470 75.910 81.750 76.190 ;
        RECT 82.790 76.430 83.070 76.710 ;
        RECT 82.790 75.910 83.070 76.190 ;
        RECT 84.110 76.430 84.390 76.710 ;
        RECT 84.110 75.910 84.390 76.190 ;
        RECT 85.430 76.430 85.710 76.710 ;
        RECT 85.430 75.910 85.710 76.190 ;
        RECT 86.750 82.470 87.030 82.750 ;
        RECT 86.750 81.950 87.030 82.230 ;
        RECT 88.070 82.470 88.350 82.750 ;
        RECT 88.070 81.950 88.350 82.230 ;
        RECT 89.390 85.490 89.670 85.770 ;
        RECT 89.390 84.970 89.670 85.250 ;
        RECT 90.710 73.410 90.990 73.690 ;
        RECT 90.710 72.890 90.990 73.170 ;
        RECT 92.030 79.450 92.310 79.730 ;
        RECT 92.030 78.930 92.310 79.210 ;
        RECT 93.350 85.490 93.630 85.770 ;
        RECT 93.350 84.970 93.630 85.250 ;
        RECT 94.670 82.470 94.950 82.750 ;
        RECT 94.670 81.950 94.950 82.230 ;
        RECT 95.990 82.470 96.270 82.750 ;
        RECT 95.990 81.950 96.270 82.230 ;
        RECT 97.310 76.430 97.590 76.710 ;
        RECT 97.310 75.910 97.590 76.190 ;
        RECT 98.630 76.430 98.910 76.710 ;
        RECT 98.630 75.910 98.910 76.190 ;
        RECT 99.950 76.430 100.230 76.710 ;
        RECT 99.950 75.910 100.230 76.190 ;
        RECT 101.270 76.430 101.550 76.710 ;
        RECT 101.270 75.910 101.550 76.190 ;
        RECT 102.590 76.430 102.870 76.710 ;
        RECT 102.590 75.910 102.870 76.190 ;
        RECT 103.910 76.430 104.190 76.710 ;
        RECT 103.910 75.910 104.190 76.190 ;
        RECT 105.230 76.430 105.510 76.710 ;
        RECT 105.230 75.910 105.510 76.190 ;
        RECT 106.550 76.430 106.830 76.710 ;
        RECT 106.550 75.910 106.830 76.190 ;
        RECT 107.870 82.470 108.150 82.750 ;
        RECT 107.870 81.950 108.150 82.230 ;
        RECT 109.190 82.470 109.470 82.750 ;
        RECT 109.190 81.950 109.470 82.230 ;
        RECT 110.510 85.490 110.790 85.770 ;
        RECT 110.510 84.970 110.790 85.250 ;
        RECT 111.830 79.450 112.110 79.730 ;
        RECT 111.830 78.930 112.110 79.210 ;
        RECT 113.150 88.510 113.430 88.790 ;
        RECT 113.150 87.990 113.430 88.270 ;
        RECT 114.470 85.490 114.750 85.770 ;
        RECT 114.470 84.970 114.750 85.250 ;
        RECT 115.790 82.470 116.070 82.750 ;
        RECT 115.790 81.950 116.070 82.230 ;
        RECT 117.110 82.470 117.390 82.750 ;
        RECT 117.110 81.950 117.390 82.230 ;
        RECT 118.430 76.430 118.710 76.710 ;
        RECT 118.430 75.910 118.710 76.190 ;
        RECT 119.750 76.430 120.030 76.710 ;
        RECT 119.750 75.910 120.030 76.190 ;
        RECT 121.070 76.430 121.350 76.710 ;
        RECT 121.070 75.910 121.350 76.190 ;
        RECT 122.390 76.430 122.670 76.710 ;
        RECT 122.390 75.910 122.670 76.190 ;
        RECT 123.710 80.500 123.990 80.780 ;
        RECT 123.710 79.980 123.990 80.260 ;
        RECT 79.280 71.250 79.560 71.530 ;
        RECT 79.800 71.250 80.080 71.530 ;
        RECT 79.280 68.230 79.560 68.510 ;
        RECT 79.800 68.230 80.080 68.510 ;
        RECT 79.280 65.210 79.560 65.490 ;
        RECT 79.800 65.210 80.080 65.490 ;
        RECT 79.280 62.190 79.560 62.470 ;
        RECT 79.800 62.190 80.080 62.470 ;
        RECT 79.280 59.170 79.560 59.450 ;
        RECT 79.800 59.170 80.080 59.450 ;
        RECT 81.470 59.430 81.750 59.710 ;
        RECT 81.470 58.910 81.750 59.190 ;
        RECT 77.110 54.510 77.390 54.790 ;
        RECT 82.790 59.430 83.070 59.710 ;
        RECT 82.790 58.910 83.070 59.190 ;
        RECT 84.110 59.430 84.390 59.710 ;
        RECT 84.110 58.910 84.390 59.190 ;
        RECT 85.430 59.430 85.710 59.710 ;
        RECT 85.430 58.910 85.710 59.190 ;
        RECT 86.750 65.470 87.030 65.750 ;
        RECT 86.750 64.950 87.030 65.230 ;
        RECT 88.070 65.470 88.350 65.750 ;
        RECT 88.070 64.950 88.350 65.230 ;
        RECT 89.390 68.490 89.670 68.770 ;
        RECT 89.390 67.970 89.670 68.250 ;
        RECT 90.710 56.410 90.990 56.690 ;
        RECT 90.710 55.890 90.990 56.170 ;
        RECT 92.030 62.450 92.310 62.730 ;
        RECT 92.030 61.930 92.310 62.210 ;
        RECT 93.350 68.490 93.630 68.770 ;
        RECT 93.350 67.970 93.630 68.250 ;
        RECT 94.670 65.470 94.950 65.750 ;
        RECT 94.670 64.950 94.950 65.230 ;
        RECT 95.990 65.470 96.270 65.750 ;
        RECT 95.990 64.950 96.270 65.230 ;
        RECT 97.310 59.430 97.590 59.710 ;
        RECT 97.310 58.910 97.590 59.190 ;
        RECT 98.630 59.430 98.910 59.710 ;
        RECT 98.630 58.910 98.910 59.190 ;
        RECT 99.950 59.430 100.230 59.710 ;
        RECT 99.950 58.910 100.230 59.190 ;
        RECT 101.270 59.430 101.550 59.710 ;
        RECT 101.270 58.910 101.550 59.190 ;
        RECT 102.590 59.430 102.870 59.710 ;
        RECT 102.590 58.910 102.870 59.190 ;
        RECT 103.910 59.430 104.190 59.710 ;
        RECT 103.910 58.910 104.190 59.190 ;
        RECT 105.230 59.430 105.510 59.710 ;
        RECT 105.230 58.910 105.510 59.190 ;
        RECT 106.550 59.430 106.830 59.710 ;
        RECT 106.550 58.910 106.830 59.190 ;
        RECT 107.870 65.470 108.150 65.750 ;
        RECT 107.870 64.950 108.150 65.230 ;
        RECT 109.190 65.470 109.470 65.750 ;
        RECT 109.190 64.950 109.470 65.230 ;
        RECT 110.510 68.490 110.790 68.770 ;
        RECT 110.510 67.970 110.790 68.250 ;
        RECT 111.830 62.450 112.110 62.730 ;
        RECT 111.830 61.930 112.110 62.210 ;
        RECT 113.150 71.510 113.430 71.790 ;
        RECT 113.150 70.990 113.430 71.270 ;
        RECT 114.470 68.490 114.750 68.770 ;
        RECT 114.470 67.970 114.750 68.250 ;
        RECT 115.790 65.470 116.070 65.750 ;
        RECT 115.790 64.950 116.070 65.230 ;
        RECT 117.110 65.470 117.390 65.750 ;
        RECT 117.110 64.950 117.390 65.230 ;
        RECT 118.430 59.430 118.710 59.710 ;
        RECT 118.430 58.910 118.710 59.190 ;
        RECT 119.750 59.430 120.030 59.710 ;
        RECT 119.750 58.910 120.030 59.190 ;
        RECT 121.070 59.430 121.350 59.710 ;
        RECT 121.070 58.910 121.350 59.190 ;
        RECT 122.390 59.430 122.670 59.710 ;
        RECT 122.390 58.910 122.670 59.190 ;
        RECT 123.710 63.500 123.990 63.780 ;
        RECT 123.710 62.980 123.990 63.260 ;
        RECT 77.110 53.990 77.390 54.270 ;
        RECT 79.280 54.250 79.560 54.530 ;
        RECT 79.800 54.250 80.080 54.530 ;
        RECT 77.110 51.490 77.390 51.770 ;
        RECT 77.110 50.970 77.390 51.250 ;
        RECT 79.280 51.230 79.560 51.510 ;
        RECT 79.800 51.230 80.080 51.510 ;
        RECT 77.110 48.470 77.390 48.750 ;
        RECT 77.110 47.950 77.390 48.230 ;
        RECT 79.280 48.210 79.560 48.490 ;
        RECT 79.800 48.210 80.080 48.490 ;
        RECT 77.110 45.450 77.390 45.730 ;
        RECT 77.110 44.930 77.390 45.210 ;
        RECT 79.280 45.190 79.560 45.470 ;
        RECT 79.800 45.190 80.080 45.470 ;
        RECT 77.110 42.430 77.390 42.710 ;
        RECT 77.110 41.910 77.390 42.190 ;
        RECT 79.280 42.170 79.560 42.450 ;
        RECT 79.800 42.170 80.080 42.450 ;
        RECT 77.110 39.410 77.390 39.690 ;
        RECT 77.110 38.890 77.390 39.170 ;
        RECT 79.280 39.150 79.560 39.430 ;
        RECT 79.800 39.150 80.080 39.430 ;
        RECT 81.470 42.430 81.750 42.710 ;
        RECT 81.470 41.910 81.750 42.190 ;
        RECT 82.790 42.430 83.070 42.710 ;
        RECT 82.790 41.910 83.070 42.190 ;
        RECT 84.110 42.430 84.390 42.710 ;
        RECT 84.110 41.910 84.390 42.190 ;
        RECT 85.430 42.430 85.710 42.710 ;
        RECT 85.430 41.910 85.710 42.190 ;
        RECT 86.750 48.470 87.030 48.750 ;
        RECT 86.750 47.950 87.030 48.230 ;
        RECT 88.070 48.470 88.350 48.750 ;
        RECT 88.070 47.950 88.350 48.230 ;
        RECT 89.390 51.490 89.670 51.770 ;
        RECT 89.390 50.970 89.670 51.250 ;
        RECT 90.710 39.410 90.990 39.690 ;
        RECT 90.710 38.890 90.990 39.170 ;
        RECT 92.030 45.450 92.310 45.730 ;
        RECT 92.030 44.930 92.310 45.210 ;
        RECT 93.350 51.490 93.630 51.770 ;
        RECT 93.350 50.970 93.630 51.250 ;
        RECT 94.670 48.470 94.950 48.750 ;
        RECT 94.670 47.950 94.950 48.230 ;
        RECT 95.990 48.470 96.270 48.750 ;
        RECT 95.990 47.950 96.270 48.230 ;
        RECT 97.310 42.430 97.590 42.710 ;
        RECT 97.310 41.910 97.590 42.190 ;
        RECT 98.630 42.430 98.910 42.710 ;
        RECT 98.630 41.910 98.910 42.190 ;
        RECT 99.950 42.430 100.230 42.710 ;
        RECT 99.950 41.910 100.230 42.190 ;
        RECT 101.270 42.430 101.550 42.710 ;
        RECT 101.270 41.910 101.550 42.190 ;
        RECT 102.590 42.430 102.870 42.710 ;
        RECT 102.590 41.910 102.870 42.190 ;
        RECT 103.910 42.430 104.190 42.710 ;
        RECT 103.910 41.910 104.190 42.190 ;
        RECT 105.230 42.430 105.510 42.710 ;
        RECT 105.230 41.910 105.510 42.190 ;
        RECT 106.550 42.430 106.830 42.710 ;
        RECT 106.550 41.910 106.830 42.190 ;
        RECT 107.870 48.470 108.150 48.750 ;
        RECT 107.870 47.950 108.150 48.230 ;
        RECT 109.190 48.470 109.470 48.750 ;
        RECT 109.190 47.950 109.470 48.230 ;
        RECT 110.510 51.490 110.790 51.770 ;
        RECT 110.510 50.970 110.790 51.250 ;
        RECT 111.830 45.450 112.110 45.730 ;
        RECT 111.830 44.930 112.110 45.210 ;
        RECT 113.150 54.510 113.430 54.790 ;
        RECT 113.150 53.990 113.430 54.270 ;
        RECT 114.470 51.490 114.750 51.770 ;
        RECT 114.470 50.970 114.750 51.250 ;
        RECT 115.790 48.470 116.070 48.750 ;
        RECT 115.790 47.950 116.070 48.230 ;
        RECT 117.110 48.470 117.390 48.750 ;
        RECT 117.110 47.950 117.390 48.230 ;
        RECT 118.430 42.430 118.710 42.710 ;
        RECT 118.430 41.910 118.710 42.190 ;
        RECT 119.750 42.430 120.030 42.710 ;
        RECT 119.750 41.910 120.030 42.190 ;
        RECT 121.070 42.430 121.350 42.710 ;
        RECT 121.070 41.910 121.350 42.190 ;
        RECT 122.390 42.430 122.670 42.710 ;
        RECT 122.390 41.910 122.670 42.190 ;
        RECT 123.710 46.500 123.990 46.780 ;
        RECT 123.710 45.980 123.990 46.260 ;
        RECT 44.550 36.280 45.630 36.600 ;
        RECT 11.790 35.480 12.870 35.800 ;
        RECT 44.550 34.680 45.630 35.000 ;
        RECT 11.790 33.880 12.870 34.200 ;
        RECT 44.550 33.080 45.630 33.400 ;
        RECT 90.630 36.280 91.710 36.600 ;
        RECT 123.390 35.480 124.470 35.800 ;
        RECT 90.630 34.680 91.710 35.000 ;
        RECT 123.390 33.880 124.470 34.200 ;
        RECT 90.630 33.080 91.710 33.400 ;
        RECT 11.790 32.280 12.870 32.600 ;
        RECT 123.390 32.280 124.470 32.600 ;
        RECT 44.550 31.480 45.630 31.800 ;
        RECT 11.790 30.680 12.870 31.000 ;
        RECT 44.550 29.880 45.630 30.200 ;
        RECT 11.790 29.080 12.870 29.400 ;
        RECT 90.630 31.480 91.710 31.800 ;
        RECT 123.390 30.680 124.470 31.000 ;
        RECT 90.630 29.880 91.710 30.200 ;
        RECT 52.330 29.380 52.610 29.660 ;
        RECT 52.850 29.380 53.130 29.660 ;
        RECT 56.290 29.380 56.570 29.660 ;
        RECT 56.810 29.380 57.090 29.660 ;
        RECT 79.170 29.380 79.450 29.660 ;
        RECT 79.690 29.380 79.970 29.660 ;
        RECT 83.130 29.380 83.410 29.660 ;
        RECT 83.650 29.380 83.930 29.660 ;
        RECT 44.550 28.280 45.630 28.600 ;
        RECT 52.330 28.500 52.610 28.780 ;
        RECT 52.850 28.500 53.130 28.780 ;
        RECT 56.290 28.500 56.570 28.780 ;
        RECT 56.810 28.500 57.090 28.780 ;
        RECT 79.170 28.500 79.450 28.780 ;
        RECT 79.690 28.500 79.970 28.780 ;
        RECT 83.130 28.500 83.410 28.780 ;
        RECT 83.650 28.500 83.930 28.780 ;
        RECT 123.390 29.080 124.470 29.400 ;
        RECT 90.630 28.280 91.710 28.600 ;
        RECT 11.790 27.480 12.870 27.800 ;
        RECT 58.890 27.620 59.170 27.900 ;
        RECT 59.410 27.620 59.690 27.900 ;
        RECT 44.550 26.680 45.630 27.000 ;
        RECT 52.330 26.740 52.610 27.020 ;
        RECT 52.850 26.740 53.130 27.020 ;
        RECT 56.290 26.740 56.570 27.020 ;
        RECT 56.810 26.740 57.090 27.020 ;
        RECT 11.790 25.880 12.870 26.200 ;
        RECT 76.570 27.620 76.850 27.900 ;
        RECT 77.090 27.620 77.370 27.900 ;
        RECT 123.390 27.480 124.470 27.800 ;
        RECT 79.170 26.740 79.450 27.020 ;
        RECT 79.690 26.740 79.970 27.020 ;
        RECT 83.130 26.740 83.410 27.020 ;
        RECT 83.650 26.740 83.930 27.020 ;
        RECT 90.630 26.680 91.710 27.000 ;
        RECT 52.330 25.860 52.610 26.140 ;
        RECT 52.850 25.860 53.130 26.140 ;
        RECT 56.290 25.860 56.570 26.140 ;
        RECT 56.810 25.860 57.090 26.140 ;
        RECT 63.330 25.860 63.610 26.140 ;
        RECT 63.850 25.860 64.130 26.140 ;
        RECT 71.970 25.860 72.250 26.140 ;
        RECT 72.490 25.860 72.770 26.140 ;
        RECT 79.170 25.860 79.450 26.140 ;
        RECT 79.690 25.860 79.970 26.140 ;
        RECT 83.130 25.860 83.410 26.140 ;
        RECT 83.650 25.860 83.930 26.140 ;
        RECT 44.550 25.080 45.630 25.400 ;
        RECT 123.390 25.880 124.470 26.200 ;
        RECT 11.790 24.280 12.870 24.600 ;
        RECT 52.330 24.980 52.610 25.260 ;
        RECT 52.850 24.980 53.130 25.260 ;
        RECT 56.290 24.980 56.570 25.260 ;
        RECT 56.810 24.980 57.090 25.260 ;
        RECT 79.170 24.980 79.450 25.260 ;
        RECT 79.690 24.980 79.970 25.260 ;
        RECT 83.130 24.980 83.410 25.260 ;
        RECT 83.650 24.980 83.930 25.260 ;
        RECT 90.630 25.080 91.710 25.400 ;
        RECT 44.550 23.480 45.630 23.800 ;
        RECT 52.330 23.220 52.610 23.500 ;
        RECT 52.850 23.220 53.130 23.500 ;
        RECT 56.290 23.220 56.570 23.500 ;
        RECT 56.810 23.220 57.090 23.500 ;
        RECT 11.790 22.680 12.870 23.000 ;
        RECT 52.330 22.340 52.610 22.620 ;
        RECT 52.850 22.340 53.130 22.620 ;
        RECT 56.130 22.340 56.410 22.620 ;
        RECT 56.650 22.340 56.930 22.620 ;
        RECT 44.550 21.880 45.630 22.200 ;
        RECT 123.390 24.280 124.470 24.600 ;
        RECT 79.170 23.220 79.450 23.500 ;
        RECT 79.690 23.220 79.970 23.500 ;
        RECT 83.130 23.220 83.410 23.500 ;
        RECT 83.650 23.220 83.930 23.500 ;
        RECT 90.630 23.480 91.710 23.800 ;
        RECT 123.390 22.680 124.470 23.000 ;
        RECT 79.330 22.340 79.610 22.620 ;
        RECT 79.850 22.340 80.130 22.620 ;
        RECT 83.130 22.340 83.410 22.620 ;
        RECT 83.650 22.340 83.930 22.620 ;
        RECT 90.630 21.880 91.710 22.200 ;
        RECT 11.790 21.080 12.870 21.400 ;
        RECT 50.170 21.460 50.450 21.740 ;
        RECT 50.690 21.460 50.970 21.740 ;
        RECT 85.290 21.460 85.570 21.740 ;
        RECT 85.810 21.460 86.090 21.740 ;
        RECT 58.450 21.020 58.730 21.300 ;
        RECT 58.970 21.020 59.250 21.300 ;
        RECT 77.010 21.020 77.290 21.300 ;
        RECT 77.530 21.020 77.810 21.300 ;
        RECT 44.550 20.280 45.630 20.600 ;
        RECT 56.290 20.580 56.570 20.860 ;
        RECT 56.810 20.580 57.090 20.860 ;
        RECT 79.170 20.580 79.450 20.860 ;
        RECT 79.690 20.580 79.970 20.860 ;
        RECT 123.390 21.080 124.470 21.400 ;
        RECT 11.790 19.480 12.870 19.800 ;
        RECT 90.630 20.280 91.710 20.600 ;
        RECT 44.550 18.680 45.630 19.000 ;
        RECT 52.330 18.820 52.610 19.100 ;
        RECT 52.850 18.820 53.130 19.100 ;
        RECT 50.170 18.380 50.450 18.660 ;
        RECT 50.690 18.380 50.970 18.660 ;
        RECT 63.330 18.820 63.610 19.100 ;
        RECT 63.850 18.820 64.130 19.100 ;
        RECT 71.970 18.820 72.250 19.100 ;
        RECT 72.490 18.820 72.770 19.100 ;
        RECT 83.130 18.820 83.410 19.100 ;
        RECT 83.650 18.820 83.930 19.100 ;
        RECT 123.390 19.480 124.470 19.800 ;
        RECT 85.290 18.380 85.570 18.660 ;
        RECT 85.810 18.380 86.090 18.660 ;
        RECT 90.630 18.680 91.710 19.000 ;
        RECT 11.790 17.880 12.870 18.200 ;
        RECT 52.330 17.940 52.610 18.220 ;
        RECT 52.850 17.940 53.130 18.220 ;
        RECT 56.290 17.940 56.570 18.220 ;
        RECT 56.810 17.940 57.090 18.220 ;
        RECT 79.170 17.940 79.450 18.220 ;
        RECT 79.690 17.940 79.970 18.220 ;
        RECT 83.130 17.940 83.410 18.220 ;
        RECT 83.650 17.940 83.930 18.220 ;
        RECT 123.390 17.880 124.470 18.200 ;
        RECT 65.490 17.500 65.770 17.780 ;
        RECT 66.010 17.500 66.290 17.780 ;
        RECT 69.970 17.500 70.250 17.780 ;
        RECT 70.490 17.500 70.770 17.780 ;
        RECT 44.550 17.080 45.630 17.400 ;
        RECT 11.790 16.280 12.870 16.600 ;
        RECT 56.290 16.350 56.570 16.630 ;
        RECT 56.810 16.350 57.090 16.630 ;
        RECT 79.170 16.350 79.450 16.630 ;
        RECT 79.690 16.350 79.970 16.630 ;
        RECT 90.630 17.080 91.710 17.400 ;
        RECT 44.550 15.480 45.630 15.800 ;
        RECT 123.390 16.280 124.470 16.600 ;
        RECT 11.790 14.680 12.870 15.000 ;
        RECT 52.330 15.300 52.610 15.580 ;
        RECT 52.850 15.300 53.130 15.580 ;
        RECT 56.290 15.300 56.570 15.580 ;
        RECT 56.810 15.300 57.090 15.580 ;
        RECT 52.330 14.420 52.610 14.700 ;
        RECT 52.850 14.420 53.130 14.700 ;
        RECT 56.290 14.420 56.570 14.700 ;
        RECT 56.810 14.420 57.090 14.700 ;
        RECT 44.550 13.880 45.630 14.200 ;
        RECT 52.330 13.540 52.610 13.820 ;
        RECT 52.850 13.540 53.130 13.820 ;
        RECT 56.290 13.540 56.570 13.820 ;
        RECT 56.810 13.540 57.090 13.820 ;
        RECT 11.790 13.080 12.870 13.400 ;
        RECT 56.290 10.220 56.570 10.500 ;
        RECT 56.810 10.220 57.090 10.500 ;
        RECT 56.290 9.700 56.570 9.980 ;
        RECT 56.810 9.700 57.090 9.980 ;
        RECT 52.330 6.620 52.610 6.900 ;
        RECT 52.850 6.620 53.130 6.900 ;
        RECT 52.330 6.100 52.610 6.380 ;
        RECT 52.850 6.100 53.130 6.380 ;
        RECT 63.330 14.420 63.610 14.700 ;
        RECT 63.850 14.420 64.130 14.700 ;
        RECT 72.130 14.420 72.410 14.700 ;
        RECT 72.650 14.420 72.930 14.700 ;
        RECT 79.170 15.300 79.450 15.580 ;
        RECT 79.690 15.300 79.970 15.580 ;
        RECT 83.130 15.300 83.410 15.580 ;
        RECT 83.650 15.300 83.930 15.580 ;
        RECT 90.630 15.480 91.710 15.800 ;
        RECT 79.170 14.420 79.450 14.700 ;
        RECT 79.690 14.420 79.970 14.700 ;
        RECT 83.130 14.420 83.410 14.700 ;
        RECT 83.650 14.420 83.930 14.700 ;
        RECT 123.390 14.680 124.470 15.000 ;
        RECT 90.630 13.880 91.710 14.200 ;
        RECT 79.170 13.540 79.450 13.820 ;
        RECT 79.690 13.540 79.970 13.820 ;
        RECT 83.130 13.540 83.410 13.820 ;
        RECT 83.650 13.540 83.930 13.820 ;
        RECT 123.390 13.080 124.470 13.400 ;
        RECT 79.170 10.220 79.450 10.500 ;
        RECT 79.690 10.220 79.970 10.500 ;
        RECT 79.170 9.700 79.450 9.980 ;
        RECT 79.690 9.700 79.970 9.980 ;
        RECT 83.130 6.620 83.410 6.900 ;
        RECT 83.650 6.620 83.930 6.900 ;
        RECT 83.130 6.100 83.410 6.380 ;
        RECT 83.650 6.100 83.930 6.380 ;
        RECT 58.890 3.950 59.170 4.230 ;
        RECT 59.410 3.950 59.690 4.230 ;
        RECT 76.570 3.950 76.850 4.230 ;
        RECT 77.090 3.950 77.370 4.230 ;
      LAYER met2 ;
        RECT 57.470 224.275 57.905 224.685 ;
        RECT 59.695 224.665 59.995 224.675 ;
        RECT 59.660 224.385 60.030 224.665 ;
        RECT 15.750 221.810 16.050 223.900 ;
        RECT 35.965 223.570 36.355 223.780 ;
        RECT 40.860 223.750 41.140 223.785 ;
        RECT 35.965 223.480 37.120 223.570 ;
        RECT 36.010 223.270 37.120 223.480 ;
        RECT 32.360 222.250 32.640 222.285 ;
        RECT 32.350 221.810 32.650 222.250 ;
        RECT 40.850 221.810 41.150 223.750 ;
        RECT 57.505 223.650 57.805 224.275 ;
        RECT 59.695 223.990 59.995 224.385 ;
        RECT 61.180 224.160 61.975 224.460 ;
        RECT 86.890 224.440 87.170 224.475 ;
        RECT 57.505 223.350 59.400 223.650 ;
        RECT 59.100 223.045 59.400 223.350 ;
        RECT 57.560 222.950 57.840 222.985 ;
        RECT 57.550 221.810 57.850 222.950 ;
        RECT 59.100 222.745 79.725 223.045 ;
        RECT 82.660 222.950 82.940 222.985 ;
        RECT 66.060 222.250 66.340 222.285 ;
        RECT 66.050 221.810 66.350 222.250 ;
        RECT 15.310 221.470 16.390 221.810 ;
        RECT 31.870 221.470 32.950 221.810 ;
        RECT 40.510 221.470 41.590 221.810 ;
        RECT 57.070 221.470 58.150 221.810 ;
        RECT 65.710 221.470 66.790 221.810 ;
        RECT 79.425 221.695 79.725 222.745 ;
        RECT 82.650 221.810 82.950 222.950 ;
        RECT 86.880 222.380 87.180 224.440 ;
        RECT 108.060 224.140 108.340 224.440 ;
        RECT 91.250 223.540 91.550 223.550 ;
        RECT 91.215 223.260 91.585 223.540 ;
        RECT 91.250 221.810 91.550 223.260 ;
        RECT 108.050 221.810 108.350 224.140 ;
        RECT 111.330 223.310 112.310 223.320 ;
        RECT 111.295 223.030 112.310 223.310 ;
        RECT 111.330 223.020 112.310 223.030 ;
        RECT 116.490 222.740 116.790 224.140 ;
        RECT 116.490 222.380 116.800 222.740 ;
        RECT 116.490 221.810 116.790 222.380 ;
        RECT 82.270 221.470 83.350 221.810 ;
        RECT 90.910 221.470 91.990 221.810 ;
        RECT 107.470 221.470 108.550 221.810 ;
        RECT 116.110 221.470 117.190 221.810 ;
        RECT 15.680 220.660 16.020 221.470 ;
        RECT 32.240 220.660 32.580 221.470 ;
        RECT 40.880 220.660 41.220 221.470 ;
        RECT 57.440 220.660 57.780 221.470 ;
        RECT 66.080 220.660 66.420 221.470 ;
        RECT 82.640 220.660 82.980 221.470 ;
        RECT 91.280 220.660 91.620 221.470 ;
        RECT 107.840 220.660 108.180 221.470 ;
        RECT 116.190 221.200 117.110 221.470 ;
        RECT 15.390 220.320 16.310 220.660 ;
        RECT 31.950 220.320 32.870 220.660 ;
        RECT 40.590 220.320 41.510 220.660 ;
        RECT 57.150 220.320 58.070 220.660 ;
        RECT 65.790 220.320 66.710 220.660 ;
        RECT 82.350 220.320 83.270 220.660 ;
        RECT 90.990 220.320 91.910 220.660 ;
        RECT 107.550 220.320 108.470 220.660 ;
        RECT 116.110 220.320 117.030 220.660 ;
        RECT 120.070 220.320 120.990 220.660 ;
        RECT 15.310 219.440 16.230 219.780 ;
        RECT 19.270 219.440 20.190 219.780 ;
        RECT 28.070 219.440 28.990 219.780 ;
        RECT 32.030 219.440 32.950 219.780 ;
        RECT 40.510 219.440 41.430 219.780 ;
        RECT 44.470 219.440 45.390 219.780 ;
        RECT 53.270 219.440 54.190 219.780 ;
        RECT 57.230 219.440 58.150 219.780 ;
        RECT 65.710 219.440 66.630 219.780 ;
        RECT 69.670 219.440 70.590 219.780 ;
        RECT 78.470 219.440 79.390 219.780 ;
        RECT 82.430 219.440 83.350 219.780 ;
        RECT 90.910 219.440 91.830 219.780 ;
        RECT 94.870 219.440 95.790 219.780 ;
        RECT 103.670 219.440 104.590 219.780 ;
        RECT 107.630 219.440 108.550 219.780 ;
        RECT 116.110 219.770 124.930 219.780 ;
        RECT 132.530 219.770 132.870 219.800 ;
        RECT 116.110 219.440 132.870 219.770 ;
        RECT 123.730 219.430 132.870 219.440 ;
        RECT 132.530 219.400 132.870 219.430 ;
        RECT 116.110 218.560 117.030 218.900 ;
        RECT 120.070 218.560 120.990 218.900 ;
        RECT 120.070 217.680 120.990 218.020 ;
        RECT 15.310 216.800 16.230 217.140 ;
        RECT 19.270 216.800 20.190 217.140 ;
        RECT 28.070 216.800 28.990 217.140 ;
        RECT 32.030 216.800 32.950 217.140 ;
        RECT 40.510 216.800 41.430 217.140 ;
        RECT 44.470 216.800 45.390 217.140 ;
        RECT 53.270 216.800 54.190 217.140 ;
        RECT 57.230 216.800 58.150 217.140 ;
        RECT 65.710 216.800 66.630 217.140 ;
        RECT 69.670 216.800 70.590 217.140 ;
        RECT 78.470 216.800 79.390 217.140 ;
        RECT 82.430 216.800 83.350 217.140 ;
        RECT 90.910 216.800 91.830 217.140 ;
        RECT 94.870 216.800 95.790 217.140 ;
        RECT 103.670 216.800 104.590 217.140 ;
        RECT 107.630 216.800 108.550 217.140 ;
        RECT 113.310 216.360 115.030 216.700 ;
        RECT 15.310 214.160 16.230 214.500 ;
        RECT 19.270 214.160 20.190 214.500 ;
        RECT 28.070 214.160 28.990 214.500 ;
        RECT 32.030 214.160 32.950 214.500 ;
        RECT 40.510 214.160 41.430 214.500 ;
        RECT 44.470 214.160 45.390 214.500 ;
        RECT 53.270 214.160 54.190 214.500 ;
        RECT 57.230 214.160 58.150 214.500 ;
        RECT 65.710 214.160 66.630 214.500 ;
        RECT 69.670 214.160 70.590 214.500 ;
        RECT 78.470 214.160 79.390 214.500 ;
        RECT 82.430 214.160 83.350 214.500 ;
        RECT 90.910 214.160 91.830 214.500 ;
        RECT 94.870 214.160 95.790 214.500 ;
        RECT 103.670 214.160 104.590 214.500 ;
        RECT 107.630 214.160 108.550 214.500 ;
        RECT 15.310 212.400 16.230 212.740 ;
        RECT 19.270 212.400 20.190 212.740 ;
        RECT 28.070 212.400 28.990 212.740 ;
        RECT 32.030 212.400 32.950 212.740 ;
        RECT 40.510 212.400 41.430 212.740 ;
        RECT 44.470 212.400 45.390 212.740 ;
        RECT 53.270 212.400 54.190 212.740 ;
        RECT 57.230 212.400 58.150 212.740 ;
        RECT 65.710 212.400 66.630 212.740 ;
        RECT 69.670 212.400 70.590 212.740 ;
        RECT 78.470 212.400 79.390 212.740 ;
        RECT 82.430 212.400 83.350 212.740 ;
        RECT 90.910 212.400 91.830 212.740 ;
        RECT 94.870 212.400 95.790 212.740 ;
        RECT 103.670 212.400 104.590 212.740 ;
        RECT 107.630 212.400 108.550 212.740 ;
        RECT 113.310 210.540 113.650 216.360 ;
        RECT 116.110 215.920 117.030 216.260 ;
        RECT 120.070 215.920 120.990 216.260 ;
        RECT 116.110 215.370 124.930 215.380 ;
        RECT 116.110 215.345 131.070 215.370 ;
        RECT 116.110 215.055 131.090 215.345 ;
        RECT 116.110 215.040 131.070 215.055 ;
        RECT 124.230 215.030 131.070 215.040 ;
        RECT 116.110 214.160 117.030 214.500 ;
        RECT 120.070 214.160 120.990 214.500 ;
        RECT 116.110 213.570 124.930 213.620 ;
        RECT 116.110 213.280 127.080 213.570 ;
        RECT 124.230 213.230 127.080 213.280 ;
        RECT 116.110 212.400 117.030 212.740 ;
        RECT 120.070 212.400 120.990 212.740 ;
        RECT 116.110 211.520 117.030 211.860 ;
        RECT 113.310 210.200 115.030 210.540 ;
        RECT 15.310 209.760 16.230 210.100 ;
        RECT 19.270 209.760 20.190 210.100 ;
        RECT 28.070 209.760 28.990 210.100 ;
        RECT 32.030 209.760 32.950 210.100 ;
        RECT 40.510 209.760 41.430 210.100 ;
        RECT 44.470 209.760 45.390 210.100 ;
        RECT 53.270 209.760 54.190 210.100 ;
        RECT 57.230 209.760 58.150 210.100 ;
        RECT 65.710 209.760 66.630 210.100 ;
        RECT 69.670 209.760 70.590 210.100 ;
        RECT 78.470 209.760 79.390 210.100 ;
        RECT 82.430 209.760 83.350 210.100 ;
        RECT 90.910 209.760 91.830 210.100 ;
        RECT 94.870 209.760 95.790 210.100 ;
        RECT 103.670 209.760 104.590 210.100 ;
        RECT 107.630 209.760 108.550 210.100 ;
        RECT 113.310 209.220 113.650 210.200 ;
        RECT 116.110 209.760 117.030 210.100 ;
        RECT 120.070 209.760 120.990 210.100 ;
        RECT 113.310 208.880 117.190 209.220 ;
        RECT 116.110 208.000 117.030 208.340 ;
        RECT 120.070 208.000 120.990 208.340 ;
        RECT 13.230 207.560 14.150 207.900 ;
        RECT 34.110 207.560 35.030 207.900 ;
        RECT 38.430 207.560 39.350 207.900 ;
        RECT 59.310 207.560 60.230 207.900 ;
        RECT 63.630 207.560 64.550 207.900 ;
        RECT 84.510 207.560 85.430 207.900 ;
        RECT 88.830 207.560 89.750 207.900 ;
        RECT 109.710 207.560 110.630 207.900 ;
        RECT 113.950 207.560 114.870 207.900 ;
        RECT 13.520 197.995 13.860 207.560 ;
        RECT 15.310 207.120 16.230 207.460 ;
        RECT 19.270 207.120 20.190 207.460 ;
        RECT 28.070 207.120 28.990 207.460 ;
        RECT 32.030 207.120 32.950 207.460 ;
        RECT 15.310 205.360 16.230 205.700 ;
        RECT 19.270 205.360 20.190 205.700 ;
        RECT 28.070 205.360 28.990 205.700 ;
        RECT 32.030 205.360 32.950 205.700 ;
        RECT 15.310 203.600 16.230 203.940 ;
        RECT 19.270 203.600 20.190 203.940 ;
        RECT 28.070 203.600 28.990 203.940 ;
        RECT 32.030 203.600 32.950 203.940 ;
        RECT 15.310 202.720 16.230 203.060 ;
        RECT 19.270 202.720 20.190 203.060 ;
        RECT 28.070 202.720 28.990 203.060 ;
        RECT 32.030 202.720 32.950 203.060 ;
        RECT 15.310 201.840 16.230 202.180 ;
        RECT 19.270 201.840 20.190 202.180 ;
        RECT 28.070 201.840 28.990 202.180 ;
        RECT 32.030 201.840 32.950 202.180 ;
        RECT 15.310 199.070 16.230 199.990 ;
        RECT 32.030 199.070 32.950 199.990 ;
        RECT 13.230 197.975 13.860 197.995 ;
        RECT 13.205 197.970 13.975 197.975 ;
        RECT 13.150 197.630 14.230 197.970 ;
        RECT 19.270 197.630 20.190 198.550 ;
        RECT 22.050 197.630 22.970 198.550 ;
        RECT 25.090 197.630 26.010 198.550 ;
        RECT 28.070 197.630 28.990 198.550 ;
        RECT 34.400 197.970 34.740 207.560 ;
        RECT 38.720 198.370 39.060 207.560 ;
        RECT 40.510 207.120 41.430 207.460 ;
        RECT 44.470 207.120 45.390 207.460 ;
        RECT 53.270 207.120 54.190 207.460 ;
        RECT 57.230 207.120 58.150 207.460 ;
        RECT 40.510 205.360 41.430 205.700 ;
        RECT 44.470 205.360 45.390 205.700 ;
        RECT 53.270 205.360 54.190 205.700 ;
        RECT 57.230 205.360 58.150 205.700 ;
        RECT 40.510 203.600 41.430 203.940 ;
        RECT 44.470 203.600 45.390 203.940 ;
        RECT 53.270 203.600 54.190 203.940 ;
        RECT 57.230 203.600 58.150 203.940 ;
        RECT 40.510 202.720 41.430 203.060 ;
        RECT 44.470 202.720 45.390 203.060 ;
        RECT 53.270 202.720 54.190 203.060 ;
        RECT 57.230 202.720 58.150 203.060 ;
        RECT 40.510 201.840 41.430 202.180 ;
        RECT 44.470 201.840 45.390 202.180 ;
        RECT 53.270 201.840 54.190 202.180 ;
        RECT 57.230 201.840 58.150 202.180 ;
        RECT 40.510 199.070 41.430 199.990 ;
        RECT 57.230 199.070 58.150 199.990 ;
        RECT 38.720 197.970 39.170 198.370 ;
        RECT 34.030 197.630 35.110 197.970 ;
        RECT 38.350 197.630 39.430 197.970 ;
        RECT 44.470 197.630 45.390 198.550 ;
        RECT 47.250 197.630 48.170 198.550 ;
        RECT 50.290 197.630 51.210 198.550 ;
        RECT 53.270 197.630 54.190 198.550 ;
        RECT 59.600 198.045 59.940 207.560 ;
        RECT 63.920 198.045 64.260 207.560 ;
        RECT 65.710 207.120 66.630 207.460 ;
        RECT 69.670 207.120 70.590 207.460 ;
        RECT 78.470 207.120 79.390 207.460 ;
        RECT 82.430 207.120 83.350 207.460 ;
        RECT 65.710 205.360 66.630 205.700 ;
        RECT 69.670 205.360 70.590 205.700 ;
        RECT 78.470 205.360 79.390 205.700 ;
        RECT 82.430 205.360 83.350 205.700 ;
        RECT 65.710 203.600 66.630 203.940 ;
        RECT 69.670 203.600 70.590 203.940 ;
        RECT 78.470 203.600 79.390 203.940 ;
        RECT 82.430 203.600 83.350 203.940 ;
        RECT 65.710 202.720 66.630 203.060 ;
        RECT 69.670 202.720 70.590 203.060 ;
        RECT 78.470 202.720 79.390 203.060 ;
        RECT 82.430 202.720 83.350 203.060 ;
        RECT 65.710 201.840 66.630 202.180 ;
        RECT 69.670 201.840 70.590 202.180 ;
        RECT 78.470 201.840 79.390 202.180 ;
        RECT 82.430 201.840 83.350 202.180 ;
        RECT 65.710 199.070 66.630 199.990 ;
        RECT 82.430 199.070 83.350 199.990 ;
        RECT 59.600 197.970 59.990 198.045 ;
        RECT 63.910 197.970 64.290 198.045 ;
        RECT 59.230 197.630 60.310 197.970 ;
        RECT 63.550 197.630 64.630 197.970 ;
        RECT 69.670 197.630 70.590 198.550 ;
        RECT 72.450 197.630 73.370 198.550 ;
        RECT 75.490 197.630 76.410 198.550 ;
        RECT 78.470 197.630 79.390 198.550 ;
        RECT 84.800 198.045 85.140 207.560 ;
        RECT 89.120 198.045 89.460 207.560 ;
        RECT 90.910 207.120 91.830 207.460 ;
        RECT 94.870 207.120 95.790 207.460 ;
        RECT 103.670 207.120 104.590 207.460 ;
        RECT 107.630 207.120 108.550 207.460 ;
        RECT 90.910 205.360 91.830 205.700 ;
        RECT 94.870 205.360 95.790 205.700 ;
        RECT 103.670 205.360 104.590 205.700 ;
        RECT 107.630 205.360 108.550 205.700 ;
        RECT 90.910 203.600 91.830 203.940 ;
        RECT 94.870 203.600 95.790 203.940 ;
        RECT 103.670 203.600 104.590 203.940 ;
        RECT 107.630 203.600 108.550 203.940 ;
        RECT 90.910 202.720 91.830 203.060 ;
        RECT 94.870 202.720 95.790 203.060 ;
        RECT 103.670 202.720 104.590 203.060 ;
        RECT 107.630 202.720 108.550 203.060 ;
        RECT 90.910 201.840 91.830 202.180 ;
        RECT 94.870 201.840 95.790 202.180 ;
        RECT 103.670 201.840 104.590 202.180 ;
        RECT 107.630 201.840 108.550 202.180 ;
        RECT 90.910 199.070 91.830 199.990 ;
        RECT 107.630 199.070 108.550 199.990 ;
        RECT 84.710 197.970 85.140 198.045 ;
        RECT 89.110 197.970 89.490 198.045 ;
        RECT 84.430 197.630 85.510 197.970 ;
        RECT 88.750 197.630 89.830 197.970 ;
        RECT 94.870 197.630 95.790 198.550 ;
        RECT 97.650 197.630 98.570 198.550 ;
        RECT 100.690 197.630 101.610 198.550 ;
        RECT 103.670 197.630 104.590 198.550 ;
        RECT 110.000 197.970 110.340 207.560 ;
        RECT 140.035 206.315 141.035 206.695 ;
        RECT 143.995 206.315 144.995 206.695 ;
        RECT 116.110 205.360 117.030 205.700 ;
        RECT 120.070 205.360 120.990 205.700 ;
        RECT 140.035 205.435 141.035 205.815 ;
        RECT 143.995 205.435 144.995 205.815 ;
        RECT 114.110 204.040 115.030 204.380 ;
        RECT 116.110 203.600 117.030 203.940 ;
        RECT 120.070 203.600 120.990 203.940 ;
        RECT 140.035 203.675 141.035 204.055 ;
        RECT 143.995 203.675 144.995 204.055 ;
        RECT 116.110 202.720 117.030 203.060 ;
        RECT 120.070 202.720 120.990 203.060 ;
        RECT 116.110 201.840 117.030 202.180 ;
        RECT 120.070 201.840 120.990 202.180 ;
        RECT 140.035 201.915 141.035 202.295 ;
        RECT 143.995 201.915 144.995 202.295 ;
        RECT 140.035 201.035 141.035 201.415 ;
        RECT 143.995 201.035 144.995 201.415 ;
        RECT 111.830 199.445 112.170 200.200 ;
        RECT 111.810 199.155 112.190 199.445 ;
        RECT 111.830 199.130 112.170 199.155 ;
        RECT 116.110 199.070 117.030 199.990 ;
        RECT 109.630 197.630 110.710 197.970 ;
        RECT 120.070 197.630 120.990 198.550 ;
        RECT 13.205 197.625 13.975 197.630 ;
        RECT 13.230 197.605 13.530 197.625 ;
        RECT 38.810 197.555 39.190 197.630 ;
        RECT 38.830 197.530 39.170 197.555 ;
        RECT 114.255 197.070 114.545 197.090 ;
        RECT 114.230 196.730 147.915 197.070 ;
        RECT 114.255 196.710 114.545 196.730 ;
        RECT 102.575 196.070 102.865 196.090 ;
        RECT 102.550 195.730 131.115 196.070 ;
        RECT 102.575 195.710 102.865 195.730 ;
        RECT 41.885 195.570 42.175 195.590 ;
        RECT 30.830 195.230 34.715 195.570 ;
        RECT 38.785 195.230 42.200 195.570 ;
        RECT 81.385 195.545 85.070 195.570 ;
        RECT 56.280 195.470 56.570 195.490 ;
        RECT 59.630 195.470 59.970 195.515 ;
        RECT 41.885 195.210 42.175 195.230 ;
        RECT 56.255 195.130 59.970 195.470 ;
        RECT 63.885 195.445 67.400 195.470 ;
        RECT 63.885 195.155 67.420 195.445 ;
        RECT 81.385 195.255 85.090 195.545 ;
        RECT 89.130 195.470 89.470 195.515 ;
        RECT 89.130 195.445 92.600 195.470 ;
        RECT 81.385 195.230 85.070 195.255 ;
        RECT 89.130 195.155 92.620 195.445 ;
        RECT 63.885 195.130 67.400 195.155 ;
        RECT 89.130 195.130 92.600 195.155 ;
        RECT 56.280 195.110 56.570 195.130 ;
        RECT 59.630 195.085 59.970 195.130 ;
        RECT 89.130 195.085 89.470 195.130 ;
        RECT 19.170 194.030 20.090 194.950 ;
        RECT 27.970 194.030 28.890 194.950 ;
        RECT 44.370 194.030 45.290 194.950 ;
        RECT 53.170 194.030 54.090 194.950 ;
        RECT 69.570 194.030 70.490 194.950 ;
        RECT 78.370 194.030 79.290 194.950 ;
        RECT 94.770 194.030 95.690 194.950 ;
        RECT 103.570 194.030 104.490 194.950 ;
        RECT 119.970 194.030 120.890 194.950 ;
        RECT 15.210 190.430 16.130 191.350 ;
        RECT 31.930 190.430 32.850 191.350 ;
        RECT 40.410 190.430 41.330 191.350 ;
        RECT 57.130 190.430 58.050 191.350 ;
        RECT 65.610 190.430 66.530 191.350 ;
        RECT 82.330 190.430 83.250 191.350 ;
        RECT 90.810 190.430 91.730 191.350 ;
        RECT 107.530 190.430 108.450 191.350 ;
        RECT 116.010 190.430 116.930 191.350 ;
        RECT 15.210 187.140 16.130 187.480 ;
        RECT 19.170 187.140 20.090 187.480 ;
        RECT 27.970 187.140 28.890 187.480 ;
        RECT 31.930 187.140 32.850 187.480 ;
        RECT 40.410 187.140 41.330 187.480 ;
        RECT 44.370 187.140 45.290 187.480 ;
        RECT 53.170 187.140 54.090 187.480 ;
        RECT 57.130 187.140 58.050 187.480 ;
        RECT 65.610 187.140 66.530 187.480 ;
        RECT 69.570 187.140 70.490 187.480 ;
        RECT 78.370 187.140 79.290 187.480 ;
        RECT 82.330 187.140 83.250 187.480 ;
        RECT 90.810 187.140 91.730 187.480 ;
        RECT 94.770 187.140 95.690 187.480 ;
        RECT 103.570 187.140 104.490 187.480 ;
        RECT 107.530 187.140 108.450 187.480 ;
        RECT 15.210 186.260 16.130 186.600 ;
        RECT 19.170 186.260 20.090 186.600 ;
        RECT 27.970 186.260 28.890 186.600 ;
        RECT 31.930 186.260 32.850 186.600 ;
        RECT 40.410 186.260 41.330 186.600 ;
        RECT 44.370 186.260 45.290 186.600 ;
        RECT 53.170 186.260 54.090 186.600 ;
        RECT 57.130 186.260 58.050 186.600 ;
        RECT 65.610 186.260 66.530 186.600 ;
        RECT 69.570 186.260 70.490 186.600 ;
        RECT 78.370 186.260 79.290 186.600 ;
        RECT 82.330 186.260 83.250 186.600 ;
        RECT 90.810 186.260 91.730 186.600 ;
        RECT 94.770 186.260 95.690 186.600 ;
        RECT 103.570 186.260 104.490 186.600 ;
        RECT 107.530 186.260 108.450 186.600 ;
        RECT 19.170 185.550 21.190 185.890 ;
        RECT 44.370 185.550 46.390 185.890 ;
        RECT 69.570 185.550 71.590 185.890 ;
        RECT 94.770 185.550 96.790 185.890 ;
        RECT 15.210 184.500 16.130 184.840 ;
        RECT 19.170 184.500 20.090 184.840 ;
        RECT 15.210 183.620 16.130 183.960 ;
        RECT 20.850 182.880 21.190 185.550 ;
        RECT 27.970 184.500 28.890 184.840 ;
        RECT 31.930 184.500 32.850 184.840 ;
        RECT 40.410 184.500 41.330 184.840 ;
        RECT 44.370 184.500 45.290 184.840 ;
        RECT 31.930 183.620 32.850 183.960 ;
        RECT 40.410 183.620 41.330 183.960 ;
        RECT 33.590 183.180 34.850 183.520 ;
        RECT 33.590 182.880 33.930 183.180 ;
        RECT 20.850 182.540 33.930 182.880 ;
        RECT 46.050 182.880 46.390 185.550 ;
        RECT 53.170 184.500 54.090 184.840 ;
        RECT 57.130 184.500 58.050 184.840 ;
        RECT 65.610 184.500 66.530 184.840 ;
        RECT 69.570 184.500 70.490 184.840 ;
        RECT 57.130 183.620 58.050 183.960 ;
        RECT 65.610 183.620 66.530 183.960 ;
        RECT 58.790 183.180 60.050 183.520 ;
        RECT 58.790 182.880 59.130 183.180 ;
        RECT 46.050 182.540 59.130 182.880 ;
        RECT 71.250 182.880 71.590 185.550 ;
        RECT 78.370 184.500 79.290 184.840 ;
        RECT 82.330 184.500 83.250 184.840 ;
        RECT 90.810 184.500 91.730 184.840 ;
        RECT 94.770 184.500 95.690 184.840 ;
        RECT 82.330 183.620 83.250 183.960 ;
        RECT 90.810 183.620 91.730 183.960 ;
        RECT 83.990 183.180 85.250 183.520 ;
        RECT 83.990 182.880 84.330 183.180 ;
        RECT 71.250 182.540 84.330 182.880 ;
        RECT 96.450 182.880 96.790 185.550 ;
        RECT 103.410 185.380 111.910 185.720 ;
        RECT 103.570 184.500 104.490 184.840 ;
        RECT 107.530 184.500 108.450 184.840 ;
        RECT 107.530 183.620 108.450 183.960 ;
        RECT 109.190 183.180 110.450 183.520 ;
        RECT 109.190 182.880 109.530 183.180 ;
        RECT 96.450 182.540 109.530 182.880 ;
        RECT 15.210 181.860 16.130 182.200 ;
        RECT 19.170 181.860 20.090 182.200 ;
        RECT 27.970 181.860 28.890 182.200 ;
        RECT 31.930 181.860 32.850 182.200 ;
        RECT 40.410 181.860 41.330 182.200 ;
        RECT 44.370 181.860 45.290 182.200 ;
        RECT 53.170 181.860 54.090 182.200 ;
        RECT 57.130 181.860 58.050 182.200 ;
        RECT 65.610 181.860 66.530 182.200 ;
        RECT 69.570 181.860 70.490 182.200 ;
        RECT 78.370 181.860 79.290 182.200 ;
        RECT 82.330 181.860 83.250 182.200 ;
        RECT 90.810 181.860 91.730 182.200 ;
        RECT 94.770 181.860 95.690 182.200 ;
        RECT 103.570 181.860 104.490 182.200 ;
        RECT 107.530 181.860 108.450 182.200 ;
        RECT 111.570 181.050 111.910 185.380 ;
        RECT 116.010 182.740 116.930 183.080 ;
        RECT 119.970 182.740 120.890 183.080 ;
        RECT 116.010 181.860 116.930 182.200 ;
        RECT 119.970 181.860 120.890 182.200 ;
        RECT 111.570 180.710 114.770 181.050 ;
        RECT 15.210 180.100 16.130 180.440 ;
        RECT 19.170 180.100 20.090 180.440 ;
        RECT 27.970 180.100 28.890 180.440 ;
        RECT 31.930 180.100 32.850 180.440 ;
        RECT 40.410 180.100 41.330 180.440 ;
        RECT 44.370 180.100 45.290 180.440 ;
        RECT 53.170 180.100 54.090 180.440 ;
        RECT 57.130 180.100 58.050 180.440 ;
        RECT 65.610 180.100 66.530 180.440 ;
        RECT 69.570 180.100 70.490 180.440 ;
        RECT 78.370 180.100 79.290 180.440 ;
        RECT 82.330 180.100 83.250 180.440 ;
        RECT 90.810 180.100 91.730 180.440 ;
        RECT 94.770 180.100 95.690 180.440 ;
        RECT 103.570 180.100 104.490 180.440 ;
        RECT 107.530 180.100 108.450 180.440 ;
        RECT 116.010 180.100 116.930 180.440 ;
        RECT 119.970 180.100 120.890 180.440 ;
        RECT 19.170 179.220 20.090 179.560 ;
        RECT 27.970 179.220 28.890 179.560 ;
        RECT 44.370 179.220 45.290 179.560 ;
        RECT 53.170 179.220 54.090 179.560 ;
        RECT 69.570 179.220 70.490 179.560 ;
        RECT 78.370 179.220 79.290 179.560 ;
        RECT 94.770 179.220 95.690 179.560 ;
        RECT 103.570 179.220 104.490 179.560 ;
        RECT 116.010 179.220 116.930 179.560 ;
        RECT 112.860 179.120 113.200 179.165 ;
        RECT 108.750 178.780 114.770 179.120 ;
        RECT 15.210 177.460 16.130 177.800 ;
        RECT 19.170 177.460 20.090 177.800 ;
        RECT 27.970 177.460 28.890 177.800 ;
        RECT 31.930 177.460 32.850 177.800 ;
        RECT 40.410 177.460 41.330 177.800 ;
        RECT 44.370 177.460 45.290 177.800 ;
        RECT 53.170 177.460 54.090 177.800 ;
        RECT 57.130 177.460 58.050 177.800 ;
        RECT 65.610 177.460 66.530 177.800 ;
        RECT 69.570 177.460 70.490 177.800 ;
        RECT 78.370 177.460 79.290 177.800 ;
        RECT 82.330 177.460 83.250 177.800 ;
        RECT 90.810 177.460 91.730 177.800 ;
        RECT 94.770 177.460 95.690 177.800 ;
        RECT 103.570 177.460 104.490 177.800 ;
        RECT 107.530 177.460 108.450 177.800 ;
        RECT 108.750 176.920 109.090 178.780 ;
        RECT 112.860 178.735 113.200 178.780 ;
        RECT 122.130 177.900 123.850 178.240 ;
        RECT 116.010 177.460 116.930 177.800 ;
        RECT 119.970 177.460 120.890 177.800 ;
        RECT 15.210 176.580 16.930 176.920 ;
        RECT 31.770 176.580 33.490 176.920 ;
        RECT 40.410 176.580 42.130 176.920 ;
        RECT 56.970 176.580 58.690 176.920 ;
        RECT 65.610 176.580 67.330 176.920 ;
        RECT 82.170 176.580 83.890 176.920 ;
        RECT 90.810 176.580 92.530 176.920 ;
        RECT 107.370 176.580 109.090 176.920 ;
        RECT 119.970 176.580 120.890 176.920 ;
        RECT 15.210 175.700 16.130 176.040 ;
        RECT 19.170 175.700 20.090 176.040 ;
        RECT 27.970 175.700 28.890 176.040 ;
        RECT 31.930 175.700 32.850 176.040 ;
        RECT 40.410 175.700 41.330 176.040 ;
        RECT 44.370 175.700 45.290 176.040 ;
        RECT 53.170 175.700 54.090 176.040 ;
        RECT 57.130 175.700 58.050 176.040 ;
        RECT 65.610 175.700 66.530 176.040 ;
        RECT 69.570 175.700 70.490 176.040 ;
        RECT 78.370 175.700 79.290 176.040 ;
        RECT 82.330 175.700 83.250 176.040 ;
        RECT 90.810 175.700 91.730 176.040 ;
        RECT 94.770 175.700 95.690 176.040 ;
        RECT 103.570 175.700 104.490 176.040 ;
        RECT 107.530 175.700 108.450 176.040 ;
        RECT 116.010 174.820 116.930 175.160 ;
        RECT 119.970 174.820 120.890 175.160 ;
        RECT 15.210 173.940 16.130 174.280 ;
        RECT 19.170 173.940 20.090 174.280 ;
        RECT 27.970 173.940 28.890 174.280 ;
        RECT 31.930 173.940 32.850 174.280 ;
        RECT 40.410 173.940 41.330 174.280 ;
        RECT 44.370 173.940 45.290 174.280 ;
        RECT 53.170 173.940 54.090 174.280 ;
        RECT 57.130 173.940 58.050 174.280 ;
        RECT 65.610 173.940 66.530 174.280 ;
        RECT 69.570 173.940 70.490 174.280 ;
        RECT 78.370 173.940 79.290 174.280 ;
        RECT 82.330 173.940 83.250 174.280 ;
        RECT 90.810 173.940 91.730 174.280 ;
        RECT 94.770 173.940 95.690 174.280 ;
        RECT 103.570 173.940 104.490 174.280 ;
        RECT 107.530 173.940 108.450 174.280 ;
        RECT 116.010 173.060 116.930 173.400 ;
        RECT 119.970 173.060 120.890 173.400 ;
        RECT 109.530 172.620 110.610 172.960 ;
        RECT 123.510 172.620 123.850 177.900 ;
        RECT 110.310 172.280 123.850 172.620 ;
        RECT 15.210 171.300 16.130 171.640 ;
        RECT 19.170 171.300 20.090 171.640 ;
        RECT 27.970 171.300 28.890 171.640 ;
        RECT 31.930 171.300 32.850 171.640 ;
        RECT 40.410 171.300 41.330 171.640 ;
        RECT 44.370 171.300 45.290 171.640 ;
        RECT 53.170 171.300 54.090 171.640 ;
        RECT 57.130 171.300 58.050 171.640 ;
        RECT 65.610 171.300 66.530 171.640 ;
        RECT 69.570 171.300 70.490 171.640 ;
        RECT 78.370 171.300 79.290 171.640 ;
        RECT 82.330 171.300 83.250 171.640 ;
        RECT 90.810 171.300 91.730 171.640 ;
        RECT 94.770 171.300 95.690 171.640 ;
        RECT 103.570 171.300 104.490 171.640 ;
        RECT 107.530 171.300 108.450 171.640 ;
        RECT 12.710 170.860 13.970 171.200 ;
        RECT 33.590 170.860 34.850 171.200 ;
        RECT 37.910 170.860 39.170 171.200 ;
        RECT 58.790 170.860 60.050 171.200 ;
        RECT 63.110 170.860 64.370 171.200 ;
        RECT 83.990 170.860 85.250 171.200 ;
        RECT 88.310 170.860 89.570 171.200 ;
        RECT 109.190 170.860 110.450 171.200 ;
        RECT 12.710 170.560 13.050 170.860 ;
        RECT 33.590 170.560 33.930 170.860 ;
        RECT 37.910 170.560 38.250 170.860 ;
        RECT 58.790 170.560 59.130 170.860 ;
        RECT 63.110 170.560 63.450 170.860 ;
        RECT 83.990 170.560 84.330 170.860 ;
        RECT 88.310 170.560 88.650 170.860 ;
        RECT 109.190 170.560 109.530 170.860 ;
        RECT 12.710 170.220 127.080 170.560 ;
        RECT 15.210 169.540 16.130 169.880 ;
        RECT 31.930 169.540 32.850 169.880 ;
        RECT 40.410 169.540 41.330 169.880 ;
        RECT 57.130 169.540 58.050 169.880 ;
        RECT 65.610 169.540 66.530 169.880 ;
        RECT 82.330 169.540 83.250 169.880 ;
        RECT 90.810 169.540 91.730 169.880 ;
        RECT 107.530 169.540 108.450 169.880 ;
        RECT 15.210 168.660 16.130 169.000 ;
        RECT 19.170 168.660 20.890 169.000 ;
        RECT 20.550 167.240 20.890 168.660 ;
        RECT 27.170 168.660 28.890 169.000 ;
        RECT 31.930 168.660 32.850 169.000 ;
        RECT 40.410 168.660 41.330 169.000 ;
        RECT 44.370 168.660 46.090 169.000 ;
        RECT 22.050 167.240 22.970 167.820 ;
        RECT 15.210 166.900 16.130 167.240 ;
        RECT 19.170 166.900 22.970 167.240 ;
        RECT 25.090 167.240 26.010 167.820 ;
        RECT 27.170 167.240 27.510 168.660 ;
        RECT 45.750 167.240 46.090 168.660 ;
        RECT 52.370 168.660 54.090 169.000 ;
        RECT 57.130 168.660 58.050 169.000 ;
        RECT 65.610 168.660 66.530 169.000 ;
        RECT 69.570 168.660 71.290 169.000 ;
        RECT 47.250 167.240 48.170 167.820 ;
        RECT 25.090 166.900 28.890 167.240 ;
        RECT 31.930 166.900 32.850 167.240 ;
        RECT 40.410 166.900 41.330 167.240 ;
        RECT 44.370 166.900 48.170 167.240 ;
        RECT 50.290 167.240 51.210 167.820 ;
        RECT 52.370 167.240 52.710 168.660 ;
        RECT 70.950 167.240 71.290 168.660 ;
        RECT 77.570 168.660 79.290 169.000 ;
        RECT 82.330 168.660 83.250 169.000 ;
        RECT 90.810 168.660 91.730 169.000 ;
        RECT 94.770 168.660 96.490 169.000 ;
        RECT 72.450 167.240 73.370 167.820 ;
        RECT 50.290 166.900 54.090 167.240 ;
        RECT 57.130 166.900 58.050 167.240 ;
        RECT 65.610 166.900 66.530 167.240 ;
        RECT 69.570 166.900 73.370 167.240 ;
        RECT 75.490 167.240 76.410 167.820 ;
        RECT 77.570 167.240 77.910 168.660 ;
        RECT 96.150 167.240 96.490 168.660 ;
        RECT 102.770 168.660 104.490 169.000 ;
        RECT 107.530 168.660 108.450 169.000 ;
        RECT 97.650 167.240 98.570 167.820 ;
        RECT 75.490 166.900 79.290 167.240 ;
        RECT 82.330 166.900 83.250 167.240 ;
        RECT 90.810 166.900 91.730 167.240 ;
        RECT 94.770 166.900 98.570 167.240 ;
        RECT 100.690 167.240 101.610 167.820 ;
        RECT 102.770 167.240 103.110 168.660 ;
        RECT 100.690 166.900 104.490 167.240 ;
        RECT 107.530 166.900 108.450 167.240 ;
        RECT 119.970 166.900 120.890 167.240 ;
        RECT 18.160 165.730 18.500 166.650 ;
        RECT 20.550 165.480 20.890 166.900 ;
        RECT 15.210 165.140 16.130 165.480 ;
        RECT 19.170 165.140 20.890 165.480 ;
        RECT 27.170 165.480 27.510 166.900 ;
        RECT 29.560 165.730 29.900 166.650 ;
        RECT 43.360 165.730 43.700 166.650 ;
        RECT 45.750 165.480 46.090 166.900 ;
        RECT 27.170 165.140 28.890 165.480 ;
        RECT 31.930 165.140 32.850 165.480 ;
        RECT 40.410 165.140 41.330 165.480 ;
        RECT 44.370 165.140 46.090 165.480 ;
        RECT 52.370 165.480 52.710 166.900 ;
        RECT 54.760 165.730 55.100 166.650 ;
        RECT 68.560 165.730 68.900 166.650 ;
        RECT 70.950 165.480 71.290 166.900 ;
        RECT 52.370 165.140 54.090 165.480 ;
        RECT 57.130 165.140 58.050 165.480 ;
        RECT 65.610 165.140 66.530 165.480 ;
        RECT 69.570 165.140 71.290 165.480 ;
        RECT 77.570 165.480 77.910 166.900 ;
        RECT 79.960 165.730 80.300 166.650 ;
        RECT 93.760 165.730 94.100 166.650 ;
        RECT 96.150 165.480 96.490 166.900 ;
        RECT 77.570 165.140 79.290 165.480 ;
        RECT 82.330 165.140 83.250 165.480 ;
        RECT 90.810 165.140 91.730 165.480 ;
        RECT 94.770 165.140 96.490 165.480 ;
        RECT 102.770 165.480 103.110 166.900 ;
        RECT 105.160 165.730 105.500 166.650 ;
        RECT 116.010 166.020 116.930 166.360 ;
        RECT 102.770 165.140 104.490 165.480 ;
        RECT 107.530 165.140 108.450 165.480 ;
        RECT 119.970 165.140 120.890 165.480 ;
        RECT 15.210 164.260 16.130 164.600 ;
        RECT 19.170 164.260 20.890 164.600 ;
        RECT 20.550 162.840 20.890 164.260 ;
        RECT 27.170 164.260 28.890 164.600 ;
        RECT 31.930 164.260 32.850 164.600 ;
        RECT 40.410 164.260 41.330 164.600 ;
        RECT 44.370 164.260 46.090 164.600 ;
        RECT 22.050 162.840 22.970 163.420 ;
        RECT 15.210 162.500 16.130 162.840 ;
        RECT 19.170 162.500 22.970 162.840 ;
        RECT 25.090 162.840 26.010 163.420 ;
        RECT 27.170 162.840 27.510 164.260 ;
        RECT 45.750 162.840 46.090 164.260 ;
        RECT 52.370 164.260 54.090 164.600 ;
        RECT 57.130 164.260 58.050 164.600 ;
        RECT 65.610 164.260 66.530 164.600 ;
        RECT 69.570 164.260 71.290 164.600 ;
        RECT 47.250 162.840 48.170 163.420 ;
        RECT 25.090 162.500 28.890 162.840 ;
        RECT 31.930 162.500 32.850 162.840 ;
        RECT 40.410 162.500 41.330 162.840 ;
        RECT 44.370 162.500 48.170 162.840 ;
        RECT 50.290 162.840 51.210 163.420 ;
        RECT 52.370 162.840 52.710 164.260 ;
        RECT 70.950 162.840 71.290 164.260 ;
        RECT 77.570 164.260 79.290 164.600 ;
        RECT 82.330 164.260 83.250 164.600 ;
        RECT 90.810 164.260 91.730 164.600 ;
        RECT 94.770 164.260 96.490 164.600 ;
        RECT 72.450 162.840 73.370 163.420 ;
        RECT 50.290 162.500 54.090 162.840 ;
        RECT 57.130 162.500 58.050 162.840 ;
        RECT 65.610 162.500 66.530 162.840 ;
        RECT 69.570 162.500 73.370 162.840 ;
        RECT 75.490 162.840 76.410 163.420 ;
        RECT 77.570 162.840 77.910 164.260 ;
        RECT 96.150 162.840 96.490 164.260 ;
        RECT 102.770 164.260 104.490 164.600 ;
        RECT 107.530 164.260 108.450 164.600 ;
        RECT 97.650 162.840 98.570 163.420 ;
        RECT 75.490 162.500 79.290 162.840 ;
        RECT 82.330 162.500 83.250 162.840 ;
        RECT 90.810 162.500 91.730 162.840 ;
        RECT 94.770 162.500 98.570 162.840 ;
        RECT 100.690 162.840 101.610 163.420 ;
        RECT 102.770 162.840 103.110 164.260 ;
        RECT 113.850 163.820 115.570 164.160 ;
        RECT 119.970 163.380 120.890 163.720 ;
        RECT 100.690 162.500 104.490 162.840 ;
        RECT 107.530 162.500 108.450 162.840 ;
        RECT 17.375 161.330 17.715 162.250 ;
        RECT 20.550 161.080 20.890 162.500 ;
        RECT 15.210 160.740 16.130 161.080 ;
        RECT 19.170 160.740 20.890 161.080 ;
        RECT 27.170 161.080 27.510 162.500 ;
        RECT 30.345 161.330 30.685 162.250 ;
        RECT 42.575 161.330 42.915 162.250 ;
        RECT 45.750 161.080 46.090 162.500 ;
        RECT 27.170 160.740 28.890 161.080 ;
        RECT 31.930 160.740 32.850 161.080 ;
        RECT 40.410 160.740 41.330 161.080 ;
        RECT 44.370 160.740 46.090 161.080 ;
        RECT 52.370 161.080 52.710 162.500 ;
        RECT 55.545 161.330 55.885 162.250 ;
        RECT 67.775 161.330 68.115 162.250 ;
        RECT 70.950 161.080 71.290 162.500 ;
        RECT 52.370 160.740 54.090 161.080 ;
        RECT 57.130 160.740 58.050 161.080 ;
        RECT 65.610 160.740 66.530 161.080 ;
        RECT 69.570 160.740 71.290 161.080 ;
        RECT 77.570 161.080 77.910 162.500 ;
        RECT 80.745 161.330 81.085 162.250 ;
        RECT 92.975 161.330 93.315 162.250 ;
        RECT 96.150 161.080 96.490 162.500 ;
        RECT 77.570 160.740 79.290 161.080 ;
        RECT 82.330 160.740 83.250 161.080 ;
        RECT 90.810 160.740 91.730 161.080 ;
        RECT 94.770 160.740 96.490 161.080 ;
        RECT 102.770 161.080 103.110 162.500 ;
        RECT 105.945 161.330 106.285 162.250 ;
        RECT 119.970 161.620 120.890 161.960 ;
        RECT 122.130 161.180 123.050 161.520 ;
        RECT 102.770 160.740 104.490 161.080 ;
        RECT 107.530 160.740 108.450 161.080 ;
        RECT 15.210 159.860 16.130 160.200 ;
        RECT 19.170 159.860 20.890 160.200 ;
        RECT 20.550 158.440 20.890 159.860 ;
        RECT 27.170 159.860 28.890 160.200 ;
        RECT 31.930 159.860 32.850 160.200 ;
        RECT 40.410 159.860 41.330 160.200 ;
        RECT 44.370 159.860 46.090 160.200 ;
        RECT 22.050 158.440 22.970 159.020 ;
        RECT 15.210 158.100 16.130 158.440 ;
        RECT 19.170 158.100 22.970 158.440 ;
        RECT 25.090 158.440 26.010 159.020 ;
        RECT 27.170 158.440 27.510 159.860 ;
        RECT 45.750 158.440 46.090 159.860 ;
        RECT 52.370 159.860 54.090 160.200 ;
        RECT 57.130 159.860 58.050 160.200 ;
        RECT 65.610 159.860 66.530 160.200 ;
        RECT 69.570 159.860 71.290 160.200 ;
        RECT 47.250 158.440 48.170 159.020 ;
        RECT 25.090 158.100 28.890 158.440 ;
        RECT 31.930 158.100 32.850 158.440 ;
        RECT 40.410 158.100 41.330 158.440 ;
        RECT 44.370 158.100 48.170 158.440 ;
        RECT 50.290 158.440 51.210 159.020 ;
        RECT 52.370 158.440 52.710 159.860 ;
        RECT 70.950 158.440 71.290 159.860 ;
        RECT 77.570 159.860 79.290 160.200 ;
        RECT 82.330 159.860 83.250 160.200 ;
        RECT 90.810 159.860 91.730 160.200 ;
        RECT 94.770 159.860 96.490 160.200 ;
        RECT 72.450 158.440 73.370 159.020 ;
        RECT 50.290 158.100 54.090 158.440 ;
        RECT 57.130 158.100 58.050 158.440 ;
        RECT 65.610 158.100 66.530 158.440 ;
        RECT 69.570 158.100 73.370 158.440 ;
        RECT 75.490 158.440 76.410 159.020 ;
        RECT 77.570 158.440 77.910 159.860 ;
        RECT 96.150 158.440 96.490 159.860 ;
        RECT 102.770 159.860 104.490 160.200 ;
        RECT 107.530 159.860 108.450 160.200 ;
        RECT 119.970 159.860 120.890 160.200 ;
        RECT 97.650 158.440 98.570 159.020 ;
        RECT 75.490 158.100 79.290 158.440 ;
        RECT 82.330 158.100 83.250 158.440 ;
        RECT 90.810 158.100 91.730 158.440 ;
        RECT 94.770 158.100 98.570 158.440 ;
        RECT 100.690 158.440 101.610 159.020 ;
        RECT 102.770 158.440 103.110 159.860 ;
        RECT 116.010 158.980 116.930 159.320 ;
        RECT 100.690 158.100 104.490 158.440 ;
        RECT 107.530 158.100 108.450 158.440 ;
        RECT 116.010 158.100 116.930 158.440 ;
        RECT 119.970 158.100 120.890 158.440 ;
        RECT 13.210 156.780 14.130 157.120 ;
        RECT 16.660 156.930 17.000 157.850 ;
        RECT 20.550 156.680 20.890 158.100 ;
        RECT 15.210 156.340 16.130 156.680 ;
        RECT 19.170 156.340 20.890 156.680 ;
        RECT 27.170 156.680 27.510 158.100 ;
        RECT 31.060 156.930 31.400 157.850 ;
        RECT 33.930 156.780 34.850 157.120 ;
        RECT 38.410 156.780 39.330 157.120 ;
        RECT 41.860 156.930 42.200 157.850 ;
        RECT 45.750 156.680 46.090 158.100 ;
        RECT 27.170 156.340 28.890 156.680 ;
        RECT 31.930 156.340 32.850 156.680 ;
        RECT 40.410 156.340 41.330 156.680 ;
        RECT 44.370 156.340 46.090 156.680 ;
        RECT 52.370 156.680 52.710 158.100 ;
        RECT 56.260 156.930 56.600 157.850 ;
        RECT 59.130 156.780 60.050 157.120 ;
        RECT 63.610 156.780 64.530 157.120 ;
        RECT 67.060 156.930 67.400 157.850 ;
        RECT 70.950 156.680 71.290 158.100 ;
        RECT 52.370 156.340 54.090 156.680 ;
        RECT 57.130 156.340 58.050 156.680 ;
        RECT 65.610 156.340 66.530 156.680 ;
        RECT 69.570 156.340 71.290 156.680 ;
        RECT 77.570 156.680 77.910 158.100 ;
        RECT 81.460 156.930 81.800 157.850 ;
        RECT 84.330 156.780 85.250 157.120 ;
        RECT 88.810 156.780 89.730 157.120 ;
        RECT 92.260 156.930 92.600 157.850 ;
        RECT 96.150 156.680 96.490 158.100 ;
        RECT 77.570 156.340 79.290 156.680 ;
        RECT 82.330 156.340 83.250 156.680 ;
        RECT 90.810 156.340 91.730 156.680 ;
        RECT 94.770 156.340 96.490 156.680 ;
        RECT 102.770 156.680 103.110 158.100 ;
        RECT 106.660 156.930 107.000 157.850 ;
        RECT 109.530 156.780 110.450 157.120 ;
        RECT 102.770 156.340 104.490 156.680 ;
        RECT 107.530 156.340 108.450 156.680 ;
        RECT 116.010 156.340 116.930 156.680 ;
        RECT 119.970 156.340 120.890 156.680 ;
        RECT 110.910 155.800 120.270 156.140 ;
        RECT 15.210 155.460 16.130 155.800 ;
        RECT 19.170 155.460 20.890 155.800 ;
        RECT 20.550 154.040 20.890 155.460 ;
        RECT 27.170 155.460 28.890 155.800 ;
        RECT 31.930 155.460 32.850 155.800 ;
        RECT 40.410 155.460 41.330 155.800 ;
        RECT 44.370 155.460 46.090 155.800 ;
        RECT 22.050 154.040 22.970 154.620 ;
        RECT 15.210 153.700 16.130 154.040 ;
        RECT 19.170 153.700 22.970 154.040 ;
        RECT 25.090 154.040 26.010 154.620 ;
        RECT 27.170 154.040 27.510 155.460 ;
        RECT 45.750 154.040 46.090 155.460 ;
        RECT 52.370 155.460 54.090 155.800 ;
        RECT 57.130 155.460 58.050 155.800 ;
        RECT 65.610 155.460 66.530 155.800 ;
        RECT 69.570 155.460 71.290 155.800 ;
        RECT 47.250 154.040 48.170 154.620 ;
        RECT 25.090 153.700 28.890 154.040 ;
        RECT 31.930 153.700 32.850 154.040 ;
        RECT 40.410 153.700 41.330 154.040 ;
        RECT 44.370 153.700 48.170 154.040 ;
        RECT 50.290 154.040 51.210 154.620 ;
        RECT 52.370 154.040 52.710 155.460 ;
        RECT 70.950 154.040 71.290 155.460 ;
        RECT 77.570 155.460 79.290 155.800 ;
        RECT 82.330 155.460 83.250 155.800 ;
        RECT 90.810 155.460 91.730 155.800 ;
        RECT 94.770 155.460 96.490 155.800 ;
        RECT 72.450 154.040 73.370 154.620 ;
        RECT 50.290 153.700 54.090 154.040 ;
        RECT 57.130 153.700 58.050 154.040 ;
        RECT 65.610 153.700 66.530 154.040 ;
        RECT 69.570 153.700 73.370 154.040 ;
        RECT 75.490 154.040 76.410 154.620 ;
        RECT 77.570 154.040 77.910 155.460 ;
        RECT 96.150 154.040 96.490 155.460 ;
        RECT 102.770 155.460 104.490 155.800 ;
        RECT 107.530 155.460 108.450 155.800 ;
        RECT 97.650 154.040 98.570 154.620 ;
        RECT 75.490 153.700 79.290 154.040 ;
        RECT 82.330 153.700 83.250 154.040 ;
        RECT 90.810 153.700 91.730 154.040 ;
        RECT 94.770 153.700 98.570 154.040 ;
        RECT 100.690 154.040 101.610 154.620 ;
        RECT 102.770 154.040 103.110 155.460 ;
        RECT 100.690 153.700 104.490 154.040 ;
        RECT 107.530 153.700 108.450 154.040 ;
        RECT 20.550 152.280 20.890 153.700 ;
        RECT 15.210 151.940 16.130 152.280 ;
        RECT 19.170 151.940 20.890 152.280 ;
        RECT 27.170 152.280 27.510 153.700 ;
        RECT 45.750 152.280 46.090 153.700 ;
        RECT 27.170 151.940 28.890 152.280 ;
        RECT 31.930 151.940 32.850 152.280 ;
        RECT 40.410 151.940 41.330 152.280 ;
        RECT 44.370 151.940 46.090 152.280 ;
        RECT 52.370 152.280 52.710 153.700 ;
        RECT 70.950 152.280 71.290 153.700 ;
        RECT 52.370 151.940 54.090 152.280 ;
        RECT 57.130 151.940 58.050 152.280 ;
        RECT 65.610 151.940 66.530 152.280 ;
        RECT 69.570 151.940 71.290 152.280 ;
        RECT 77.570 152.280 77.910 153.700 ;
        RECT 96.150 152.280 96.490 153.700 ;
        RECT 77.570 151.940 79.290 152.280 ;
        RECT 82.330 151.940 83.250 152.280 ;
        RECT 90.810 151.940 91.730 152.280 ;
        RECT 94.770 151.940 96.490 152.280 ;
        RECT 102.770 152.280 103.110 153.700 ;
        RECT 102.770 151.940 104.490 152.280 ;
        RECT 107.530 151.940 108.450 152.280 ;
        RECT 13.050 150.620 102.935 150.960 ;
        RECT 110.910 149.200 111.250 155.800 ;
        RECT 119.970 155.460 120.890 155.800 ;
        RECT 116.010 154.580 116.930 154.920 ;
        RECT 119.970 154.580 120.890 154.920 ;
        RECT 116.010 153.700 116.930 154.040 ;
        RECT 119.970 153.700 120.890 154.040 ;
        RECT 116.010 151.940 116.930 152.280 ;
        RECT 119.970 151.940 120.890 152.280 ;
        RECT 12.710 148.860 13.970 149.200 ;
        RECT 33.590 148.860 34.850 149.200 ;
        RECT 37.910 148.860 39.170 149.200 ;
        RECT 58.790 148.860 60.050 149.200 ;
        RECT 63.110 148.860 64.370 149.200 ;
        RECT 83.990 148.860 85.250 149.200 ;
        RECT 88.310 148.860 89.570 149.200 ;
        RECT 109.190 148.860 111.250 149.200 ;
        RECT 113.270 151.230 117.090 151.570 ;
        RECT 12.710 147.820 13.050 148.860 ;
        RECT 15.210 148.420 16.130 148.760 ;
        RECT 19.170 148.420 20.090 148.760 ;
        RECT 27.970 148.420 28.890 148.760 ;
        RECT 31.930 148.420 32.850 148.760 ;
        RECT 33.590 147.820 33.930 148.860 ;
        RECT 37.910 147.820 38.250 148.860 ;
        RECT 40.410 148.420 41.330 148.760 ;
        RECT 44.370 148.420 45.290 148.760 ;
        RECT 53.170 148.420 54.090 148.760 ;
        RECT 57.130 148.420 58.050 148.760 ;
        RECT 58.790 147.820 59.130 148.860 ;
        RECT 63.110 147.820 63.450 148.860 ;
        RECT 65.610 148.420 66.530 148.760 ;
        RECT 69.570 148.420 70.490 148.760 ;
        RECT 78.370 148.420 79.290 148.760 ;
        RECT 82.330 148.420 83.250 148.760 ;
        RECT 83.990 147.820 84.330 148.860 ;
        RECT 88.310 147.820 88.650 148.860 ;
        RECT 90.810 148.420 91.730 148.760 ;
        RECT 94.770 148.420 95.690 148.760 ;
        RECT 103.570 148.420 104.490 148.760 ;
        RECT 107.530 148.420 108.450 148.760 ;
        RECT 109.190 147.820 109.530 148.860 ;
        RECT 12.710 147.480 110.610 147.820 ;
        RECT 12.870 146.720 110.450 147.060 ;
        RECT 12.870 145.680 13.210 146.720 ;
        RECT 33.590 145.680 33.930 146.720 ;
        RECT 38.070 145.680 38.410 146.720 ;
        RECT 58.790 145.680 59.130 146.720 ;
        RECT 63.270 145.680 63.610 146.720 ;
        RECT 83.990 145.680 84.330 146.720 ;
        RECT 88.470 145.680 88.810 146.720 ;
        RECT 109.190 145.680 109.530 146.720 ;
        RECT 113.270 146.020 113.610 151.230 ;
        RECT 116.010 150.180 116.930 150.520 ;
        RECT 119.970 150.180 120.890 150.520 ;
        RECT 119.970 149.300 120.890 149.640 ;
        RECT 119.970 147.540 120.890 147.880 ;
        RECT 110.150 145.680 113.610 146.020 ;
        RECT 119.970 145.780 120.890 146.120 ;
        RECT 12.870 145.340 14.130 145.680 ;
        RECT 33.590 145.340 34.850 145.680 ;
        RECT 38.070 145.340 39.330 145.680 ;
        RECT 58.790 145.340 60.050 145.680 ;
        RECT 63.270 145.340 64.530 145.680 ;
        RECT 83.990 145.340 85.250 145.680 ;
        RECT 88.470 145.340 89.730 145.680 ;
        RECT 109.190 145.340 110.450 145.680 ;
        RECT 122.130 145.340 123.050 145.680 ;
        RECT 15.210 144.900 16.130 145.240 ;
        RECT 19.170 144.900 20.090 145.240 ;
        RECT 27.970 144.900 28.890 145.240 ;
        RECT 31.930 144.900 32.850 145.240 ;
        RECT 40.410 144.900 41.330 145.240 ;
        RECT 44.370 144.900 45.290 145.240 ;
        RECT 53.170 144.900 54.090 145.240 ;
        RECT 57.130 144.900 58.050 145.240 ;
        RECT 65.610 144.900 66.530 145.240 ;
        RECT 69.570 144.900 70.490 145.240 ;
        RECT 78.370 144.900 79.290 145.240 ;
        RECT 82.330 144.900 83.250 145.240 ;
        RECT 90.810 144.900 91.730 145.240 ;
        RECT 94.770 144.900 95.690 145.240 ;
        RECT 103.570 144.900 104.490 145.240 ;
        RECT 107.530 144.900 108.450 145.240 ;
        RECT 119.970 144.020 120.890 144.360 ;
        RECT 15.210 143.140 16.130 143.480 ;
        RECT 19.170 143.140 20.090 143.480 ;
        RECT 27.970 143.140 28.890 143.480 ;
        RECT 31.930 143.140 32.850 143.480 ;
        RECT 40.410 143.140 41.330 143.480 ;
        RECT 44.370 143.140 45.290 143.480 ;
        RECT 53.170 143.140 54.090 143.480 ;
        RECT 57.130 143.140 58.050 143.480 ;
        RECT 65.610 143.140 66.530 143.480 ;
        RECT 69.570 143.140 70.490 143.480 ;
        RECT 78.370 143.140 79.290 143.480 ;
        RECT 82.330 143.140 83.250 143.480 ;
        RECT 90.810 143.140 91.730 143.480 ;
        RECT 94.770 143.140 95.690 143.480 ;
        RECT 103.570 143.140 104.490 143.480 ;
        RECT 107.530 143.140 108.450 143.480 ;
        RECT 116.010 143.140 116.930 143.480 ;
        RECT 19.170 142.260 20.090 142.600 ;
        RECT 27.970 142.260 28.890 142.600 ;
        RECT 44.370 142.260 45.290 142.600 ;
        RECT 53.170 142.260 54.090 142.600 ;
        RECT 69.570 142.260 70.490 142.600 ;
        RECT 78.370 142.260 79.290 142.600 ;
        RECT 94.770 142.260 95.690 142.600 ;
        RECT 103.570 142.260 104.490 142.600 ;
        RECT 15.210 141.380 16.130 141.720 ;
        RECT 31.930 141.380 32.850 141.720 ;
        RECT 40.410 141.380 41.330 141.720 ;
        RECT 57.130 141.380 58.050 141.720 ;
        RECT 65.610 141.380 66.530 141.720 ;
        RECT 82.330 141.380 83.250 141.720 ;
        RECT 90.810 141.380 91.730 141.720 ;
        RECT 107.530 141.380 108.450 141.720 ;
        RECT 113.850 140.940 114.770 141.280 ;
        RECT 15.210 140.500 16.130 140.840 ;
        RECT 31.930 140.500 32.850 140.840 ;
        RECT 40.410 140.500 41.330 140.840 ;
        RECT 57.130 140.500 58.050 140.840 ;
        RECT 65.610 140.500 66.530 140.840 ;
        RECT 82.330 140.500 83.250 140.840 ;
        RECT 90.810 140.500 91.730 140.840 ;
        RECT 107.530 140.500 108.450 140.840 ;
        RECT 29.330 138.500 38.410 138.840 ;
        RECT 29.330 138.200 29.670 138.500 ;
        RECT 15.210 137.860 16.130 138.200 ;
        RECT 19.330 137.860 21.190 138.200 ;
        RECT 27.810 137.860 29.670 138.200 ;
        RECT 31.930 137.860 32.850 138.200 ;
        RECT 19.170 136.980 20.090 137.320 ;
        RECT 13.210 136.540 14.130 136.880 ;
        RECT 20.850 136.240 21.190 137.860 ;
        RECT 27.970 136.980 28.890 137.320 ;
        RECT 38.070 136.880 38.410 138.500 ;
        RECT 54.530 138.500 63.610 138.840 ;
        RECT 54.530 138.200 54.870 138.500 ;
        RECT 40.410 137.860 41.330 138.200 ;
        RECT 44.530 137.860 46.390 138.200 ;
        RECT 53.010 137.860 54.870 138.200 ;
        RECT 57.130 137.860 58.050 138.200 ;
        RECT 44.370 136.980 45.290 137.320 ;
        RECT 33.590 136.540 34.850 136.880 ;
        RECT 38.070 136.540 39.330 136.880 ;
        RECT 33.590 136.240 33.930 136.540 ;
        RECT 20.850 135.900 33.930 136.240 ;
        RECT 46.050 136.240 46.390 137.860 ;
        RECT 53.170 136.980 54.090 137.320 ;
        RECT 63.270 136.880 63.610 138.500 ;
        RECT 79.730 138.500 88.810 138.840 ;
        RECT 79.730 138.200 80.070 138.500 ;
        RECT 65.610 137.860 66.530 138.200 ;
        RECT 69.730 137.860 71.590 138.200 ;
        RECT 78.210 137.860 80.070 138.200 ;
        RECT 82.330 137.860 83.250 138.200 ;
        RECT 69.570 136.980 70.490 137.320 ;
        RECT 58.790 136.540 60.050 136.880 ;
        RECT 63.270 136.540 64.530 136.880 ;
        RECT 58.790 136.240 59.130 136.540 ;
        RECT 46.050 135.900 59.130 136.240 ;
        RECT 71.250 136.240 71.590 137.860 ;
        RECT 78.370 136.980 79.290 137.320 ;
        RECT 88.470 136.880 88.810 138.500 ;
        RECT 104.930 138.200 105.270 138.500 ;
        RECT 90.810 137.860 91.730 138.200 ;
        RECT 94.930 137.860 96.790 138.200 ;
        RECT 103.410 137.860 105.270 138.200 ;
        RECT 107.530 137.860 108.450 138.200 ;
        RECT 94.770 136.980 95.690 137.320 ;
        RECT 83.990 136.540 85.250 136.880 ;
        RECT 88.470 136.540 89.730 136.880 ;
        RECT 83.990 136.240 84.330 136.540 ;
        RECT 71.250 135.900 84.330 136.240 ;
        RECT 96.450 136.240 96.790 137.860 ;
        RECT 103.570 136.980 104.490 137.320 ;
        RECT 119.970 136.980 120.890 137.320 ;
        RECT 109.190 136.540 110.450 136.880 ;
        RECT 109.190 136.240 109.530 136.540 ;
        RECT 96.450 135.900 109.530 136.240 ;
        RECT 116.010 136.100 116.930 136.440 ;
        RECT 15.210 135.220 16.130 135.560 ;
        RECT 19.170 135.220 20.090 135.560 ;
        RECT 27.970 135.220 28.890 135.560 ;
        RECT 31.930 135.220 32.850 135.560 ;
        RECT 40.410 135.220 41.330 135.560 ;
        RECT 44.370 135.220 45.290 135.560 ;
        RECT 53.170 135.220 54.090 135.560 ;
        RECT 57.130 135.220 58.050 135.560 ;
        RECT 65.610 135.220 66.530 135.560 ;
        RECT 69.570 135.220 70.490 135.560 ;
        RECT 78.370 135.220 79.290 135.560 ;
        RECT 82.330 135.220 83.250 135.560 ;
        RECT 90.810 135.220 91.730 135.560 ;
        RECT 94.770 135.220 95.690 135.560 ;
        RECT 103.570 135.220 104.490 135.560 ;
        RECT 107.530 135.220 108.450 135.560 ;
        RECT 116.010 135.220 116.930 135.560 ;
        RECT 119.970 135.220 120.890 135.560 ;
        RECT 15.210 134.340 16.130 134.680 ;
        RECT 19.170 134.340 20.090 134.680 ;
        RECT 27.970 134.340 28.890 134.680 ;
        RECT 31.930 134.340 32.850 134.680 ;
        RECT 40.410 134.340 41.330 134.680 ;
        RECT 44.370 134.340 45.290 134.680 ;
        RECT 53.170 134.340 54.090 134.680 ;
        RECT 57.130 134.340 58.050 134.680 ;
        RECT 65.610 134.340 66.530 134.680 ;
        RECT 69.570 134.340 70.490 134.680 ;
        RECT 78.370 134.340 79.290 134.680 ;
        RECT 82.330 134.340 83.250 134.680 ;
        RECT 90.810 134.340 91.730 134.680 ;
        RECT 94.770 134.340 95.690 134.680 ;
        RECT 103.570 134.340 104.490 134.680 ;
        RECT 107.530 134.340 108.450 134.680 ;
        RECT 116.010 134.340 116.930 134.680 ;
        RECT 119.970 134.340 120.890 134.680 ;
        RECT 69.560 130.690 69.900 130.980 ;
        RECT 93.760 130.690 94.100 130.980 ;
        RECT 69.560 130.350 94.100 130.690 ;
        RECT 69.560 130.060 69.900 130.350 ;
        RECT 93.760 130.060 94.100 130.350 ;
        RECT 70.500 129.760 70.840 130.050 ;
        RECT 79.960 129.760 80.300 130.050 ;
        RECT 70.500 129.420 80.300 129.760 ;
        RECT 70.500 129.130 70.840 129.420 ;
        RECT 79.960 129.130 80.300 129.420 ;
        RECT 68.560 128.830 68.900 129.120 ;
        RECT 71.440 128.830 71.780 129.120 ;
        RECT 68.560 128.490 71.780 128.830 ;
        RECT 68.560 128.200 68.900 128.490 ;
        RECT 71.440 128.200 71.780 128.490 ;
        RECT 54.760 127.900 55.100 128.190 ;
        RECT 72.380 127.900 72.720 128.190 ;
        RECT 54.760 127.560 72.720 127.900 ;
        RECT 54.760 127.270 55.100 127.560 ;
        RECT 72.380 127.270 72.720 127.560 ;
        RECT 43.360 126.970 43.700 127.260 ;
        RECT 73.320 126.970 73.660 127.260 ;
        RECT 43.360 126.630 73.660 126.970 ;
        RECT 43.360 126.340 43.700 126.630 ;
        RECT 73.320 126.340 73.660 126.630 ;
        RECT 29.560 126.040 29.900 126.330 ;
        RECT 75.200 126.040 75.540 126.330 ;
        RECT 29.560 125.700 75.540 126.040 ;
        RECT 29.560 125.410 29.900 125.700 ;
        RECT 75.200 125.410 75.540 125.700 ;
        RECT 18.160 125.110 18.500 125.400 ;
        RECT 77.080 125.110 77.420 125.400 ;
        RECT 18.160 124.770 77.420 125.110 ;
        RECT 18.160 124.480 18.500 124.770 ;
        RECT 77.080 124.480 77.420 124.770 ;
        RECT 42.575 124.180 42.915 124.470 ;
        RECT 62.600 124.180 62.940 124.470 ;
        RECT 42.575 123.840 62.940 124.180 ;
        RECT 42.575 123.550 42.915 123.840 ;
        RECT 62.600 123.550 62.940 123.840 ;
        RECT 30.340 123.250 30.680 123.540 ;
        RECT 60.720 123.250 61.060 123.540 ;
        RECT 30.340 122.910 61.060 123.250 ;
        RECT 30.340 122.620 30.680 122.910 ;
        RECT 60.720 122.620 61.060 122.910 ;
        RECT 17.375 122.320 17.715 122.610 ;
        RECT 58.840 122.320 59.180 122.610 ;
        RECT 17.375 121.980 59.180 122.320 ;
        RECT 17.375 121.690 17.715 121.980 ;
        RECT 58.840 121.690 59.180 121.980 ;
        RECT 66.360 121.390 66.700 121.680 ;
        RECT 92.260 121.390 92.600 121.680 ;
        RECT 66.360 121.050 92.600 121.390 ;
        RECT 66.360 120.760 66.700 121.050 ;
        RECT 92.260 120.760 92.600 121.050 ;
        RECT 65.420 120.460 65.760 120.750 ;
        RECT 81.455 120.460 81.795 120.750 ;
        RECT 65.420 120.120 81.795 120.460 ;
        RECT 65.420 119.830 65.760 120.120 ;
        RECT 81.455 119.830 81.795 120.120 ;
        RECT 64.480 119.530 64.820 119.820 ;
        RECT 67.060 119.530 67.400 119.820 ;
        RECT 64.480 119.190 67.400 119.530 ;
        RECT 64.480 118.900 64.820 119.190 ;
        RECT 67.060 118.900 67.400 119.190 ;
        RECT 56.255 118.600 56.595 118.890 ;
        RECT 63.540 118.600 63.880 118.890 ;
        RECT 56.255 118.260 63.880 118.600 ;
        RECT 56.255 117.970 56.595 118.260 ;
        RECT 63.540 117.970 63.880 118.260 ;
        RECT 41.860 117.670 42.200 117.960 ;
        RECT 61.660 117.670 62.000 117.960 ;
        RECT 41.860 117.330 62.000 117.670 ;
        RECT 41.860 117.040 42.200 117.330 ;
        RECT 61.660 117.040 62.000 117.330 ;
        RECT 31.055 116.740 31.395 117.030 ;
        RECT 59.780 116.740 60.120 117.030 ;
        RECT 31.055 116.400 60.120 116.740 ;
        RECT 31.055 116.110 31.395 116.400 ;
        RECT 59.780 116.110 60.120 116.400 ;
        RECT 16.660 115.810 17.000 116.100 ;
        RECT 57.900 115.810 58.240 116.100 ;
        RECT 16.660 115.470 58.240 115.810 ;
        RECT 16.660 115.180 17.000 115.470 ;
        RECT 57.900 115.180 58.240 115.470 ;
        RECT 38.410 114.880 38.750 115.170 ;
        RECT 74.260 114.880 74.600 115.170 ;
        RECT 38.410 114.540 74.600 114.880 ;
        RECT 38.410 114.250 38.750 114.540 ;
        RECT 74.260 114.250 74.600 114.540 ;
        RECT 33.930 113.950 34.270 114.240 ;
        RECT 76.140 113.950 76.480 114.240 ;
        RECT 33.930 113.610 76.480 113.950 ;
        RECT 33.930 113.320 34.270 113.610 ;
        RECT 76.140 113.320 76.480 113.610 ;
        RECT 13.210 113.020 13.550 113.310 ;
        RECT 78.020 113.020 78.360 113.310 ;
        RECT 13.210 112.680 78.360 113.020 ;
        RECT 13.210 112.390 13.550 112.680 ;
        RECT 78.020 112.390 78.360 112.680 ;
        RECT 113.850 111.160 114.190 113.440 ;
        RECT 55.140 110.820 56.060 111.160 ;
        RECT 113.850 110.820 114.770 111.160 ;
        RECT 55.140 106.510 55.480 110.820 ;
        RECT 115.230 109.300 115.570 113.440 ;
        RECT 80.780 108.960 81.700 109.300 ;
        RECT 115.230 108.960 116.150 109.300 ;
        RECT 80.780 106.510 81.120 108.960 ;
        RECT 12.240 38.170 12.580 106.510 ;
        RECT 22.800 104.930 23.140 105.850 ;
        RECT 57.900 105.560 58.240 105.850 ;
        RECT 56.120 105.220 58.240 105.560 ;
        RECT 57.900 104.930 58.240 105.220 ;
        RECT 78.020 105.560 78.360 105.850 ;
        RECT 78.020 105.220 80.140 105.560 ;
        RECT 78.020 104.930 78.360 105.220 ;
        RECT 113.120 104.930 113.460 105.850 ;
        RECT 21.480 101.910 21.820 102.830 ;
        RECT 25.440 101.910 25.780 102.830 ;
        RECT 42.600 101.910 42.940 102.830 ;
        RECT 46.560 101.910 46.900 102.830 ;
        RECT 57.900 102.540 58.240 102.830 ;
        RECT 56.120 102.200 58.240 102.540 ;
        RECT 57.900 101.910 58.240 102.200 ;
        RECT 78.020 102.540 78.360 102.830 ;
        RECT 78.020 102.200 80.140 102.540 ;
        RECT 78.020 101.910 78.360 102.200 ;
        RECT 89.360 101.910 89.700 102.830 ;
        RECT 93.320 101.910 93.660 102.830 ;
        RECT 110.480 101.910 110.820 102.830 ;
        RECT 114.440 101.910 114.780 102.830 ;
        RECT 18.840 98.890 19.180 99.810 ;
        RECT 20.160 98.890 20.500 99.810 ;
        RECT 26.760 98.890 27.100 99.810 ;
        RECT 28.080 98.890 28.420 99.810 ;
        RECT 39.960 98.890 40.300 99.810 ;
        RECT 41.280 98.890 41.620 99.810 ;
        RECT 47.880 98.890 48.220 99.810 ;
        RECT 49.200 98.890 49.540 99.810 ;
        RECT 57.900 99.520 58.240 99.810 ;
        RECT 56.120 99.180 58.240 99.520 ;
        RECT 57.900 98.890 58.240 99.180 ;
        RECT 78.020 99.520 78.360 99.810 ;
        RECT 78.020 99.180 80.140 99.520 ;
        RECT 78.020 98.890 78.360 99.180 ;
        RECT 86.720 98.890 87.060 99.810 ;
        RECT 88.040 98.890 88.380 99.810 ;
        RECT 94.640 98.890 94.980 99.810 ;
        RECT 95.960 98.890 96.300 99.810 ;
        RECT 107.840 98.890 108.180 99.810 ;
        RECT 109.160 98.890 109.500 99.810 ;
        RECT 115.760 98.890 116.100 99.810 ;
        RECT 117.080 98.890 117.420 99.810 ;
        RECT 24.120 95.870 24.460 96.790 ;
        RECT 43.920 95.870 44.260 96.790 ;
        RECT 57.900 96.500 58.240 96.790 ;
        RECT 56.120 96.160 58.240 96.500 ;
        RECT 57.900 95.870 58.240 96.160 ;
        RECT 78.020 96.500 78.360 96.790 ;
        RECT 78.020 96.160 80.140 96.500 ;
        RECT 78.020 95.870 78.360 96.160 ;
        RECT 92.000 95.870 92.340 96.790 ;
        RECT 111.800 95.870 112.140 96.790 ;
        RECT 13.560 92.850 13.900 93.770 ;
        RECT 14.880 92.850 15.220 93.770 ;
        RECT 16.200 92.850 16.540 93.770 ;
        RECT 17.520 92.850 17.860 93.770 ;
        RECT 29.400 92.850 29.740 93.770 ;
        RECT 30.720 92.850 31.060 93.770 ;
        RECT 32.040 92.850 32.380 93.770 ;
        RECT 33.360 92.850 33.700 93.770 ;
        RECT 34.680 92.850 35.020 93.770 ;
        RECT 36.000 92.850 36.340 93.770 ;
        RECT 37.320 92.850 37.660 93.770 ;
        RECT 38.640 92.850 38.980 93.770 ;
        RECT 50.520 92.850 50.860 93.770 ;
        RECT 51.840 92.850 52.180 93.770 ;
        RECT 53.160 92.850 53.500 93.770 ;
        RECT 54.480 92.850 54.820 93.770 ;
        RECT 57.900 93.480 58.240 93.770 ;
        RECT 56.120 93.140 58.240 93.480 ;
        RECT 57.900 92.850 58.240 93.140 ;
        RECT 78.020 93.480 78.360 93.770 ;
        RECT 78.020 93.140 80.140 93.480 ;
        RECT 78.020 92.850 78.360 93.140 ;
        RECT 81.440 92.850 81.780 93.770 ;
        RECT 82.760 92.850 83.100 93.770 ;
        RECT 84.080 92.850 84.420 93.770 ;
        RECT 85.400 92.850 85.740 93.770 ;
        RECT 97.280 92.850 97.620 93.770 ;
        RECT 98.600 92.850 98.940 93.770 ;
        RECT 99.920 92.850 100.260 93.770 ;
        RECT 101.240 92.850 101.580 93.770 ;
        RECT 102.560 92.850 102.900 93.770 ;
        RECT 103.880 92.850 104.220 93.770 ;
        RECT 105.200 92.850 105.540 93.770 ;
        RECT 106.520 92.850 106.860 93.770 ;
        RECT 118.400 92.850 118.740 93.770 ;
        RECT 119.720 92.850 120.060 93.770 ;
        RECT 121.040 92.850 121.380 93.770 ;
        RECT 122.360 92.850 122.700 93.770 ;
        RECT 45.240 89.830 45.580 90.750 ;
        RECT 57.900 90.460 58.240 90.750 ;
        RECT 56.120 90.120 58.240 90.460 ;
        RECT 57.900 89.830 58.240 90.120 ;
        RECT 78.020 90.460 78.360 90.750 ;
        RECT 78.020 90.120 80.140 90.460 ;
        RECT 78.020 89.830 78.360 90.120 ;
        RECT 90.680 89.830 91.020 90.750 ;
        RECT 22.800 87.930 23.140 88.850 ;
        RECT 61.660 88.560 62.000 88.850 ;
        RECT 56.120 88.220 62.000 88.560 ;
        RECT 61.660 87.930 62.000 88.220 ;
        RECT 74.260 88.560 74.600 88.850 ;
        RECT 74.260 88.220 80.140 88.560 ;
        RECT 74.260 87.930 74.600 88.220 ;
        RECT 113.120 87.930 113.460 88.850 ;
        RECT 21.480 84.910 21.820 85.830 ;
        RECT 25.440 84.910 25.780 85.830 ;
        RECT 42.600 84.910 42.940 85.830 ;
        RECT 46.560 84.910 46.900 85.830 ;
        RECT 61.660 85.540 62.000 85.830 ;
        RECT 56.120 85.200 62.000 85.540 ;
        RECT 61.660 84.910 62.000 85.200 ;
        RECT 74.260 85.540 74.600 85.830 ;
        RECT 74.260 85.200 80.140 85.540 ;
        RECT 74.260 84.910 74.600 85.200 ;
        RECT 89.360 84.910 89.700 85.830 ;
        RECT 93.320 84.910 93.660 85.830 ;
        RECT 110.480 84.910 110.820 85.830 ;
        RECT 114.440 84.910 114.780 85.830 ;
        RECT 18.840 81.890 19.180 82.810 ;
        RECT 20.160 81.890 20.500 82.810 ;
        RECT 26.760 81.890 27.100 82.810 ;
        RECT 28.080 81.890 28.420 82.810 ;
        RECT 39.960 81.890 40.300 82.810 ;
        RECT 41.280 81.890 41.620 82.810 ;
        RECT 47.880 81.890 48.220 82.810 ;
        RECT 49.200 81.890 49.540 82.810 ;
        RECT 62.600 82.520 62.940 82.810 ;
        RECT 56.120 82.180 62.940 82.520 ;
        RECT 62.600 81.890 62.940 82.180 ;
        RECT 73.320 82.520 73.660 82.810 ;
        RECT 73.320 82.180 80.140 82.520 ;
        RECT 73.320 81.890 73.660 82.180 ;
        RECT 86.720 81.890 87.060 82.810 ;
        RECT 88.040 81.890 88.380 82.810 ;
        RECT 94.640 81.890 94.980 82.810 ;
        RECT 95.960 81.890 96.300 82.810 ;
        RECT 107.840 81.890 108.180 82.810 ;
        RECT 109.160 81.890 109.500 82.810 ;
        RECT 115.760 81.890 116.100 82.810 ;
        RECT 117.080 81.890 117.420 82.810 ;
        RECT 24.120 78.870 24.460 79.790 ;
        RECT 43.920 78.870 44.260 79.790 ;
        RECT 61.660 79.500 62.000 79.790 ;
        RECT 56.120 79.160 62.000 79.500 ;
        RECT 61.660 78.870 62.000 79.160 ;
        RECT 74.260 79.500 74.600 79.790 ;
        RECT 74.260 79.160 80.140 79.500 ;
        RECT 74.260 78.870 74.600 79.160 ;
        RECT 92.000 78.870 92.340 79.790 ;
        RECT 111.800 78.870 112.140 79.790 ;
        RECT 13.560 75.850 13.900 76.770 ;
        RECT 14.880 75.850 15.220 76.770 ;
        RECT 16.200 75.850 16.540 76.770 ;
        RECT 17.520 75.850 17.860 76.770 ;
        RECT 29.400 75.850 29.740 76.770 ;
        RECT 30.720 75.850 31.060 76.770 ;
        RECT 32.040 75.850 32.380 76.770 ;
        RECT 33.360 75.850 33.700 76.770 ;
        RECT 34.680 75.850 35.020 76.770 ;
        RECT 36.000 75.850 36.340 76.770 ;
        RECT 37.320 75.850 37.660 76.770 ;
        RECT 38.640 75.850 38.980 76.770 ;
        RECT 50.520 75.850 50.860 76.770 ;
        RECT 51.840 75.850 52.180 76.770 ;
        RECT 53.160 75.850 53.500 76.770 ;
        RECT 54.480 75.850 54.820 76.770 ;
        RECT 60.720 76.480 61.060 76.770 ;
        RECT 56.120 76.140 61.060 76.480 ;
        RECT 60.720 75.850 61.060 76.140 ;
        RECT 75.200 76.480 75.540 76.770 ;
        RECT 75.200 76.140 80.140 76.480 ;
        RECT 75.200 75.850 75.540 76.140 ;
        RECT 81.440 75.850 81.780 76.770 ;
        RECT 82.760 75.850 83.100 76.770 ;
        RECT 84.080 75.850 84.420 76.770 ;
        RECT 85.400 75.850 85.740 76.770 ;
        RECT 97.280 75.850 97.620 76.770 ;
        RECT 98.600 75.850 98.940 76.770 ;
        RECT 99.920 75.850 100.260 76.770 ;
        RECT 101.240 75.850 101.580 76.770 ;
        RECT 102.560 75.850 102.900 76.770 ;
        RECT 103.880 75.850 104.220 76.770 ;
        RECT 105.200 75.850 105.540 76.770 ;
        RECT 106.520 75.850 106.860 76.770 ;
        RECT 118.400 75.850 118.740 76.770 ;
        RECT 119.720 75.850 120.060 76.770 ;
        RECT 121.040 75.850 121.380 76.770 ;
        RECT 122.360 75.850 122.700 76.770 ;
        RECT 45.240 72.830 45.580 73.750 ;
        RECT 61.660 73.460 62.000 73.750 ;
        RECT 56.120 73.120 62.000 73.460 ;
        RECT 61.660 72.830 62.000 73.120 ;
        RECT 74.260 73.460 74.600 73.750 ;
        RECT 74.260 73.120 80.140 73.460 ;
        RECT 74.260 72.830 74.600 73.120 ;
        RECT 90.680 72.830 91.020 73.750 ;
        RECT 22.800 70.930 23.140 71.850 ;
        RECT 66.360 71.560 66.700 71.850 ;
        RECT 56.120 71.220 66.700 71.560 ;
        RECT 66.360 70.930 66.700 71.220 ;
        RECT 69.560 71.560 69.900 71.850 ;
        RECT 69.560 71.220 80.140 71.560 ;
        RECT 69.560 70.930 69.900 71.220 ;
        RECT 113.120 70.930 113.460 71.850 ;
        RECT 21.480 67.910 21.820 68.830 ;
        RECT 25.440 67.910 25.780 68.830 ;
        RECT 42.600 67.910 42.940 68.830 ;
        RECT 46.560 67.910 46.900 68.830 ;
        RECT 64.480 68.540 64.820 68.830 ;
        RECT 56.120 68.200 64.820 68.540 ;
        RECT 64.480 67.910 64.820 68.200 ;
        RECT 71.440 68.540 71.780 68.830 ;
        RECT 71.440 68.200 80.140 68.540 ;
        RECT 71.440 67.910 71.780 68.200 ;
        RECT 89.360 67.910 89.700 68.830 ;
        RECT 93.320 67.910 93.660 68.830 ;
        RECT 110.480 67.910 110.820 68.830 ;
        RECT 114.440 67.910 114.780 68.830 ;
        RECT 18.840 64.890 19.180 65.810 ;
        RECT 20.160 64.890 20.500 65.810 ;
        RECT 26.760 64.890 27.100 65.810 ;
        RECT 28.080 64.890 28.420 65.810 ;
        RECT 39.960 64.890 40.300 65.810 ;
        RECT 41.280 64.890 41.620 65.810 ;
        RECT 47.880 64.890 48.220 65.810 ;
        RECT 49.200 64.890 49.540 65.810 ;
        RECT 63.540 65.520 63.880 65.810 ;
        RECT 56.120 65.180 63.880 65.520 ;
        RECT 63.540 64.890 63.880 65.180 ;
        RECT 72.380 65.520 72.720 65.810 ;
        RECT 72.380 65.180 80.140 65.520 ;
        RECT 72.380 64.890 72.720 65.180 ;
        RECT 86.720 64.890 87.060 65.810 ;
        RECT 88.040 64.890 88.380 65.810 ;
        RECT 94.640 64.890 94.980 65.810 ;
        RECT 95.960 64.890 96.300 65.810 ;
        RECT 107.840 64.890 108.180 65.810 ;
        RECT 109.160 64.890 109.500 65.810 ;
        RECT 115.760 64.890 116.100 65.810 ;
        RECT 117.080 64.890 117.420 65.810 ;
        RECT 24.120 61.870 24.460 62.790 ;
        RECT 43.920 61.870 44.260 62.790 ;
        RECT 65.420 62.500 65.760 62.790 ;
        RECT 56.120 62.160 65.760 62.500 ;
        RECT 65.420 61.870 65.760 62.160 ;
        RECT 70.500 62.500 70.840 62.790 ;
        RECT 70.500 62.160 80.140 62.500 ;
        RECT 70.500 61.870 70.840 62.160 ;
        RECT 92.000 61.870 92.340 62.790 ;
        RECT 111.800 61.870 112.140 62.790 ;
        RECT 13.560 58.850 13.900 59.770 ;
        RECT 14.880 58.850 15.220 59.770 ;
        RECT 16.200 58.850 16.540 59.770 ;
        RECT 17.520 58.850 17.860 59.770 ;
        RECT 29.400 58.850 29.740 59.770 ;
        RECT 30.720 58.850 31.060 59.770 ;
        RECT 32.040 58.850 32.380 59.770 ;
        RECT 33.360 58.850 33.700 59.770 ;
        RECT 34.680 58.850 35.020 59.770 ;
        RECT 36.000 58.850 36.340 59.770 ;
        RECT 37.320 58.850 37.660 59.770 ;
        RECT 38.640 58.850 38.980 59.770 ;
        RECT 50.520 58.850 50.860 59.770 ;
        RECT 51.840 58.850 52.180 59.770 ;
        RECT 53.160 58.850 53.500 59.770 ;
        RECT 54.480 58.850 54.820 59.770 ;
        RECT 59.780 59.480 60.120 59.770 ;
        RECT 56.120 59.140 60.120 59.480 ;
        RECT 59.780 58.850 60.120 59.140 ;
        RECT 76.140 59.480 76.480 59.770 ;
        RECT 76.140 59.140 80.140 59.480 ;
        RECT 76.140 58.850 76.480 59.140 ;
        RECT 81.440 58.850 81.780 59.770 ;
        RECT 82.760 58.850 83.100 59.770 ;
        RECT 84.080 58.850 84.420 59.770 ;
        RECT 85.400 58.850 85.740 59.770 ;
        RECT 97.280 58.850 97.620 59.770 ;
        RECT 98.600 58.850 98.940 59.770 ;
        RECT 99.920 58.850 100.260 59.770 ;
        RECT 101.240 58.850 101.580 59.770 ;
        RECT 102.560 58.850 102.900 59.770 ;
        RECT 103.880 58.850 104.220 59.770 ;
        RECT 105.200 58.850 105.540 59.770 ;
        RECT 106.520 58.850 106.860 59.770 ;
        RECT 118.400 58.850 118.740 59.770 ;
        RECT 119.720 58.850 120.060 59.770 ;
        RECT 121.040 58.850 121.380 59.770 ;
        RECT 122.360 58.850 122.700 59.770 ;
        RECT 45.240 55.830 45.580 56.750 ;
        RECT 90.680 55.830 91.020 56.750 ;
        RECT 22.800 53.930 23.140 54.850 ;
        RECT 58.840 54.560 59.180 54.850 ;
        RECT 56.120 54.220 59.180 54.560 ;
        RECT 58.840 53.930 59.180 54.220 ;
        RECT 77.080 54.560 77.420 54.850 ;
        RECT 77.080 54.220 80.140 54.560 ;
        RECT 77.080 53.930 77.420 54.220 ;
        RECT 113.120 53.930 113.460 54.850 ;
        RECT 21.480 50.910 21.820 51.830 ;
        RECT 25.440 50.910 25.780 51.830 ;
        RECT 42.600 50.910 42.940 51.830 ;
        RECT 46.560 50.910 46.900 51.830 ;
        RECT 58.840 51.540 59.180 51.830 ;
        RECT 56.120 51.200 59.180 51.540 ;
        RECT 58.840 50.910 59.180 51.200 ;
        RECT 77.080 51.540 77.420 51.830 ;
        RECT 77.080 51.200 80.140 51.540 ;
        RECT 77.080 50.910 77.420 51.200 ;
        RECT 89.360 50.910 89.700 51.830 ;
        RECT 93.320 50.910 93.660 51.830 ;
        RECT 110.480 50.910 110.820 51.830 ;
        RECT 114.440 50.910 114.780 51.830 ;
        RECT 18.840 47.890 19.180 48.810 ;
        RECT 20.160 47.890 20.500 48.810 ;
        RECT 26.760 47.890 27.100 48.810 ;
        RECT 28.080 47.890 28.420 48.810 ;
        RECT 39.960 47.890 40.300 48.810 ;
        RECT 41.280 47.890 41.620 48.810 ;
        RECT 47.880 47.890 48.220 48.810 ;
        RECT 49.200 47.890 49.540 48.810 ;
        RECT 58.840 48.520 59.180 48.810 ;
        RECT 56.120 48.180 59.180 48.520 ;
        RECT 58.840 47.890 59.180 48.180 ;
        RECT 77.080 48.520 77.420 48.810 ;
        RECT 77.080 48.180 80.140 48.520 ;
        RECT 77.080 47.890 77.420 48.180 ;
        RECT 86.720 47.890 87.060 48.810 ;
        RECT 88.040 47.890 88.380 48.810 ;
        RECT 94.640 47.890 94.980 48.810 ;
        RECT 95.960 47.890 96.300 48.810 ;
        RECT 107.840 47.890 108.180 48.810 ;
        RECT 109.160 47.890 109.500 48.810 ;
        RECT 115.760 47.890 116.100 48.810 ;
        RECT 117.080 47.890 117.420 48.810 ;
        RECT 24.120 44.870 24.460 45.790 ;
        RECT 43.920 44.870 44.260 45.790 ;
        RECT 58.840 45.500 59.180 45.790 ;
        RECT 56.120 45.160 59.180 45.500 ;
        RECT 58.840 44.870 59.180 45.160 ;
        RECT 77.080 45.500 77.420 45.790 ;
        RECT 77.080 45.160 80.140 45.500 ;
        RECT 77.080 44.870 77.420 45.160 ;
        RECT 92.000 44.870 92.340 45.790 ;
        RECT 111.800 44.870 112.140 45.790 ;
        RECT 13.560 41.850 13.900 42.770 ;
        RECT 14.880 41.850 15.220 42.770 ;
        RECT 16.200 41.850 16.540 42.770 ;
        RECT 17.520 41.850 17.860 42.770 ;
        RECT 29.400 41.850 29.740 42.770 ;
        RECT 30.720 41.850 31.060 42.770 ;
        RECT 32.040 41.850 32.380 42.770 ;
        RECT 33.360 41.850 33.700 42.770 ;
        RECT 34.680 41.850 35.020 42.770 ;
        RECT 36.000 41.850 36.340 42.770 ;
        RECT 37.320 41.850 37.660 42.770 ;
        RECT 38.640 41.850 38.980 42.770 ;
        RECT 50.520 41.850 50.860 42.770 ;
        RECT 51.840 41.850 52.180 42.770 ;
        RECT 53.160 41.850 53.500 42.770 ;
        RECT 54.480 41.850 54.820 42.770 ;
        RECT 58.840 42.480 59.180 42.770 ;
        RECT 56.120 42.140 59.180 42.480 ;
        RECT 58.840 41.850 59.180 42.140 ;
        RECT 77.080 42.480 77.420 42.770 ;
        RECT 77.080 42.140 80.140 42.480 ;
        RECT 77.080 41.850 77.420 42.140 ;
        RECT 81.440 41.850 81.780 42.770 ;
        RECT 82.760 41.850 83.100 42.770 ;
        RECT 84.080 41.850 84.420 42.770 ;
        RECT 85.400 41.850 85.740 42.770 ;
        RECT 97.280 41.850 97.620 42.770 ;
        RECT 98.600 41.850 98.940 42.770 ;
        RECT 99.920 41.850 100.260 42.770 ;
        RECT 101.240 41.850 101.580 42.770 ;
        RECT 102.560 41.850 102.900 42.770 ;
        RECT 103.880 41.850 104.220 42.770 ;
        RECT 105.200 41.850 105.540 42.770 ;
        RECT 106.520 41.850 106.860 42.770 ;
        RECT 118.400 41.850 118.740 42.770 ;
        RECT 119.720 41.850 120.060 42.770 ;
        RECT 121.040 41.850 121.380 42.770 ;
        RECT 122.360 41.850 122.700 42.770 ;
        RECT 45.240 38.830 45.580 39.750 ;
        RECT 58.840 39.460 59.180 39.750 ;
        RECT 56.120 39.120 59.180 39.460 ;
        RECT 58.840 38.830 59.180 39.120 ;
        RECT 77.080 39.460 77.420 39.750 ;
        RECT 77.080 39.120 80.140 39.460 ;
        RECT 77.080 38.830 77.420 39.120 ;
        RECT 90.680 38.830 91.020 39.750 ;
        RECT 123.680 38.170 124.020 106.510 ;
        RECT 11.070 36.240 46.710 36.640 ;
        RECT 11.070 35.440 45.990 35.840 ;
        RECT 11.070 34.240 11.430 35.440 ;
        RECT 46.350 35.040 46.710 36.240 ;
        RECT 11.790 34.640 46.710 35.040 ;
        RECT 11.070 33.840 45.990 34.240 ;
        RECT 11.070 32.640 11.430 33.840 ;
        RECT 46.350 33.440 46.710 34.640 ;
        RECT 11.790 33.040 46.710 33.440 ;
        RECT 89.550 36.240 125.190 36.640 ;
        RECT 89.550 35.040 89.910 36.240 ;
        RECT 90.270 35.440 125.190 35.840 ;
        RECT 89.550 34.640 124.470 35.040 ;
        RECT 89.550 33.440 89.910 34.640 ;
        RECT 124.830 34.240 125.190 35.440 ;
        RECT 90.270 33.840 125.190 34.240 ;
        RECT 89.550 33.040 124.470 33.440 ;
        RECT 124.830 32.640 125.190 33.840 ;
        RECT 11.070 32.240 46.710 32.640 ;
        RECT 89.550 32.240 125.190 32.640 ;
        RECT 11.070 31.440 46.710 31.840 ;
        RECT 11.070 30.640 45.990 31.040 ;
        RECT 11.070 29.440 11.430 30.640 ;
        RECT 46.350 30.240 46.710 31.440 ;
        RECT 11.790 29.840 46.710 30.240 ;
        RECT 11.070 29.040 45.990 29.440 ;
        RECT 11.070 27.840 11.430 29.040 ;
        RECT 46.350 28.640 46.710 29.840 ;
        RECT 89.550 31.440 125.190 31.840 ;
        RECT 89.550 30.240 89.910 31.440 ;
        RECT 90.270 30.640 125.190 31.040 ;
        RECT 89.550 29.840 124.470 30.240 ;
        RECT 52.270 29.350 53.190 29.690 ;
        RECT 56.230 29.350 57.150 29.690 ;
        RECT 79.110 29.350 80.030 29.690 ;
        RECT 83.070 29.350 83.990 29.690 ;
        RECT 11.790 28.240 46.710 28.640 ;
        RECT 52.270 28.470 53.190 28.810 ;
        RECT 56.230 28.470 57.150 28.810 ;
        RECT 79.110 28.470 80.030 28.810 ;
        RECT 83.070 28.470 83.990 28.810 ;
        RECT 89.550 28.640 89.910 29.840 ;
        RECT 124.830 29.440 125.190 30.640 ;
        RECT 90.270 29.040 125.190 29.440 ;
        RECT 89.550 28.240 124.470 28.640 ;
        RECT 11.070 27.440 46.710 27.840 ;
        RECT 58.830 27.590 59.750 27.930 ;
        RECT 76.510 27.590 77.430 27.930 ;
        RECT 124.830 27.840 125.190 29.040 ;
        RECT 89.550 27.440 125.190 27.840 ;
        RECT 11.070 26.640 46.710 27.040 ;
        RECT 52.270 26.710 53.190 27.050 ;
        RECT 56.230 26.710 57.150 27.050 ;
        RECT 79.110 26.710 80.030 27.050 ;
        RECT 83.070 26.710 83.990 27.050 ;
        RECT 11.070 25.840 45.990 26.240 ;
        RECT 11.070 24.640 11.430 25.840 ;
        RECT 46.350 25.440 46.710 26.640 ;
        RECT 89.550 26.640 125.190 27.040 ;
        RECT 52.270 25.830 53.190 26.170 ;
        RECT 56.230 25.830 57.150 26.170 ;
        RECT 63.270 25.830 64.990 26.170 ;
        RECT 71.910 25.830 72.830 26.170 ;
        RECT 79.110 25.830 80.030 26.170 ;
        RECT 83.070 25.830 83.990 26.170 ;
        RECT 11.790 25.040 46.710 25.440 ;
        RECT 11.070 24.240 45.990 24.640 ;
        RECT 11.070 23.040 11.430 24.240 ;
        RECT 46.350 23.840 46.710 25.040 ;
        RECT 52.270 24.950 53.190 25.290 ;
        RECT 56.230 24.950 57.150 25.290 ;
        RECT 11.790 23.440 46.710 23.840 ;
        RECT 52.270 23.190 53.190 23.530 ;
        RECT 56.230 23.190 57.150 23.530 ;
        RECT 11.070 22.640 46.710 23.040 ;
        RECT 52.270 22.310 53.190 22.650 ;
        RECT 56.070 22.310 60.970 22.650 ;
        RECT 11.070 21.840 46.710 22.240 ;
        RECT 11.070 21.040 45.990 21.440 ;
        RECT 11.070 19.840 11.430 21.040 ;
        RECT 46.350 20.640 46.710 21.840 ;
        RECT 50.110 21.430 51.030 21.770 ;
        RECT 57.590 20.990 59.310 21.330 ;
        RECT 11.790 20.240 46.710 20.640 ;
        RECT 56.230 20.550 57.150 20.890 ;
        RECT 11.070 19.440 45.990 19.840 ;
        RECT 11.070 18.240 11.430 19.440 ;
        RECT 46.350 19.040 46.710 20.240 ;
        RECT 11.790 18.640 46.710 19.040 ;
        RECT 51.470 18.790 53.190 19.130 ;
        RECT 50.110 18.350 51.030 18.690 ;
        RECT 11.070 17.840 46.710 18.240 ;
        RECT 11.070 17.040 46.710 17.440 ;
        RECT 11.070 16.240 45.990 16.640 ;
        RECT 11.070 15.040 11.430 16.240 ;
        RECT 46.350 15.840 46.710 17.040 ;
        RECT 11.790 15.440 46.710 15.840 ;
        RECT 11.070 14.640 45.990 15.040 ;
        RECT 11.070 13.440 11.430 14.640 ;
        RECT 46.350 14.240 46.710 15.440 ;
        RECT 11.790 13.840 46.710 14.240 ;
        RECT 11.070 13.380 46.710 13.440 ;
        RECT 51.470 13.380 51.810 18.790 ;
        RECT 52.270 17.910 53.190 18.250 ;
        RECT 56.230 17.910 57.150 18.250 ;
        RECT 57.590 16.660 57.930 20.990 ;
        RECT 60.630 17.810 60.970 22.310 ;
        RECT 64.650 19.130 64.990 25.830 ;
        RECT 89.550 25.440 89.910 26.640 ;
        RECT 90.270 25.840 125.190 26.240 ;
        RECT 79.110 24.950 80.030 25.290 ;
        RECT 83.070 24.950 83.990 25.290 ;
        RECT 89.550 25.040 124.470 25.440 ;
        RECT 89.550 23.840 89.910 25.040 ;
        RECT 124.830 24.640 125.190 25.840 ;
        RECT 90.270 24.240 125.190 24.640 ;
        RECT 79.110 23.190 80.030 23.530 ;
        RECT 83.070 23.190 83.990 23.530 ;
        RECT 89.550 23.440 124.470 23.840 ;
        RECT 124.830 23.040 125.190 24.240 ;
        RECT 75.290 22.310 80.190 22.650 ;
        RECT 83.070 22.310 83.990 22.650 ;
        RECT 89.550 22.640 125.190 23.040 ;
        RECT 63.270 18.790 64.190 19.130 ;
        RECT 64.650 18.790 72.830 19.130 ;
        RECT 75.290 17.810 75.630 22.310 ;
        RECT 89.550 21.840 125.190 22.240 ;
        RECT 85.230 21.430 86.150 21.770 ;
        RECT 76.950 20.990 78.670 21.330 ;
        RECT 60.630 17.470 66.350 17.810 ;
        RECT 69.910 17.470 75.630 17.810 ;
        RECT 56.230 16.320 57.930 16.660 ;
        RECT 78.330 16.660 78.670 20.990 ;
        RECT 79.110 20.550 80.030 20.890 ;
        RECT 89.550 20.640 89.910 21.840 ;
        RECT 90.270 21.040 125.190 21.440 ;
        RECT 89.550 20.240 124.470 20.640 ;
        RECT 83.070 18.790 84.790 19.130 ;
        RECT 79.110 17.910 80.030 18.250 ;
        RECT 83.070 17.910 83.990 18.250 ;
        RECT 78.330 16.320 80.030 16.660 ;
        RECT 52.270 15.270 53.190 15.610 ;
        RECT 56.230 15.270 57.150 15.610 ;
        RECT 79.110 15.270 80.030 15.610 ;
        RECT 83.070 15.270 83.990 15.610 ;
        RECT 52.270 14.390 53.190 14.730 ;
        RECT 56.230 14.390 57.150 14.730 ;
        RECT 63.270 14.390 64.190 14.730 ;
        RECT 72.070 14.660 72.990 14.730 ;
        RECT 72.070 14.390 73.090 14.660 ;
        RECT 79.110 14.390 80.030 14.730 ;
        RECT 83.070 14.390 83.990 14.730 ;
        RECT 52.270 13.510 53.190 13.850 ;
        RECT 56.230 13.510 57.150 13.850 ;
        RECT 11.070 13.040 51.810 13.380 ;
        RECT 56.230 9.640 57.150 10.560 ;
        RECT 52.270 6.040 53.190 6.960 ;
        RECT 58.830 3.920 59.750 4.260 ;
        RECT 63.470 2.065 64.070 14.390 ;
        RECT 72.490 2.900 73.090 14.390 ;
        RECT 79.110 13.510 80.030 13.850 ;
        RECT 83.070 13.510 83.990 13.850 ;
        RECT 84.450 13.380 84.790 18.790 ;
        RECT 89.550 19.040 89.910 20.240 ;
        RECT 124.830 19.840 125.190 21.040 ;
        RECT 90.270 19.440 125.190 19.840 ;
        RECT 85.230 18.350 86.150 18.690 ;
        RECT 89.550 18.640 124.470 19.040 ;
        RECT 124.830 18.240 125.190 19.440 ;
        RECT 89.550 17.840 125.190 18.240 ;
        RECT 89.550 17.040 125.190 17.440 ;
        RECT 89.550 15.840 89.910 17.040 ;
        RECT 90.270 16.240 125.190 16.640 ;
        RECT 89.550 15.440 124.470 15.840 ;
        RECT 89.550 14.240 89.910 15.440 ;
        RECT 124.830 15.040 125.190 16.240 ;
        RECT 90.270 14.640 125.190 15.040 ;
        RECT 89.550 13.840 124.470 14.240 ;
        RECT 124.830 13.440 125.190 14.640 ;
        RECT 89.550 13.380 125.190 13.440 ;
        RECT 84.450 13.040 125.190 13.380 ;
        RECT 79.110 9.640 80.030 10.560 ;
        RECT 83.070 6.040 83.990 6.960 ;
        RECT 76.510 3.920 77.430 4.260 ;
        RECT 72.515 2.880 73.065 2.900 ;
        RECT 63.450 1.515 64.090 2.065 ;
        RECT 63.470 1.490 64.070 1.515 ;
      LAYER via2 ;
        RECT 57.515 224.325 57.795 224.605 ;
        RECT 59.705 224.385 59.985 224.665 ;
        RECT 36.010 223.480 36.310 223.780 ;
        RECT 40.860 223.460 41.140 223.740 ;
        RECT 15.760 222.660 16.040 222.940 ;
        RECT 32.360 221.960 32.640 222.240 ;
        RECT 61.630 224.160 61.930 224.460 ;
        RECT 86.890 224.150 87.170 224.430 ;
        RECT 57.560 222.660 57.840 222.940 ;
        RECT 66.060 221.960 66.340 222.240 ;
        RECT 79.425 221.740 79.725 222.040 ;
        RECT 82.660 222.660 82.940 222.940 ;
        RECT 108.060 223.960 108.340 224.240 ;
        RECT 91.260 223.260 91.540 223.540 ;
        RECT 111.340 223.030 111.620 223.310 ;
        RECT 116.170 220.350 116.450 220.630 ;
        RECT 116.690 220.350 116.970 220.630 ;
        RECT 120.130 220.350 120.410 220.630 ;
        RECT 120.650 220.350 120.930 220.630 ;
        RECT 15.370 219.470 15.650 219.750 ;
        RECT 15.890 219.470 16.170 219.750 ;
        RECT 19.330 219.470 19.610 219.750 ;
        RECT 19.850 219.470 20.130 219.750 ;
        RECT 28.130 219.470 28.410 219.750 ;
        RECT 28.650 219.470 28.930 219.750 ;
        RECT 32.090 219.470 32.370 219.750 ;
        RECT 32.610 219.470 32.890 219.750 ;
        RECT 40.570 219.470 40.850 219.750 ;
        RECT 41.090 219.470 41.370 219.750 ;
        RECT 44.530 219.470 44.810 219.750 ;
        RECT 45.050 219.470 45.330 219.750 ;
        RECT 53.330 219.470 53.610 219.750 ;
        RECT 53.850 219.470 54.130 219.750 ;
        RECT 57.290 219.470 57.570 219.750 ;
        RECT 57.810 219.470 58.090 219.750 ;
        RECT 65.770 219.470 66.050 219.750 ;
        RECT 66.290 219.470 66.570 219.750 ;
        RECT 69.730 219.470 70.010 219.750 ;
        RECT 70.250 219.470 70.530 219.750 ;
        RECT 78.530 219.470 78.810 219.750 ;
        RECT 79.050 219.470 79.330 219.750 ;
        RECT 82.490 219.470 82.770 219.750 ;
        RECT 83.010 219.470 83.290 219.750 ;
        RECT 90.970 219.470 91.250 219.750 ;
        RECT 91.490 219.470 91.770 219.750 ;
        RECT 94.930 219.470 95.210 219.750 ;
        RECT 95.450 219.470 95.730 219.750 ;
        RECT 103.730 219.470 104.010 219.750 ;
        RECT 104.250 219.470 104.530 219.750 ;
        RECT 107.690 219.470 107.970 219.750 ;
        RECT 108.210 219.470 108.490 219.750 ;
        RECT 116.170 218.590 116.450 218.870 ;
        RECT 116.690 218.590 116.970 218.870 ;
        RECT 120.130 218.590 120.410 218.870 ;
        RECT 120.650 218.590 120.930 218.870 ;
        RECT 120.130 217.710 120.410 217.990 ;
        RECT 120.650 217.710 120.930 217.990 ;
        RECT 15.370 216.830 15.650 217.110 ;
        RECT 15.890 216.830 16.170 217.110 ;
        RECT 19.330 216.830 19.610 217.110 ;
        RECT 19.850 216.830 20.130 217.110 ;
        RECT 28.130 216.830 28.410 217.110 ;
        RECT 28.650 216.830 28.930 217.110 ;
        RECT 32.090 216.830 32.370 217.110 ;
        RECT 32.610 216.830 32.890 217.110 ;
        RECT 40.570 216.830 40.850 217.110 ;
        RECT 41.090 216.830 41.370 217.110 ;
        RECT 44.530 216.830 44.810 217.110 ;
        RECT 45.050 216.830 45.330 217.110 ;
        RECT 53.330 216.830 53.610 217.110 ;
        RECT 53.850 216.830 54.130 217.110 ;
        RECT 57.290 216.830 57.570 217.110 ;
        RECT 57.810 216.830 58.090 217.110 ;
        RECT 65.770 216.830 66.050 217.110 ;
        RECT 66.290 216.830 66.570 217.110 ;
        RECT 69.730 216.830 70.010 217.110 ;
        RECT 70.250 216.830 70.530 217.110 ;
        RECT 78.530 216.830 78.810 217.110 ;
        RECT 79.050 216.830 79.330 217.110 ;
        RECT 82.490 216.830 82.770 217.110 ;
        RECT 83.010 216.830 83.290 217.110 ;
        RECT 90.970 216.830 91.250 217.110 ;
        RECT 91.490 216.830 91.770 217.110 ;
        RECT 94.930 216.830 95.210 217.110 ;
        RECT 95.450 216.830 95.730 217.110 ;
        RECT 103.730 216.830 104.010 217.110 ;
        RECT 104.250 216.830 104.530 217.110 ;
        RECT 107.690 216.830 107.970 217.110 ;
        RECT 108.210 216.830 108.490 217.110 ;
        RECT 15.370 214.190 15.650 214.470 ;
        RECT 15.890 214.190 16.170 214.470 ;
        RECT 19.330 214.190 19.610 214.470 ;
        RECT 19.850 214.190 20.130 214.470 ;
        RECT 28.130 214.190 28.410 214.470 ;
        RECT 28.650 214.190 28.930 214.470 ;
        RECT 32.090 214.190 32.370 214.470 ;
        RECT 32.610 214.190 32.890 214.470 ;
        RECT 40.570 214.190 40.850 214.470 ;
        RECT 41.090 214.190 41.370 214.470 ;
        RECT 44.530 214.190 44.810 214.470 ;
        RECT 45.050 214.190 45.330 214.470 ;
        RECT 53.330 214.190 53.610 214.470 ;
        RECT 53.850 214.190 54.130 214.470 ;
        RECT 57.290 214.190 57.570 214.470 ;
        RECT 57.810 214.190 58.090 214.470 ;
        RECT 65.770 214.190 66.050 214.470 ;
        RECT 66.290 214.190 66.570 214.470 ;
        RECT 69.730 214.190 70.010 214.470 ;
        RECT 70.250 214.190 70.530 214.470 ;
        RECT 78.530 214.190 78.810 214.470 ;
        RECT 79.050 214.190 79.330 214.470 ;
        RECT 82.490 214.190 82.770 214.470 ;
        RECT 83.010 214.190 83.290 214.470 ;
        RECT 90.970 214.190 91.250 214.470 ;
        RECT 91.490 214.190 91.770 214.470 ;
        RECT 94.930 214.190 95.210 214.470 ;
        RECT 95.450 214.190 95.730 214.470 ;
        RECT 103.730 214.190 104.010 214.470 ;
        RECT 104.250 214.190 104.530 214.470 ;
        RECT 107.690 214.190 107.970 214.470 ;
        RECT 108.210 214.190 108.490 214.470 ;
        RECT 15.370 212.430 15.650 212.710 ;
        RECT 15.890 212.430 16.170 212.710 ;
        RECT 19.330 212.430 19.610 212.710 ;
        RECT 19.850 212.430 20.130 212.710 ;
        RECT 28.130 212.430 28.410 212.710 ;
        RECT 28.650 212.430 28.930 212.710 ;
        RECT 32.090 212.430 32.370 212.710 ;
        RECT 32.610 212.430 32.890 212.710 ;
        RECT 40.570 212.430 40.850 212.710 ;
        RECT 41.090 212.430 41.370 212.710 ;
        RECT 44.530 212.430 44.810 212.710 ;
        RECT 45.050 212.430 45.330 212.710 ;
        RECT 53.330 212.430 53.610 212.710 ;
        RECT 53.850 212.430 54.130 212.710 ;
        RECT 57.290 212.430 57.570 212.710 ;
        RECT 57.810 212.430 58.090 212.710 ;
        RECT 65.770 212.430 66.050 212.710 ;
        RECT 66.290 212.430 66.570 212.710 ;
        RECT 69.730 212.430 70.010 212.710 ;
        RECT 70.250 212.430 70.530 212.710 ;
        RECT 78.530 212.430 78.810 212.710 ;
        RECT 79.050 212.430 79.330 212.710 ;
        RECT 82.490 212.430 82.770 212.710 ;
        RECT 83.010 212.430 83.290 212.710 ;
        RECT 90.970 212.430 91.250 212.710 ;
        RECT 91.490 212.430 91.770 212.710 ;
        RECT 94.930 212.430 95.210 212.710 ;
        RECT 95.450 212.430 95.730 212.710 ;
        RECT 103.730 212.430 104.010 212.710 ;
        RECT 104.250 212.430 104.530 212.710 ;
        RECT 107.690 212.430 107.970 212.710 ;
        RECT 108.210 212.430 108.490 212.710 ;
        RECT 116.170 215.950 116.450 216.230 ;
        RECT 116.690 215.950 116.970 216.230 ;
        RECT 120.130 215.950 120.410 216.230 ;
        RECT 120.650 215.950 120.930 216.230 ;
        RECT 130.755 215.055 131.045 215.345 ;
        RECT 116.170 214.190 116.450 214.470 ;
        RECT 116.690 214.190 116.970 214.470 ;
        RECT 120.130 214.190 120.410 214.470 ;
        RECT 120.650 214.190 120.930 214.470 ;
        RECT 116.170 212.430 116.450 212.710 ;
        RECT 116.690 212.430 116.970 212.710 ;
        RECT 120.130 212.430 120.410 212.710 ;
        RECT 120.650 212.430 120.930 212.710 ;
        RECT 116.170 211.550 116.450 211.830 ;
        RECT 116.690 211.550 116.970 211.830 ;
        RECT 15.370 209.790 15.650 210.070 ;
        RECT 15.890 209.790 16.170 210.070 ;
        RECT 19.330 209.790 19.610 210.070 ;
        RECT 19.850 209.790 20.130 210.070 ;
        RECT 28.130 209.790 28.410 210.070 ;
        RECT 28.650 209.790 28.930 210.070 ;
        RECT 32.090 209.790 32.370 210.070 ;
        RECT 32.610 209.790 32.890 210.070 ;
        RECT 40.570 209.790 40.850 210.070 ;
        RECT 41.090 209.790 41.370 210.070 ;
        RECT 44.530 209.790 44.810 210.070 ;
        RECT 45.050 209.790 45.330 210.070 ;
        RECT 53.330 209.790 53.610 210.070 ;
        RECT 53.850 209.790 54.130 210.070 ;
        RECT 57.290 209.790 57.570 210.070 ;
        RECT 57.810 209.790 58.090 210.070 ;
        RECT 65.770 209.790 66.050 210.070 ;
        RECT 66.290 209.790 66.570 210.070 ;
        RECT 69.730 209.790 70.010 210.070 ;
        RECT 70.250 209.790 70.530 210.070 ;
        RECT 78.530 209.790 78.810 210.070 ;
        RECT 79.050 209.790 79.330 210.070 ;
        RECT 82.490 209.790 82.770 210.070 ;
        RECT 83.010 209.790 83.290 210.070 ;
        RECT 90.970 209.790 91.250 210.070 ;
        RECT 91.490 209.790 91.770 210.070 ;
        RECT 94.930 209.790 95.210 210.070 ;
        RECT 95.450 209.790 95.730 210.070 ;
        RECT 103.730 209.790 104.010 210.070 ;
        RECT 104.250 209.790 104.530 210.070 ;
        RECT 107.690 209.790 107.970 210.070 ;
        RECT 108.210 209.790 108.490 210.070 ;
        RECT 116.170 209.790 116.450 210.070 ;
        RECT 116.690 209.790 116.970 210.070 ;
        RECT 120.130 209.790 120.410 210.070 ;
        RECT 120.650 209.790 120.930 210.070 ;
        RECT 116.170 208.030 116.450 208.310 ;
        RECT 116.690 208.030 116.970 208.310 ;
        RECT 120.130 208.030 120.410 208.310 ;
        RECT 120.650 208.030 120.930 208.310 ;
        RECT 114.010 207.590 114.290 207.870 ;
        RECT 114.530 207.590 114.810 207.870 ;
        RECT 15.370 207.150 15.650 207.430 ;
        RECT 15.890 207.150 16.170 207.430 ;
        RECT 19.330 207.150 19.610 207.430 ;
        RECT 19.850 207.150 20.130 207.430 ;
        RECT 28.130 207.150 28.410 207.430 ;
        RECT 28.650 207.150 28.930 207.430 ;
        RECT 32.090 207.150 32.370 207.430 ;
        RECT 32.610 207.150 32.890 207.430 ;
        RECT 15.370 205.390 15.650 205.670 ;
        RECT 15.890 205.390 16.170 205.670 ;
        RECT 19.330 205.390 19.610 205.670 ;
        RECT 19.850 205.390 20.130 205.670 ;
        RECT 28.130 205.390 28.410 205.670 ;
        RECT 28.650 205.390 28.930 205.670 ;
        RECT 32.090 205.390 32.370 205.670 ;
        RECT 32.610 205.390 32.890 205.670 ;
        RECT 15.370 203.630 15.650 203.910 ;
        RECT 15.890 203.630 16.170 203.910 ;
        RECT 19.330 203.630 19.610 203.910 ;
        RECT 19.850 203.630 20.130 203.910 ;
        RECT 28.130 203.630 28.410 203.910 ;
        RECT 28.650 203.630 28.930 203.910 ;
        RECT 32.090 203.630 32.370 203.910 ;
        RECT 32.610 203.630 32.890 203.910 ;
        RECT 15.370 202.750 15.650 203.030 ;
        RECT 15.890 202.750 16.170 203.030 ;
        RECT 19.330 202.750 19.610 203.030 ;
        RECT 19.850 202.750 20.130 203.030 ;
        RECT 28.130 202.750 28.410 203.030 ;
        RECT 28.650 202.750 28.930 203.030 ;
        RECT 32.090 202.750 32.370 203.030 ;
        RECT 32.610 202.750 32.890 203.030 ;
        RECT 15.370 201.870 15.650 202.150 ;
        RECT 15.890 201.870 16.170 202.150 ;
        RECT 19.330 201.870 19.610 202.150 ;
        RECT 19.850 201.870 20.130 202.150 ;
        RECT 28.130 201.870 28.410 202.150 ;
        RECT 28.650 201.870 28.930 202.150 ;
        RECT 32.090 201.870 32.370 202.150 ;
        RECT 32.610 201.870 32.890 202.150 ;
        RECT 15.370 199.650 15.650 199.930 ;
        RECT 15.890 199.650 16.170 199.930 ;
        RECT 15.370 199.130 15.650 199.410 ;
        RECT 15.890 199.130 16.170 199.410 ;
        RECT 32.090 199.650 32.370 199.930 ;
        RECT 32.610 199.650 32.890 199.930 ;
        RECT 32.090 199.130 32.370 199.410 ;
        RECT 32.610 199.130 32.890 199.410 ;
        RECT 19.330 198.210 19.610 198.490 ;
        RECT 19.850 198.210 20.130 198.490 ;
        RECT 13.230 197.650 13.530 197.950 ;
        RECT 19.330 197.690 19.610 197.970 ;
        RECT 19.850 197.690 20.130 197.970 ;
        RECT 22.110 198.210 22.390 198.490 ;
        RECT 22.630 198.210 22.910 198.490 ;
        RECT 22.110 197.690 22.390 197.970 ;
        RECT 22.630 197.690 22.910 197.970 ;
        RECT 25.150 198.210 25.430 198.490 ;
        RECT 25.670 198.210 25.950 198.490 ;
        RECT 25.150 197.690 25.430 197.970 ;
        RECT 25.670 197.690 25.950 197.970 ;
        RECT 28.130 198.210 28.410 198.490 ;
        RECT 28.650 198.210 28.930 198.490 ;
        RECT 40.570 207.150 40.850 207.430 ;
        RECT 41.090 207.150 41.370 207.430 ;
        RECT 44.530 207.150 44.810 207.430 ;
        RECT 45.050 207.150 45.330 207.430 ;
        RECT 53.330 207.150 53.610 207.430 ;
        RECT 53.850 207.150 54.130 207.430 ;
        RECT 57.290 207.150 57.570 207.430 ;
        RECT 57.810 207.150 58.090 207.430 ;
        RECT 40.570 205.390 40.850 205.670 ;
        RECT 41.090 205.390 41.370 205.670 ;
        RECT 44.530 205.390 44.810 205.670 ;
        RECT 45.050 205.390 45.330 205.670 ;
        RECT 53.330 205.390 53.610 205.670 ;
        RECT 53.850 205.390 54.130 205.670 ;
        RECT 57.290 205.390 57.570 205.670 ;
        RECT 57.810 205.390 58.090 205.670 ;
        RECT 40.570 203.630 40.850 203.910 ;
        RECT 41.090 203.630 41.370 203.910 ;
        RECT 44.530 203.630 44.810 203.910 ;
        RECT 45.050 203.630 45.330 203.910 ;
        RECT 53.330 203.630 53.610 203.910 ;
        RECT 53.850 203.630 54.130 203.910 ;
        RECT 57.290 203.630 57.570 203.910 ;
        RECT 57.810 203.630 58.090 203.910 ;
        RECT 40.570 202.750 40.850 203.030 ;
        RECT 41.090 202.750 41.370 203.030 ;
        RECT 44.530 202.750 44.810 203.030 ;
        RECT 45.050 202.750 45.330 203.030 ;
        RECT 53.330 202.750 53.610 203.030 ;
        RECT 53.850 202.750 54.130 203.030 ;
        RECT 57.290 202.750 57.570 203.030 ;
        RECT 57.810 202.750 58.090 203.030 ;
        RECT 40.570 201.870 40.850 202.150 ;
        RECT 41.090 201.870 41.370 202.150 ;
        RECT 44.530 201.870 44.810 202.150 ;
        RECT 45.050 201.870 45.330 202.150 ;
        RECT 53.330 201.870 53.610 202.150 ;
        RECT 53.850 201.870 54.130 202.150 ;
        RECT 57.290 201.870 57.570 202.150 ;
        RECT 57.810 201.870 58.090 202.150 ;
        RECT 40.570 199.650 40.850 199.930 ;
        RECT 41.090 199.650 41.370 199.930 ;
        RECT 40.570 199.130 40.850 199.410 ;
        RECT 41.090 199.130 41.370 199.410 ;
        RECT 57.290 199.650 57.570 199.930 ;
        RECT 57.810 199.650 58.090 199.930 ;
        RECT 57.290 199.130 57.570 199.410 ;
        RECT 57.810 199.130 58.090 199.410 ;
        RECT 44.530 198.210 44.810 198.490 ;
        RECT 45.050 198.210 45.330 198.490 ;
        RECT 28.130 197.690 28.410 197.970 ;
        RECT 28.650 197.690 28.930 197.970 ;
        RECT 34.355 197.655 34.645 197.945 ;
        RECT 38.855 197.555 39.145 197.845 ;
        RECT 44.530 197.690 44.810 197.970 ;
        RECT 45.050 197.690 45.330 197.970 ;
        RECT 47.310 198.210 47.590 198.490 ;
        RECT 47.830 198.210 48.110 198.490 ;
        RECT 47.310 197.690 47.590 197.970 ;
        RECT 47.830 197.690 48.110 197.970 ;
        RECT 50.350 198.210 50.630 198.490 ;
        RECT 50.870 198.210 51.150 198.490 ;
        RECT 50.350 197.690 50.630 197.970 ;
        RECT 50.870 197.690 51.150 197.970 ;
        RECT 53.330 198.210 53.610 198.490 ;
        RECT 53.850 198.210 54.130 198.490 ;
        RECT 65.770 207.150 66.050 207.430 ;
        RECT 66.290 207.150 66.570 207.430 ;
        RECT 69.730 207.150 70.010 207.430 ;
        RECT 70.250 207.150 70.530 207.430 ;
        RECT 78.530 207.150 78.810 207.430 ;
        RECT 79.050 207.150 79.330 207.430 ;
        RECT 82.490 207.150 82.770 207.430 ;
        RECT 83.010 207.150 83.290 207.430 ;
        RECT 65.770 205.390 66.050 205.670 ;
        RECT 66.290 205.390 66.570 205.670 ;
        RECT 69.730 205.390 70.010 205.670 ;
        RECT 70.250 205.390 70.530 205.670 ;
        RECT 78.530 205.390 78.810 205.670 ;
        RECT 79.050 205.390 79.330 205.670 ;
        RECT 82.490 205.390 82.770 205.670 ;
        RECT 83.010 205.390 83.290 205.670 ;
        RECT 65.770 203.630 66.050 203.910 ;
        RECT 66.290 203.630 66.570 203.910 ;
        RECT 69.730 203.630 70.010 203.910 ;
        RECT 70.250 203.630 70.530 203.910 ;
        RECT 78.530 203.630 78.810 203.910 ;
        RECT 79.050 203.630 79.330 203.910 ;
        RECT 82.490 203.630 82.770 203.910 ;
        RECT 83.010 203.630 83.290 203.910 ;
        RECT 65.770 202.750 66.050 203.030 ;
        RECT 66.290 202.750 66.570 203.030 ;
        RECT 69.730 202.750 70.010 203.030 ;
        RECT 70.250 202.750 70.530 203.030 ;
        RECT 78.530 202.750 78.810 203.030 ;
        RECT 79.050 202.750 79.330 203.030 ;
        RECT 82.490 202.750 82.770 203.030 ;
        RECT 83.010 202.750 83.290 203.030 ;
        RECT 65.770 201.870 66.050 202.150 ;
        RECT 66.290 201.870 66.570 202.150 ;
        RECT 69.730 201.870 70.010 202.150 ;
        RECT 70.250 201.870 70.530 202.150 ;
        RECT 78.530 201.870 78.810 202.150 ;
        RECT 79.050 201.870 79.330 202.150 ;
        RECT 82.490 201.870 82.770 202.150 ;
        RECT 83.010 201.870 83.290 202.150 ;
        RECT 65.770 199.650 66.050 199.930 ;
        RECT 66.290 199.650 66.570 199.930 ;
        RECT 65.770 199.130 66.050 199.410 ;
        RECT 66.290 199.130 66.570 199.410 ;
        RECT 82.490 199.650 82.770 199.930 ;
        RECT 83.010 199.650 83.290 199.930 ;
        RECT 82.490 199.130 82.770 199.410 ;
        RECT 83.010 199.130 83.290 199.410 ;
        RECT 69.730 198.210 70.010 198.490 ;
        RECT 70.250 198.210 70.530 198.490 ;
        RECT 53.330 197.690 53.610 197.970 ;
        RECT 53.850 197.690 54.130 197.970 ;
        RECT 59.655 197.755 59.945 198.045 ;
        RECT 63.955 197.755 64.245 198.045 ;
        RECT 69.730 197.690 70.010 197.970 ;
        RECT 70.250 197.690 70.530 197.970 ;
        RECT 72.510 198.210 72.790 198.490 ;
        RECT 73.030 198.210 73.310 198.490 ;
        RECT 72.510 197.690 72.790 197.970 ;
        RECT 73.030 197.690 73.310 197.970 ;
        RECT 75.550 198.210 75.830 198.490 ;
        RECT 76.070 198.210 76.350 198.490 ;
        RECT 75.550 197.690 75.830 197.970 ;
        RECT 76.070 197.690 76.350 197.970 ;
        RECT 78.530 198.210 78.810 198.490 ;
        RECT 79.050 198.210 79.330 198.490 ;
        RECT 90.970 207.150 91.250 207.430 ;
        RECT 91.490 207.150 91.770 207.430 ;
        RECT 94.930 207.150 95.210 207.430 ;
        RECT 95.450 207.150 95.730 207.430 ;
        RECT 103.730 207.150 104.010 207.430 ;
        RECT 104.250 207.150 104.530 207.430 ;
        RECT 107.690 207.150 107.970 207.430 ;
        RECT 108.210 207.150 108.490 207.430 ;
        RECT 90.970 205.390 91.250 205.670 ;
        RECT 91.490 205.390 91.770 205.670 ;
        RECT 94.930 205.390 95.210 205.670 ;
        RECT 95.450 205.390 95.730 205.670 ;
        RECT 103.730 205.390 104.010 205.670 ;
        RECT 104.250 205.390 104.530 205.670 ;
        RECT 107.690 205.390 107.970 205.670 ;
        RECT 108.210 205.390 108.490 205.670 ;
        RECT 90.970 203.630 91.250 203.910 ;
        RECT 91.490 203.630 91.770 203.910 ;
        RECT 94.930 203.630 95.210 203.910 ;
        RECT 95.450 203.630 95.730 203.910 ;
        RECT 103.730 203.630 104.010 203.910 ;
        RECT 104.250 203.630 104.530 203.910 ;
        RECT 107.690 203.630 107.970 203.910 ;
        RECT 108.210 203.630 108.490 203.910 ;
        RECT 90.970 202.750 91.250 203.030 ;
        RECT 91.490 202.750 91.770 203.030 ;
        RECT 94.930 202.750 95.210 203.030 ;
        RECT 95.450 202.750 95.730 203.030 ;
        RECT 103.730 202.750 104.010 203.030 ;
        RECT 104.250 202.750 104.530 203.030 ;
        RECT 107.690 202.750 107.970 203.030 ;
        RECT 108.210 202.750 108.490 203.030 ;
        RECT 90.970 201.870 91.250 202.150 ;
        RECT 91.490 201.870 91.770 202.150 ;
        RECT 94.930 201.870 95.210 202.150 ;
        RECT 95.450 201.870 95.730 202.150 ;
        RECT 103.730 201.870 104.010 202.150 ;
        RECT 104.250 201.870 104.530 202.150 ;
        RECT 107.690 201.870 107.970 202.150 ;
        RECT 108.210 201.870 108.490 202.150 ;
        RECT 90.970 199.650 91.250 199.930 ;
        RECT 91.490 199.650 91.770 199.930 ;
        RECT 90.970 199.130 91.250 199.410 ;
        RECT 91.490 199.130 91.770 199.410 ;
        RECT 107.690 199.650 107.970 199.930 ;
        RECT 108.210 199.650 108.490 199.930 ;
        RECT 107.690 199.130 107.970 199.410 ;
        RECT 108.210 199.130 108.490 199.410 ;
        RECT 94.930 198.210 95.210 198.490 ;
        RECT 95.450 198.210 95.730 198.490 ;
        RECT 78.530 197.690 78.810 197.970 ;
        RECT 79.050 197.690 79.330 197.970 ;
        RECT 84.755 197.755 85.045 198.045 ;
        RECT 89.155 197.755 89.445 198.045 ;
        RECT 94.930 197.690 95.210 197.970 ;
        RECT 95.450 197.690 95.730 197.970 ;
        RECT 97.710 198.210 97.990 198.490 ;
        RECT 98.230 198.210 98.510 198.490 ;
        RECT 97.710 197.690 97.990 197.970 ;
        RECT 98.230 197.690 98.510 197.970 ;
        RECT 100.750 198.210 101.030 198.490 ;
        RECT 101.270 198.210 101.550 198.490 ;
        RECT 100.750 197.690 101.030 197.970 ;
        RECT 101.270 197.690 101.550 197.970 ;
        RECT 103.730 198.210 104.010 198.490 ;
        RECT 104.250 198.210 104.530 198.490 ;
        RECT 140.095 206.345 140.415 206.665 ;
        RECT 140.655 206.345 140.975 206.665 ;
        RECT 144.055 206.345 144.375 206.665 ;
        RECT 144.615 206.345 144.935 206.665 ;
        RECT 116.170 205.390 116.450 205.670 ;
        RECT 116.690 205.390 116.970 205.670 ;
        RECT 120.130 205.390 120.410 205.670 ;
        RECT 120.650 205.390 120.930 205.670 ;
        RECT 140.095 205.465 140.415 205.785 ;
        RECT 140.655 205.465 140.975 205.785 ;
        RECT 144.055 205.465 144.375 205.785 ;
        RECT 144.615 205.465 144.935 205.785 ;
        RECT 114.170 204.070 114.450 204.350 ;
        RECT 114.690 204.070 114.970 204.350 ;
        RECT 116.170 203.630 116.450 203.910 ;
        RECT 116.690 203.630 116.970 203.910 ;
        RECT 120.130 203.630 120.410 203.910 ;
        RECT 120.650 203.630 120.930 203.910 ;
        RECT 140.095 203.705 140.415 204.025 ;
        RECT 140.655 203.705 140.975 204.025 ;
        RECT 144.055 203.705 144.375 204.025 ;
        RECT 144.615 203.705 144.935 204.025 ;
        RECT 116.170 202.750 116.450 203.030 ;
        RECT 116.690 202.750 116.970 203.030 ;
        RECT 120.130 202.750 120.410 203.030 ;
        RECT 120.650 202.750 120.930 203.030 ;
        RECT 116.170 201.870 116.450 202.150 ;
        RECT 116.690 201.870 116.970 202.150 ;
        RECT 120.130 201.870 120.410 202.150 ;
        RECT 120.650 201.870 120.930 202.150 ;
        RECT 140.095 201.945 140.415 202.265 ;
        RECT 140.655 201.945 140.975 202.265 ;
        RECT 144.055 201.945 144.375 202.265 ;
        RECT 144.615 201.945 144.935 202.265 ;
        RECT 140.095 201.065 140.415 201.385 ;
        RECT 140.655 201.065 140.975 201.385 ;
        RECT 144.055 201.065 144.375 201.385 ;
        RECT 144.615 201.065 144.935 201.385 ;
        RECT 116.170 199.650 116.450 199.930 ;
        RECT 116.690 199.650 116.970 199.930 ;
        RECT 111.855 199.155 112.145 199.445 ;
        RECT 116.170 199.130 116.450 199.410 ;
        RECT 116.690 199.130 116.970 199.410 ;
        RECT 120.130 198.210 120.410 198.490 ;
        RECT 120.650 198.210 120.930 198.490 ;
        RECT 103.730 197.690 104.010 197.970 ;
        RECT 104.250 197.690 104.530 197.970 ;
        RECT 109.955 197.655 110.245 197.945 ;
        RECT 120.130 197.690 120.410 197.970 ;
        RECT 120.650 197.690 120.930 197.970 ;
        RECT 114.255 196.755 114.545 197.045 ;
        RECT 147.530 196.730 147.870 197.070 ;
        RECT 102.575 195.755 102.865 196.045 ;
        RECT 130.730 195.730 131.070 196.070 ;
        RECT 31.080 195.255 31.370 195.545 ;
        RECT 34.330 195.230 34.670 195.570 ;
        RECT 38.830 195.230 39.170 195.570 ;
        RECT 41.885 195.255 42.175 195.545 ;
        RECT 56.280 195.155 56.570 195.445 ;
        RECT 59.630 195.130 59.970 195.470 ;
        RECT 63.930 195.130 64.270 195.470 ;
        RECT 67.085 195.155 67.375 195.445 ;
        RECT 81.430 195.230 81.770 195.570 ;
        RECT 84.755 195.255 85.045 195.545 ;
        RECT 92.285 195.155 92.575 195.445 ;
        RECT 19.230 194.610 19.510 194.890 ;
        RECT 19.750 194.610 20.030 194.890 ;
        RECT 19.230 194.090 19.510 194.370 ;
        RECT 19.750 194.090 20.030 194.370 ;
        RECT 28.030 194.610 28.310 194.890 ;
        RECT 28.550 194.610 28.830 194.890 ;
        RECT 28.030 194.090 28.310 194.370 ;
        RECT 28.550 194.090 28.830 194.370 ;
        RECT 44.430 194.610 44.710 194.890 ;
        RECT 44.950 194.610 45.230 194.890 ;
        RECT 44.430 194.090 44.710 194.370 ;
        RECT 44.950 194.090 45.230 194.370 ;
        RECT 53.230 194.610 53.510 194.890 ;
        RECT 53.750 194.610 54.030 194.890 ;
        RECT 53.230 194.090 53.510 194.370 ;
        RECT 53.750 194.090 54.030 194.370 ;
        RECT 69.630 194.610 69.910 194.890 ;
        RECT 70.150 194.610 70.430 194.890 ;
        RECT 69.630 194.090 69.910 194.370 ;
        RECT 70.150 194.090 70.430 194.370 ;
        RECT 78.430 194.610 78.710 194.890 ;
        RECT 78.950 194.610 79.230 194.890 ;
        RECT 78.430 194.090 78.710 194.370 ;
        RECT 78.950 194.090 79.230 194.370 ;
        RECT 94.830 194.610 95.110 194.890 ;
        RECT 95.350 194.610 95.630 194.890 ;
        RECT 94.830 194.090 95.110 194.370 ;
        RECT 95.350 194.090 95.630 194.370 ;
        RECT 103.630 194.610 103.910 194.890 ;
        RECT 104.150 194.610 104.430 194.890 ;
        RECT 103.630 194.090 103.910 194.370 ;
        RECT 104.150 194.090 104.430 194.370 ;
        RECT 120.030 194.610 120.310 194.890 ;
        RECT 120.550 194.610 120.830 194.890 ;
        RECT 120.030 194.090 120.310 194.370 ;
        RECT 120.550 194.090 120.830 194.370 ;
        RECT 15.270 191.010 15.550 191.290 ;
        RECT 15.790 191.010 16.070 191.290 ;
        RECT 15.270 190.490 15.550 190.770 ;
        RECT 15.790 190.490 16.070 190.770 ;
        RECT 31.990 191.010 32.270 191.290 ;
        RECT 32.510 191.010 32.790 191.290 ;
        RECT 31.990 190.490 32.270 190.770 ;
        RECT 32.510 190.490 32.790 190.770 ;
        RECT 40.470 191.010 40.750 191.290 ;
        RECT 40.990 191.010 41.270 191.290 ;
        RECT 40.470 190.490 40.750 190.770 ;
        RECT 40.990 190.490 41.270 190.770 ;
        RECT 57.190 191.010 57.470 191.290 ;
        RECT 57.710 191.010 57.990 191.290 ;
        RECT 57.190 190.490 57.470 190.770 ;
        RECT 57.710 190.490 57.990 190.770 ;
        RECT 65.670 191.010 65.950 191.290 ;
        RECT 66.190 191.010 66.470 191.290 ;
        RECT 65.670 190.490 65.950 190.770 ;
        RECT 66.190 190.490 66.470 190.770 ;
        RECT 82.390 191.010 82.670 191.290 ;
        RECT 82.910 191.010 83.190 191.290 ;
        RECT 82.390 190.490 82.670 190.770 ;
        RECT 82.910 190.490 83.190 190.770 ;
        RECT 90.870 191.010 91.150 191.290 ;
        RECT 91.390 191.010 91.670 191.290 ;
        RECT 90.870 190.490 91.150 190.770 ;
        RECT 91.390 190.490 91.670 190.770 ;
        RECT 107.590 191.010 107.870 191.290 ;
        RECT 108.110 191.010 108.390 191.290 ;
        RECT 107.590 190.490 107.870 190.770 ;
        RECT 108.110 190.490 108.390 190.770 ;
        RECT 116.070 191.010 116.350 191.290 ;
        RECT 116.590 191.010 116.870 191.290 ;
        RECT 116.070 190.490 116.350 190.770 ;
        RECT 116.590 190.490 116.870 190.770 ;
        RECT 15.270 187.170 15.550 187.450 ;
        RECT 15.790 187.170 16.070 187.450 ;
        RECT 19.230 187.170 19.510 187.450 ;
        RECT 19.750 187.170 20.030 187.450 ;
        RECT 28.030 187.170 28.310 187.450 ;
        RECT 28.550 187.170 28.830 187.450 ;
        RECT 31.990 187.170 32.270 187.450 ;
        RECT 32.510 187.170 32.790 187.450 ;
        RECT 40.470 187.170 40.750 187.450 ;
        RECT 40.990 187.170 41.270 187.450 ;
        RECT 44.430 187.170 44.710 187.450 ;
        RECT 44.950 187.170 45.230 187.450 ;
        RECT 53.230 187.170 53.510 187.450 ;
        RECT 53.750 187.170 54.030 187.450 ;
        RECT 57.190 187.170 57.470 187.450 ;
        RECT 57.710 187.170 57.990 187.450 ;
        RECT 65.670 187.170 65.950 187.450 ;
        RECT 66.190 187.170 66.470 187.450 ;
        RECT 69.630 187.170 69.910 187.450 ;
        RECT 70.150 187.170 70.430 187.450 ;
        RECT 78.430 187.170 78.710 187.450 ;
        RECT 78.950 187.170 79.230 187.450 ;
        RECT 82.390 187.170 82.670 187.450 ;
        RECT 82.910 187.170 83.190 187.450 ;
        RECT 90.870 187.170 91.150 187.450 ;
        RECT 91.390 187.170 91.670 187.450 ;
        RECT 94.830 187.170 95.110 187.450 ;
        RECT 95.350 187.170 95.630 187.450 ;
        RECT 103.630 187.170 103.910 187.450 ;
        RECT 104.150 187.170 104.430 187.450 ;
        RECT 107.590 187.170 107.870 187.450 ;
        RECT 108.110 187.170 108.390 187.450 ;
        RECT 15.270 186.290 15.550 186.570 ;
        RECT 15.790 186.290 16.070 186.570 ;
        RECT 19.230 186.290 19.510 186.570 ;
        RECT 19.750 186.290 20.030 186.570 ;
        RECT 28.030 186.290 28.310 186.570 ;
        RECT 28.550 186.290 28.830 186.570 ;
        RECT 31.990 186.290 32.270 186.570 ;
        RECT 32.510 186.290 32.790 186.570 ;
        RECT 40.470 186.290 40.750 186.570 ;
        RECT 40.990 186.290 41.270 186.570 ;
        RECT 44.430 186.290 44.710 186.570 ;
        RECT 44.950 186.290 45.230 186.570 ;
        RECT 53.230 186.290 53.510 186.570 ;
        RECT 53.750 186.290 54.030 186.570 ;
        RECT 57.190 186.290 57.470 186.570 ;
        RECT 57.710 186.290 57.990 186.570 ;
        RECT 65.670 186.290 65.950 186.570 ;
        RECT 66.190 186.290 66.470 186.570 ;
        RECT 69.630 186.290 69.910 186.570 ;
        RECT 70.150 186.290 70.430 186.570 ;
        RECT 78.430 186.290 78.710 186.570 ;
        RECT 78.950 186.290 79.230 186.570 ;
        RECT 82.390 186.290 82.670 186.570 ;
        RECT 82.910 186.290 83.190 186.570 ;
        RECT 90.870 186.290 91.150 186.570 ;
        RECT 91.390 186.290 91.670 186.570 ;
        RECT 94.830 186.290 95.110 186.570 ;
        RECT 95.350 186.290 95.630 186.570 ;
        RECT 103.630 186.290 103.910 186.570 ;
        RECT 104.150 186.290 104.430 186.570 ;
        RECT 107.590 186.290 107.870 186.570 ;
        RECT 108.110 186.290 108.390 186.570 ;
        RECT 15.270 184.530 15.550 184.810 ;
        RECT 15.790 184.530 16.070 184.810 ;
        RECT 19.230 184.530 19.510 184.810 ;
        RECT 19.750 184.530 20.030 184.810 ;
        RECT 15.270 183.650 15.550 183.930 ;
        RECT 15.790 183.650 16.070 183.930 ;
        RECT 28.030 184.530 28.310 184.810 ;
        RECT 28.550 184.530 28.830 184.810 ;
        RECT 31.990 184.530 32.270 184.810 ;
        RECT 32.510 184.530 32.790 184.810 ;
        RECT 40.470 184.530 40.750 184.810 ;
        RECT 40.990 184.530 41.270 184.810 ;
        RECT 44.430 184.530 44.710 184.810 ;
        RECT 44.950 184.530 45.230 184.810 ;
        RECT 31.990 183.650 32.270 183.930 ;
        RECT 32.510 183.650 32.790 183.930 ;
        RECT 40.470 183.650 40.750 183.930 ;
        RECT 40.990 183.650 41.270 183.930 ;
        RECT 53.230 184.530 53.510 184.810 ;
        RECT 53.750 184.530 54.030 184.810 ;
        RECT 57.190 184.530 57.470 184.810 ;
        RECT 57.710 184.530 57.990 184.810 ;
        RECT 65.670 184.530 65.950 184.810 ;
        RECT 66.190 184.530 66.470 184.810 ;
        RECT 69.630 184.530 69.910 184.810 ;
        RECT 70.150 184.530 70.430 184.810 ;
        RECT 57.190 183.650 57.470 183.930 ;
        RECT 57.710 183.650 57.990 183.930 ;
        RECT 65.670 183.650 65.950 183.930 ;
        RECT 66.190 183.650 66.470 183.930 ;
        RECT 78.430 184.530 78.710 184.810 ;
        RECT 78.950 184.530 79.230 184.810 ;
        RECT 82.390 184.530 82.670 184.810 ;
        RECT 82.910 184.530 83.190 184.810 ;
        RECT 90.870 184.530 91.150 184.810 ;
        RECT 91.390 184.530 91.670 184.810 ;
        RECT 94.830 184.530 95.110 184.810 ;
        RECT 95.350 184.530 95.630 184.810 ;
        RECT 82.390 183.650 82.670 183.930 ;
        RECT 82.910 183.650 83.190 183.930 ;
        RECT 90.870 183.650 91.150 183.930 ;
        RECT 91.390 183.650 91.670 183.930 ;
        RECT 103.630 184.530 103.910 184.810 ;
        RECT 104.150 184.530 104.430 184.810 ;
        RECT 107.590 184.530 107.870 184.810 ;
        RECT 108.110 184.530 108.390 184.810 ;
        RECT 107.590 183.650 107.870 183.930 ;
        RECT 108.110 183.650 108.390 183.930 ;
        RECT 15.270 181.890 15.550 182.170 ;
        RECT 15.790 181.890 16.070 182.170 ;
        RECT 19.230 181.890 19.510 182.170 ;
        RECT 19.750 181.890 20.030 182.170 ;
        RECT 28.030 181.890 28.310 182.170 ;
        RECT 28.550 181.890 28.830 182.170 ;
        RECT 31.990 181.890 32.270 182.170 ;
        RECT 32.510 181.890 32.790 182.170 ;
        RECT 40.470 181.890 40.750 182.170 ;
        RECT 40.990 181.890 41.270 182.170 ;
        RECT 44.430 181.890 44.710 182.170 ;
        RECT 44.950 181.890 45.230 182.170 ;
        RECT 53.230 181.890 53.510 182.170 ;
        RECT 53.750 181.890 54.030 182.170 ;
        RECT 57.190 181.890 57.470 182.170 ;
        RECT 57.710 181.890 57.990 182.170 ;
        RECT 65.670 181.890 65.950 182.170 ;
        RECT 66.190 181.890 66.470 182.170 ;
        RECT 69.630 181.890 69.910 182.170 ;
        RECT 70.150 181.890 70.430 182.170 ;
        RECT 78.430 181.890 78.710 182.170 ;
        RECT 78.950 181.890 79.230 182.170 ;
        RECT 82.390 181.890 82.670 182.170 ;
        RECT 82.910 181.890 83.190 182.170 ;
        RECT 90.870 181.890 91.150 182.170 ;
        RECT 91.390 181.890 91.670 182.170 ;
        RECT 94.830 181.890 95.110 182.170 ;
        RECT 95.350 181.890 95.630 182.170 ;
        RECT 103.630 181.890 103.910 182.170 ;
        RECT 104.150 181.890 104.430 182.170 ;
        RECT 107.590 181.890 107.870 182.170 ;
        RECT 108.110 181.890 108.390 182.170 ;
        RECT 116.070 182.770 116.350 183.050 ;
        RECT 116.590 182.770 116.870 183.050 ;
        RECT 120.030 182.770 120.310 183.050 ;
        RECT 120.550 182.770 120.830 183.050 ;
        RECT 116.070 181.890 116.350 182.170 ;
        RECT 116.590 181.890 116.870 182.170 ;
        RECT 120.030 181.890 120.310 182.170 ;
        RECT 120.550 181.890 120.830 182.170 ;
        RECT 15.270 180.130 15.550 180.410 ;
        RECT 15.790 180.130 16.070 180.410 ;
        RECT 19.230 180.130 19.510 180.410 ;
        RECT 19.750 180.130 20.030 180.410 ;
        RECT 28.030 180.130 28.310 180.410 ;
        RECT 28.550 180.130 28.830 180.410 ;
        RECT 31.990 180.130 32.270 180.410 ;
        RECT 32.510 180.130 32.790 180.410 ;
        RECT 40.470 180.130 40.750 180.410 ;
        RECT 40.990 180.130 41.270 180.410 ;
        RECT 44.430 180.130 44.710 180.410 ;
        RECT 44.950 180.130 45.230 180.410 ;
        RECT 53.230 180.130 53.510 180.410 ;
        RECT 53.750 180.130 54.030 180.410 ;
        RECT 57.190 180.130 57.470 180.410 ;
        RECT 57.710 180.130 57.990 180.410 ;
        RECT 65.670 180.130 65.950 180.410 ;
        RECT 66.190 180.130 66.470 180.410 ;
        RECT 69.630 180.130 69.910 180.410 ;
        RECT 70.150 180.130 70.430 180.410 ;
        RECT 78.430 180.130 78.710 180.410 ;
        RECT 78.950 180.130 79.230 180.410 ;
        RECT 82.390 180.130 82.670 180.410 ;
        RECT 82.910 180.130 83.190 180.410 ;
        RECT 90.870 180.130 91.150 180.410 ;
        RECT 91.390 180.130 91.670 180.410 ;
        RECT 94.830 180.130 95.110 180.410 ;
        RECT 95.350 180.130 95.630 180.410 ;
        RECT 103.630 180.130 103.910 180.410 ;
        RECT 104.150 180.130 104.430 180.410 ;
        RECT 107.590 180.130 107.870 180.410 ;
        RECT 108.110 180.130 108.390 180.410 ;
        RECT 116.070 180.130 116.350 180.410 ;
        RECT 116.590 180.130 116.870 180.410 ;
        RECT 120.030 180.130 120.310 180.410 ;
        RECT 120.550 180.130 120.830 180.410 ;
        RECT 19.230 179.250 19.510 179.530 ;
        RECT 19.750 179.250 20.030 179.530 ;
        RECT 28.030 179.250 28.310 179.530 ;
        RECT 28.550 179.250 28.830 179.530 ;
        RECT 44.430 179.250 44.710 179.530 ;
        RECT 44.950 179.250 45.230 179.530 ;
        RECT 53.230 179.250 53.510 179.530 ;
        RECT 53.750 179.250 54.030 179.530 ;
        RECT 69.630 179.250 69.910 179.530 ;
        RECT 70.150 179.250 70.430 179.530 ;
        RECT 78.430 179.250 78.710 179.530 ;
        RECT 78.950 179.250 79.230 179.530 ;
        RECT 94.830 179.250 95.110 179.530 ;
        RECT 95.350 179.250 95.630 179.530 ;
        RECT 103.630 179.250 103.910 179.530 ;
        RECT 104.150 179.250 104.430 179.530 ;
        RECT 116.070 179.250 116.350 179.530 ;
        RECT 116.590 179.250 116.870 179.530 ;
        RECT 112.860 178.780 113.200 179.120 ;
        RECT 15.270 177.490 15.550 177.770 ;
        RECT 15.790 177.490 16.070 177.770 ;
        RECT 19.230 177.490 19.510 177.770 ;
        RECT 19.750 177.490 20.030 177.770 ;
        RECT 28.030 177.490 28.310 177.770 ;
        RECT 28.550 177.490 28.830 177.770 ;
        RECT 31.990 177.490 32.270 177.770 ;
        RECT 32.510 177.490 32.790 177.770 ;
        RECT 40.470 177.490 40.750 177.770 ;
        RECT 40.990 177.490 41.270 177.770 ;
        RECT 44.430 177.490 44.710 177.770 ;
        RECT 44.950 177.490 45.230 177.770 ;
        RECT 53.230 177.490 53.510 177.770 ;
        RECT 53.750 177.490 54.030 177.770 ;
        RECT 57.190 177.490 57.470 177.770 ;
        RECT 57.710 177.490 57.990 177.770 ;
        RECT 65.670 177.490 65.950 177.770 ;
        RECT 66.190 177.490 66.470 177.770 ;
        RECT 69.630 177.490 69.910 177.770 ;
        RECT 70.150 177.490 70.430 177.770 ;
        RECT 78.430 177.490 78.710 177.770 ;
        RECT 78.950 177.490 79.230 177.770 ;
        RECT 82.390 177.490 82.670 177.770 ;
        RECT 82.910 177.490 83.190 177.770 ;
        RECT 90.870 177.490 91.150 177.770 ;
        RECT 91.390 177.490 91.670 177.770 ;
        RECT 94.830 177.490 95.110 177.770 ;
        RECT 95.350 177.490 95.630 177.770 ;
        RECT 103.630 177.490 103.910 177.770 ;
        RECT 104.150 177.490 104.430 177.770 ;
        RECT 107.590 177.490 107.870 177.770 ;
        RECT 108.110 177.490 108.390 177.770 ;
        RECT 116.070 177.490 116.350 177.770 ;
        RECT 116.590 177.490 116.870 177.770 ;
        RECT 120.030 177.490 120.310 177.770 ;
        RECT 120.550 177.490 120.830 177.770 ;
        RECT 120.030 176.610 120.310 176.890 ;
        RECT 120.550 176.610 120.830 176.890 ;
        RECT 15.270 175.730 15.550 176.010 ;
        RECT 15.790 175.730 16.070 176.010 ;
        RECT 19.230 175.730 19.510 176.010 ;
        RECT 19.750 175.730 20.030 176.010 ;
        RECT 28.030 175.730 28.310 176.010 ;
        RECT 28.550 175.730 28.830 176.010 ;
        RECT 31.990 175.730 32.270 176.010 ;
        RECT 32.510 175.730 32.790 176.010 ;
        RECT 40.470 175.730 40.750 176.010 ;
        RECT 40.990 175.730 41.270 176.010 ;
        RECT 44.430 175.730 44.710 176.010 ;
        RECT 44.950 175.730 45.230 176.010 ;
        RECT 53.230 175.730 53.510 176.010 ;
        RECT 53.750 175.730 54.030 176.010 ;
        RECT 57.190 175.730 57.470 176.010 ;
        RECT 57.710 175.730 57.990 176.010 ;
        RECT 65.670 175.730 65.950 176.010 ;
        RECT 66.190 175.730 66.470 176.010 ;
        RECT 69.630 175.730 69.910 176.010 ;
        RECT 70.150 175.730 70.430 176.010 ;
        RECT 78.430 175.730 78.710 176.010 ;
        RECT 78.950 175.730 79.230 176.010 ;
        RECT 82.390 175.730 82.670 176.010 ;
        RECT 82.910 175.730 83.190 176.010 ;
        RECT 90.870 175.730 91.150 176.010 ;
        RECT 91.390 175.730 91.670 176.010 ;
        RECT 94.830 175.730 95.110 176.010 ;
        RECT 95.350 175.730 95.630 176.010 ;
        RECT 103.630 175.730 103.910 176.010 ;
        RECT 104.150 175.730 104.430 176.010 ;
        RECT 107.590 175.730 107.870 176.010 ;
        RECT 108.110 175.730 108.390 176.010 ;
        RECT 116.070 174.850 116.350 175.130 ;
        RECT 116.590 174.850 116.870 175.130 ;
        RECT 120.030 174.850 120.310 175.130 ;
        RECT 120.550 174.850 120.830 175.130 ;
        RECT 15.270 173.970 15.550 174.250 ;
        RECT 15.790 173.970 16.070 174.250 ;
        RECT 19.230 173.970 19.510 174.250 ;
        RECT 19.750 173.970 20.030 174.250 ;
        RECT 28.030 173.970 28.310 174.250 ;
        RECT 28.550 173.970 28.830 174.250 ;
        RECT 31.990 173.970 32.270 174.250 ;
        RECT 32.510 173.970 32.790 174.250 ;
        RECT 40.470 173.970 40.750 174.250 ;
        RECT 40.990 173.970 41.270 174.250 ;
        RECT 44.430 173.970 44.710 174.250 ;
        RECT 44.950 173.970 45.230 174.250 ;
        RECT 53.230 173.970 53.510 174.250 ;
        RECT 53.750 173.970 54.030 174.250 ;
        RECT 57.190 173.970 57.470 174.250 ;
        RECT 57.710 173.970 57.990 174.250 ;
        RECT 65.670 173.970 65.950 174.250 ;
        RECT 66.190 173.970 66.470 174.250 ;
        RECT 69.630 173.970 69.910 174.250 ;
        RECT 70.150 173.970 70.430 174.250 ;
        RECT 78.430 173.970 78.710 174.250 ;
        RECT 78.950 173.970 79.230 174.250 ;
        RECT 82.390 173.970 82.670 174.250 ;
        RECT 82.910 173.970 83.190 174.250 ;
        RECT 90.870 173.970 91.150 174.250 ;
        RECT 91.390 173.970 91.670 174.250 ;
        RECT 94.830 173.970 95.110 174.250 ;
        RECT 95.350 173.970 95.630 174.250 ;
        RECT 103.630 173.970 103.910 174.250 ;
        RECT 104.150 173.970 104.430 174.250 ;
        RECT 107.590 173.970 107.870 174.250 ;
        RECT 108.110 173.970 108.390 174.250 ;
        RECT 116.070 173.090 116.350 173.370 ;
        RECT 116.590 173.090 116.870 173.370 ;
        RECT 120.030 173.090 120.310 173.370 ;
        RECT 120.550 173.090 120.830 173.370 ;
        RECT 15.270 171.330 15.550 171.610 ;
        RECT 15.790 171.330 16.070 171.610 ;
        RECT 19.230 171.330 19.510 171.610 ;
        RECT 19.750 171.330 20.030 171.610 ;
        RECT 28.030 171.330 28.310 171.610 ;
        RECT 28.550 171.330 28.830 171.610 ;
        RECT 31.990 171.330 32.270 171.610 ;
        RECT 32.510 171.330 32.790 171.610 ;
        RECT 40.470 171.330 40.750 171.610 ;
        RECT 40.990 171.330 41.270 171.610 ;
        RECT 44.430 171.330 44.710 171.610 ;
        RECT 44.950 171.330 45.230 171.610 ;
        RECT 53.230 171.330 53.510 171.610 ;
        RECT 53.750 171.330 54.030 171.610 ;
        RECT 57.190 171.330 57.470 171.610 ;
        RECT 57.710 171.330 57.990 171.610 ;
        RECT 65.670 171.330 65.950 171.610 ;
        RECT 66.190 171.330 66.470 171.610 ;
        RECT 69.630 171.330 69.910 171.610 ;
        RECT 70.150 171.330 70.430 171.610 ;
        RECT 78.430 171.330 78.710 171.610 ;
        RECT 78.950 171.330 79.230 171.610 ;
        RECT 82.390 171.330 82.670 171.610 ;
        RECT 82.910 171.330 83.190 171.610 ;
        RECT 90.870 171.330 91.150 171.610 ;
        RECT 91.390 171.330 91.670 171.610 ;
        RECT 94.830 171.330 95.110 171.610 ;
        RECT 95.350 171.330 95.630 171.610 ;
        RECT 103.630 171.330 103.910 171.610 ;
        RECT 104.150 171.330 104.430 171.610 ;
        RECT 107.590 171.330 107.870 171.610 ;
        RECT 108.110 171.330 108.390 171.610 ;
        RECT 15.270 169.570 15.550 169.850 ;
        RECT 15.790 169.570 16.070 169.850 ;
        RECT 31.990 169.570 32.270 169.850 ;
        RECT 32.510 169.570 32.790 169.850 ;
        RECT 40.470 169.570 40.750 169.850 ;
        RECT 40.990 169.570 41.270 169.850 ;
        RECT 57.190 169.570 57.470 169.850 ;
        RECT 57.710 169.570 57.990 169.850 ;
        RECT 65.670 169.570 65.950 169.850 ;
        RECT 66.190 169.570 66.470 169.850 ;
        RECT 82.390 169.570 82.670 169.850 ;
        RECT 82.910 169.570 83.190 169.850 ;
        RECT 90.870 169.570 91.150 169.850 ;
        RECT 91.390 169.570 91.670 169.850 ;
        RECT 107.590 169.570 107.870 169.850 ;
        RECT 108.110 169.570 108.390 169.850 ;
        RECT 15.270 168.690 15.550 168.970 ;
        RECT 15.790 168.690 16.070 168.970 ;
        RECT 31.990 168.690 32.270 168.970 ;
        RECT 32.510 168.690 32.790 168.970 ;
        RECT 40.470 168.690 40.750 168.970 ;
        RECT 40.990 168.690 41.270 168.970 ;
        RECT 22.110 167.480 22.390 167.760 ;
        RECT 22.630 167.480 22.910 167.760 ;
        RECT 15.270 166.930 15.550 167.210 ;
        RECT 15.790 166.930 16.070 167.210 ;
        RECT 22.110 166.960 22.390 167.240 ;
        RECT 22.630 166.960 22.910 167.240 ;
        RECT 25.150 167.480 25.430 167.760 ;
        RECT 25.670 167.480 25.950 167.760 ;
        RECT 57.190 168.690 57.470 168.970 ;
        RECT 57.710 168.690 57.990 168.970 ;
        RECT 65.670 168.690 65.950 168.970 ;
        RECT 66.190 168.690 66.470 168.970 ;
        RECT 47.310 167.480 47.590 167.760 ;
        RECT 47.830 167.480 48.110 167.760 ;
        RECT 25.150 166.960 25.430 167.240 ;
        RECT 25.670 166.960 25.950 167.240 ;
        RECT 31.990 166.930 32.270 167.210 ;
        RECT 32.510 166.930 32.790 167.210 ;
        RECT 40.470 166.930 40.750 167.210 ;
        RECT 40.990 166.930 41.270 167.210 ;
        RECT 47.310 166.960 47.590 167.240 ;
        RECT 47.830 166.960 48.110 167.240 ;
        RECT 50.350 167.480 50.630 167.760 ;
        RECT 50.870 167.480 51.150 167.760 ;
        RECT 82.390 168.690 82.670 168.970 ;
        RECT 82.910 168.690 83.190 168.970 ;
        RECT 90.870 168.690 91.150 168.970 ;
        RECT 91.390 168.690 91.670 168.970 ;
        RECT 72.510 167.480 72.790 167.760 ;
        RECT 73.030 167.480 73.310 167.760 ;
        RECT 50.350 166.960 50.630 167.240 ;
        RECT 50.870 166.960 51.150 167.240 ;
        RECT 57.190 166.930 57.470 167.210 ;
        RECT 57.710 166.930 57.990 167.210 ;
        RECT 65.670 166.930 65.950 167.210 ;
        RECT 66.190 166.930 66.470 167.210 ;
        RECT 72.510 166.960 72.790 167.240 ;
        RECT 73.030 166.960 73.310 167.240 ;
        RECT 75.550 167.480 75.830 167.760 ;
        RECT 76.070 167.480 76.350 167.760 ;
        RECT 107.590 168.690 107.870 168.970 ;
        RECT 108.110 168.690 108.390 168.970 ;
        RECT 97.710 167.480 97.990 167.760 ;
        RECT 98.230 167.480 98.510 167.760 ;
        RECT 75.550 166.960 75.830 167.240 ;
        RECT 76.070 166.960 76.350 167.240 ;
        RECT 82.390 166.930 82.670 167.210 ;
        RECT 82.910 166.930 83.190 167.210 ;
        RECT 90.870 166.930 91.150 167.210 ;
        RECT 91.390 166.930 91.670 167.210 ;
        RECT 97.710 166.960 97.990 167.240 ;
        RECT 98.230 166.960 98.510 167.240 ;
        RECT 100.750 167.480 101.030 167.760 ;
        RECT 101.270 167.480 101.550 167.760 ;
        RECT 100.750 166.960 101.030 167.240 ;
        RECT 101.270 166.960 101.550 167.240 ;
        RECT 107.590 166.930 107.870 167.210 ;
        RECT 108.110 166.930 108.390 167.210 ;
        RECT 120.030 166.930 120.310 167.210 ;
        RECT 120.550 166.930 120.830 167.210 ;
        RECT 18.190 166.310 18.470 166.590 ;
        RECT 18.190 165.790 18.470 166.070 ;
        RECT 15.270 165.170 15.550 165.450 ;
        RECT 15.790 165.170 16.070 165.450 ;
        RECT 29.590 166.310 29.870 166.590 ;
        RECT 29.590 165.790 29.870 166.070 ;
        RECT 43.390 166.310 43.670 166.590 ;
        RECT 43.390 165.790 43.670 166.070 ;
        RECT 31.990 165.170 32.270 165.450 ;
        RECT 32.510 165.170 32.790 165.450 ;
        RECT 40.470 165.170 40.750 165.450 ;
        RECT 40.990 165.170 41.270 165.450 ;
        RECT 54.790 166.310 55.070 166.590 ;
        RECT 54.790 165.790 55.070 166.070 ;
        RECT 68.590 166.310 68.870 166.590 ;
        RECT 68.590 165.790 68.870 166.070 ;
        RECT 57.190 165.170 57.470 165.450 ;
        RECT 57.710 165.170 57.990 165.450 ;
        RECT 65.670 165.170 65.950 165.450 ;
        RECT 66.190 165.170 66.470 165.450 ;
        RECT 79.990 166.310 80.270 166.590 ;
        RECT 79.990 165.790 80.270 166.070 ;
        RECT 93.790 166.310 94.070 166.590 ;
        RECT 93.790 165.790 94.070 166.070 ;
        RECT 82.390 165.170 82.670 165.450 ;
        RECT 82.910 165.170 83.190 165.450 ;
        RECT 90.870 165.170 91.150 165.450 ;
        RECT 91.390 165.170 91.670 165.450 ;
        RECT 105.190 166.310 105.470 166.590 ;
        RECT 105.190 165.790 105.470 166.070 ;
        RECT 116.070 166.050 116.350 166.330 ;
        RECT 116.590 166.050 116.870 166.330 ;
        RECT 107.590 165.170 107.870 165.450 ;
        RECT 108.110 165.170 108.390 165.450 ;
        RECT 120.030 165.170 120.310 165.450 ;
        RECT 120.550 165.170 120.830 165.450 ;
        RECT 15.270 164.290 15.550 164.570 ;
        RECT 15.790 164.290 16.070 164.570 ;
        RECT 31.990 164.290 32.270 164.570 ;
        RECT 32.510 164.290 32.790 164.570 ;
        RECT 40.470 164.290 40.750 164.570 ;
        RECT 40.990 164.290 41.270 164.570 ;
        RECT 22.110 163.080 22.390 163.360 ;
        RECT 22.630 163.080 22.910 163.360 ;
        RECT 15.270 162.530 15.550 162.810 ;
        RECT 15.790 162.530 16.070 162.810 ;
        RECT 22.110 162.560 22.390 162.840 ;
        RECT 22.630 162.560 22.910 162.840 ;
        RECT 25.150 163.080 25.430 163.360 ;
        RECT 25.670 163.080 25.950 163.360 ;
        RECT 57.190 164.290 57.470 164.570 ;
        RECT 57.710 164.290 57.990 164.570 ;
        RECT 65.670 164.290 65.950 164.570 ;
        RECT 66.190 164.290 66.470 164.570 ;
        RECT 47.310 163.080 47.590 163.360 ;
        RECT 47.830 163.080 48.110 163.360 ;
        RECT 25.150 162.560 25.430 162.840 ;
        RECT 25.670 162.560 25.950 162.840 ;
        RECT 31.990 162.530 32.270 162.810 ;
        RECT 32.510 162.530 32.790 162.810 ;
        RECT 40.470 162.530 40.750 162.810 ;
        RECT 40.990 162.530 41.270 162.810 ;
        RECT 47.310 162.560 47.590 162.840 ;
        RECT 47.830 162.560 48.110 162.840 ;
        RECT 50.350 163.080 50.630 163.360 ;
        RECT 50.870 163.080 51.150 163.360 ;
        RECT 82.390 164.290 82.670 164.570 ;
        RECT 82.910 164.290 83.190 164.570 ;
        RECT 90.870 164.290 91.150 164.570 ;
        RECT 91.390 164.290 91.670 164.570 ;
        RECT 72.510 163.080 72.790 163.360 ;
        RECT 73.030 163.080 73.310 163.360 ;
        RECT 50.350 162.560 50.630 162.840 ;
        RECT 50.870 162.560 51.150 162.840 ;
        RECT 57.190 162.530 57.470 162.810 ;
        RECT 57.710 162.530 57.990 162.810 ;
        RECT 65.670 162.530 65.950 162.810 ;
        RECT 66.190 162.530 66.470 162.810 ;
        RECT 72.510 162.560 72.790 162.840 ;
        RECT 73.030 162.560 73.310 162.840 ;
        RECT 75.550 163.080 75.830 163.360 ;
        RECT 76.070 163.080 76.350 163.360 ;
        RECT 107.590 164.290 107.870 164.570 ;
        RECT 108.110 164.290 108.390 164.570 ;
        RECT 97.710 163.080 97.990 163.360 ;
        RECT 98.230 163.080 98.510 163.360 ;
        RECT 75.550 162.560 75.830 162.840 ;
        RECT 76.070 162.560 76.350 162.840 ;
        RECT 82.390 162.530 82.670 162.810 ;
        RECT 82.910 162.530 83.190 162.810 ;
        RECT 90.870 162.530 91.150 162.810 ;
        RECT 91.390 162.530 91.670 162.810 ;
        RECT 97.710 162.560 97.990 162.840 ;
        RECT 98.230 162.560 98.510 162.840 ;
        RECT 100.750 163.080 101.030 163.360 ;
        RECT 101.270 163.080 101.550 163.360 ;
        RECT 114.710 163.850 114.990 164.130 ;
        RECT 115.230 163.850 115.510 164.130 ;
        RECT 120.030 163.410 120.310 163.690 ;
        RECT 120.550 163.410 120.830 163.690 ;
        RECT 100.750 162.560 101.030 162.840 ;
        RECT 101.270 162.560 101.550 162.840 ;
        RECT 107.590 162.530 107.870 162.810 ;
        RECT 108.110 162.530 108.390 162.810 ;
        RECT 17.405 161.910 17.685 162.190 ;
        RECT 17.405 161.390 17.685 161.670 ;
        RECT 15.270 160.770 15.550 161.050 ;
        RECT 15.790 160.770 16.070 161.050 ;
        RECT 30.375 161.910 30.655 162.190 ;
        RECT 30.375 161.390 30.655 161.670 ;
        RECT 42.605 161.910 42.885 162.190 ;
        RECT 42.605 161.390 42.885 161.670 ;
        RECT 31.990 160.770 32.270 161.050 ;
        RECT 32.510 160.770 32.790 161.050 ;
        RECT 40.470 160.770 40.750 161.050 ;
        RECT 40.990 160.770 41.270 161.050 ;
        RECT 55.575 161.910 55.855 162.190 ;
        RECT 55.575 161.390 55.855 161.670 ;
        RECT 67.805 161.910 68.085 162.190 ;
        RECT 67.805 161.390 68.085 161.670 ;
        RECT 57.190 160.770 57.470 161.050 ;
        RECT 57.710 160.770 57.990 161.050 ;
        RECT 65.670 160.770 65.950 161.050 ;
        RECT 66.190 160.770 66.470 161.050 ;
        RECT 80.775 161.910 81.055 162.190 ;
        RECT 80.775 161.390 81.055 161.670 ;
        RECT 93.005 161.910 93.285 162.190 ;
        RECT 93.005 161.390 93.285 161.670 ;
        RECT 82.390 160.770 82.670 161.050 ;
        RECT 82.910 160.770 83.190 161.050 ;
        RECT 90.870 160.770 91.150 161.050 ;
        RECT 91.390 160.770 91.670 161.050 ;
        RECT 105.975 161.910 106.255 162.190 ;
        RECT 105.975 161.390 106.255 161.670 ;
        RECT 120.030 161.650 120.310 161.930 ;
        RECT 120.550 161.650 120.830 161.930 ;
        RECT 122.190 161.210 122.470 161.490 ;
        RECT 122.710 161.210 122.990 161.490 ;
        RECT 107.590 160.770 107.870 161.050 ;
        RECT 108.110 160.770 108.390 161.050 ;
        RECT 15.270 159.890 15.550 160.170 ;
        RECT 15.790 159.890 16.070 160.170 ;
        RECT 31.990 159.890 32.270 160.170 ;
        RECT 32.510 159.890 32.790 160.170 ;
        RECT 40.470 159.890 40.750 160.170 ;
        RECT 40.990 159.890 41.270 160.170 ;
        RECT 22.110 158.680 22.390 158.960 ;
        RECT 22.630 158.680 22.910 158.960 ;
        RECT 15.270 158.130 15.550 158.410 ;
        RECT 15.790 158.130 16.070 158.410 ;
        RECT 22.110 158.160 22.390 158.440 ;
        RECT 22.630 158.160 22.910 158.440 ;
        RECT 25.150 158.680 25.430 158.960 ;
        RECT 25.670 158.680 25.950 158.960 ;
        RECT 57.190 159.890 57.470 160.170 ;
        RECT 57.710 159.890 57.990 160.170 ;
        RECT 65.670 159.890 65.950 160.170 ;
        RECT 66.190 159.890 66.470 160.170 ;
        RECT 47.310 158.680 47.590 158.960 ;
        RECT 47.830 158.680 48.110 158.960 ;
        RECT 25.150 158.160 25.430 158.440 ;
        RECT 25.670 158.160 25.950 158.440 ;
        RECT 31.990 158.130 32.270 158.410 ;
        RECT 32.510 158.130 32.790 158.410 ;
        RECT 40.470 158.130 40.750 158.410 ;
        RECT 40.990 158.130 41.270 158.410 ;
        RECT 47.310 158.160 47.590 158.440 ;
        RECT 47.830 158.160 48.110 158.440 ;
        RECT 50.350 158.680 50.630 158.960 ;
        RECT 50.870 158.680 51.150 158.960 ;
        RECT 82.390 159.890 82.670 160.170 ;
        RECT 82.910 159.890 83.190 160.170 ;
        RECT 90.870 159.890 91.150 160.170 ;
        RECT 91.390 159.890 91.670 160.170 ;
        RECT 72.510 158.680 72.790 158.960 ;
        RECT 73.030 158.680 73.310 158.960 ;
        RECT 50.350 158.160 50.630 158.440 ;
        RECT 50.870 158.160 51.150 158.440 ;
        RECT 57.190 158.130 57.470 158.410 ;
        RECT 57.710 158.130 57.990 158.410 ;
        RECT 65.670 158.130 65.950 158.410 ;
        RECT 66.190 158.130 66.470 158.410 ;
        RECT 72.510 158.160 72.790 158.440 ;
        RECT 73.030 158.160 73.310 158.440 ;
        RECT 75.550 158.680 75.830 158.960 ;
        RECT 76.070 158.680 76.350 158.960 ;
        RECT 107.590 159.890 107.870 160.170 ;
        RECT 108.110 159.890 108.390 160.170 ;
        RECT 120.030 159.890 120.310 160.170 ;
        RECT 120.550 159.890 120.830 160.170 ;
        RECT 97.710 158.680 97.990 158.960 ;
        RECT 98.230 158.680 98.510 158.960 ;
        RECT 75.550 158.160 75.830 158.440 ;
        RECT 76.070 158.160 76.350 158.440 ;
        RECT 82.390 158.130 82.670 158.410 ;
        RECT 82.910 158.130 83.190 158.410 ;
        RECT 90.870 158.130 91.150 158.410 ;
        RECT 91.390 158.130 91.670 158.410 ;
        RECT 97.710 158.160 97.990 158.440 ;
        RECT 98.230 158.160 98.510 158.440 ;
        RECT 100.750 158.680 101.030 158.960 ;
        RECT 101.270 158.680 101.550 158.960 ;
        RECT 116.070 159.010 116.350 159.290 ;
        RECT 116.590 159.010 116.870 159.290 ;
        RECT 100.750 158.160 101.030 158.440 ;
        RECT 101.270 158.160 101.550 158.440 ;
        RECT 107.590 158.130 107.870 158.410 ;
        RECT 108.110 158.130 108.390 158.410 ;
        RECT 116.070 158.130 116.350 158.410 ;
        RECT 116.590 158.130 116.870 158.410 ;
        RECT 120.030 158.130 120.310 158.410 ;
        RECT 120.550 158.130 120.830 158.410 ;
        RECT 16.690 157.510 16.970 157.790 ;
        RECT 13.270 156.810 13.550 157.090 ;
        RECT 13.790 156.810 14.070 157.090 ;
        RECT 16.690 156.990 16.970 157.270 ;
        RECT 15.270 156.370 15.550 156.650 ;
        RECT 15.790 156.370 16.070 156.650 ;
        RECT 31.090 157.510 31.370 157.790 ;
        RECT 31.090 156.990 31.370 157.270 ;
        RECT 41.890 157.510 42.170 157.790 ;
        RECT 33.990 156.810 34.270 157.090 ;
        RECT 34.510 156.810 34.790 157.090 ;
        RECT 38.470 156.810 38.750 157.090 ;
        RECT 38.990 156.810 39.270 157.090 ;
        RECT 41.890 156.990 42.170 157.270 ;
        RECT 31.990 156.370 32.270 156.650 ;
        RECT 32.510 156.370 32.790 156.650 ;
        RECT 40.470 156.370 40.750 156.650 ;
        RECT 40.990 156.370 41.270 156.650 ;
        RECT 56.290 157.510 56.570 157.790 ;
        RECT 56.290 156.990 56.570 157.270 ;
        RECT 67.090 157.510 67.370 157.790 ;
        RECT 59.190 156.810 59.470 157.090 ;
        RECT 59.710 156.810 59.990 157.090 ;
        RECT 63.670 156.810 63.950 157.090 ;
        RECT 64.190 156.810 64.470 157.090 ;
        RECT 67.090 156.990 67.370 157.270 ;
        RECT 57.190 156.370 57.470 156.650 ;
        RECT 57.710 156.370 57.990 156.650 ;
        RECT 65.670 156.370 65.950 156.650 ;
        RECT 66.190 156.370 66.470 156.650 ;
        RECT 81.490 157.510 81.770 157.790 ;
        RECT 81.490 156.990 81.770 157.270 ;
        RECT 92.290 157.510 92.570 157.790 ;
        RECT 84.390 156.810 84.670 157.090 ;
        RECT 84.910 156.810 85.190 157.090 ;
        RECT 88.870 156.810 89.150 157.090 ;
        RECT 89.390 156.810 89.670 157.090 ;
        RECT 92.290 156.990 92.570 157.270 ;
        RECT 82.390 156.370 82.670 156.650 ;
        RECT 82.910 156.370 83.190 156.650 ;
        RECT 90.870 156.370 91.150 156.650 ;
        RECT 91.390 156.370 91.670 156.650 ;
        RECT 106.690 157.510 106.970 157.790 ;
        RECT 106.690 156.990 106.970 157.270 ;
        RECT 109.590 156.810 109.870 157.090 ;
        RECT 110.110 156.810 110.390 157.090 ;
        RECT 107.590 156.370 107.870 156.650 ;
        RECT 108.110 156.370 108.390 156.650 ;
        RECT 116.070 156.370 116.350 156.650 ;
        RECT 116.590 156.370 116.870 156.650 ;
        RECT 120.030 156.370 120.310 156.650 ;
        RECT 120.550 156.370 120.830 156.650 ;
        RECT 15.270 155.490 15.550 155.770 ;
        RECT 15.790 155.490 16.070 155.770 ;
        RECT 31.990 155.490 32.270 155.770 ;
        RECT 32.510 155.490 32.790 155.770 ;
        RECT 40.470 155.490 40.750 155.770 ;
        RECT 40.990 155.490 41.270 155.770 ;
        RECT 22.110 154.280 22.390 154.560 ;
        RECT 22.630 154.280 22.910 154.560 ;
        RECT 15.270 153.730 15.550 154.010 ;
        RECT 15.790 153.730 16.070 154.010 ;
        RECT 22.110 153.760 22.390 154.040 ;
        RECT 22.630 153.760 22.910 154.040 ;
        RECT 25.150 154.280 25.430 154.560 ;
        RECT 25.670 154.280 25.950 154.560 ;
        RECT 57.190 155.490 57.470 155.770 ;
        RECT 57.710 155.490 57.990 155.770 ;
        RECT 65.670 155.490 65.950 155.770 ;
        RECT 66.190 155.490 66.470 155.770 ;
        RECT 47.310 154.280 47.590 154.560 ;
        RECT 47.830 154.280 48.110 154.560 ;
        RECT 25.150 153.760 25.430 154.040 ;
        RECT 25.670 153.760 25.950 154.040 ;
        RECT 31.990 153.730 32.270 154.010 ;
        RECT 32.510 153.730 32.790 154.010 ;
        RECT 40.470 153.730 40.750 154.010 ;
        RECT 40.990 153.730 41.270 154.010 ;
        RECT 47.310 153.760 47.590 154.040 ;
        RECT 47.830 153.760 48.110 154.040 ;
        RECT 50.350 154.280 50.630 154.560 ;
        RECT 50.870 154.280 51.150 154.560 ;
        RECT 82.390 155.490 82.670 155.770 ;
        RECT 82.910 155.490 83.190 155.770 ;
        RECT 90.870 155.490 91.150 155.770 ;
        RECT 91.390 155.490 91.670 155.770 ;
        RECT 72.510 154.280 72.790 154.560 ;
        RECT 73.030 154.280 73.310 154.560 ;
        RECT 50.350 153.760 50.630 154.040 ;
        RECT 50.870 153.760 51.150 154.040 ;
        RECT 57.190 153.730 57.470 154.010 ;
        RECT 57.710 153.730 57.990 154.010 ;
        RECT 65.670 153.730 65.950 154.010 ;
        RECT 66.190 153.730 66.470 154.010 ;
        RECT 72.510 153.760 72.790 154.040 ;
        RECT 73.030 153.760 73.310 154.040 ;
        RECT 75.550 154.280 75.830 154.560 ;
        RECT 76.070 154.280 76.350 154.560 ;
        RECT 107.590 155.490 107.870 155.770 ;
        RECT 108.110 155.490 108.390 155.770 ;
        RECT 97.710 154.280 97.990 154.560 ;
        RECT 98.230 154.280 98.510 154.560 ;
        RECT 75.550 153.760 75.830 154.040 ;
        RECT 76.070 153.760 76.350 154.040 ;
        RECT 82.390 153.730 82.670 154.010 ;
        RECT 82.910 153.730 83.190 154.010 ;
        RECT 90.870 153.730 91.150 154.010 ;
        RECT 91.390 153.730 91.670 154.010 ;
        RECT 97.710 153.760 97.990 154.040 ;
        RECT 98.230 153.760 98.510 154.040 ;
        RECT 100.750 154.280 101.030 154.560 ;
        RECT 101.270 154.280 101.550 154.560 ;
        RECT 100.750 153.760 101.030 154.040 ;
        RECT 101.270 153.760 101.550 154.040 ;
        RECT 107.590 153.730 107.870 154.010 ;
        RECT 108.110 153.730 108.390 154.010 ;
        RECT 15.270 151.970 15.550 152.250 ;
        RECT 15.790 151.970 16.070 152.250 ;
        RECT 31.990 151.970 32.270 152.250 ;
        RECT 32.510 151.970 32.790 152.250 ;
        RECT 40.470 151.970 40.750 152.250 ;
        RECT 40.990 151.970 41.270 152.250 ;
        RECT 57.190 151.970 57.470 152.250 ;
        RECT 57.710 151.970 57.990 152.250 ;
        RECT 65.670 151.970 65.950 152.250 ;
        RECT 66.190 151.970 66.470 152.250 ;
        RECT 82.390 151.970 82.670 152.250 ;
        RECT 82.910 151.970 83.190 152.250 ;
        RECT 90.870 151.970 91.150 152.250 ;
        RECT 91.390 151.970 91.670 152.250 ;
        RECT 107.590 151.970 107.870 152.250 ;
        RECT 108.110 151.970 108.390 152.250 ;
        RECT 102.550 150.620 102.890 150.960 ;
        RECT 116.070 154.610 116.350 154.890 ;
        RECT 116.590 154.610 116.870 154.890 ;
        RECT 120.030 154.610 120.310 154.890 ;
        RECT 120.550 154.610 120.830 154.890 ;
        RECT 116.070 153.730 116.350 154.010 ;
        RECT 116.590 153.730 116.870 154.010 ;
        RECT 120.030 153.730 120.310 154.010 ;
        RECT 120.550 153.730 120.830 154.010 ;
        RECT 116.070 151.970 116.350 152.250 ;
        RECT 116.590 151.970 116.870 152.250 ;
        RECT 120.030 151.970 120.310 152.250 ;
        RECT 120.550 151.970 120.830 152.250 ;
        RECT 15.270 148.450 15.550 148.730 ;
        RECT 15.790 148.450 16.070 148.730 ;
        RECT 19.230 148.450 19.510 148.730 ;
        RECT 19.750 148.450 20.030 148.730 ;
        RECT 28.030 148.450 28.310 148.730 ;
        RECT 28.550 148.450 28.830 148.730 ;
        RECT 31.990 148.450 32.270 148.730 ;
        RECT 32.510 148.450 32.790 148.730 ;
        RECT 40.470 148.450 40.750 148.730 ;
        RECT 40.990 148.450 41.270 148.730 ;
        RECT 44.430 148.450 44.710 148.730 ;
        RECT 44.950 148.450 45.230 148.730 ;
        RECT 53.230 148.450 53.510 148.730 ;
        RECT 53.750 148.450 54.030 148.730 ;
        RECT 57.190 148.450 57.470 148.730 ;
        RECT 57.710 148.450 57.990 148.730 ;
        RECT 65.670 148.450 65.950 148.730 ;
        RECT 66.190 148.450 66.470 148.730 ;
        RECT 69.630 148.450 69.910 148.730 ;
        RECT 70.150 148.450 70.430 148.730 ;
        RECT 78.430 148.450 78.710 148.730 ;
        RECT 78.950 148.450 79.230 148.730 ;
        RECT 82.390 148.450 82.670 148.730 ;
        RECT 82.910 148.450 83.190 148.730 ;
        RECT 90.870 148.450 91.150 148.730 ;
        RECT 91.390 148.450 91.670 148.730 ;
        RECT 94.830 148.450 95.110 148.730 ;
        RECT 95.350 148.450 95.630 148.730 ;
        RECT 103.630 148.450 103.910 148.730 ;
        RECT 104.150 148.450 104.430 148.730 ;
        RECT 107.590 148.450 107.870 148.730 ;
        RECT 108.110 148.450 108.390 148.730 ;
        RECT 116.070 150.210 116.350 150.490 ;
        RECT 116.590 150.210 116.870 150.490 ;
        RECT 120.030 150.210 120.310 150.490 ;
        RECT 120.550 150.210 120.830 150.490 ;
        RECT 120.030 149.330 120.310 149.610 ;
        RECT 120.550 149.330 120.830 149.610 ;
        RECT 120.030 147.570 120.310 147.850 ;
        RECT 120.550 147.570 120.830 147.850 ;
        RECT 120.030 145.810 120.310 146.090 ;
        RECT 120.550 145.810 120.830 146.090 ;
        RECT 122.190 145.370 122.470 145.650 ;
        RECT 122.710 145.370 122.990 145.650 ;
        RECT 15.270 144.930 15.550 145.210 ;
        RECT 15.790 144.930 16.070 145.210 ;
        RECT 19.230 144.930 19.510 145.210 ;
        RECT 19.750 144.930 20.030 145.210 ;
        RECT 28.030 144.930 28.310 145.210 ;
        RECT 28.550 144.930 28.830 145.210 ;
        RECT 31.990 144.930 32.270 145.210 ;
        RECT 32.510 144.930 32.790 145.210 ;
        RECT 40.470 144.930 40.750 145.210 ;
        RECT 40.990 144.930 41.270 145.210 ;
        RECT 44.430 144.930 44.710 145.210 ;
        RECT 44.950 144.930 45.230 145.210 ;
        RECT 53.230 144.930 53.510 145.210 ;
        RECT 53.750 144.930 54.030 145.210 ;
        RECT 57.190 144.930 57.470 145.210 ;
        RECT 57.710 144.930 57.990 145.210 ;
        RECT 65.670 144.930 65.950 145.210 ;
        RECT 66.190 144.930 66.470 145.210 ;
        RECT 69.630 144.930 69.910 145.210 ;
        RECT 70.150 144.930 70.430 145.210 ;
        RECT 78.430 144.930 78.710 145.210 ;
        RECT 78.950 144.930 79.230 145.210 ;
        RECT 82.390 144.930 82.670 145.210 ;
        RECT 82.910 144.930 83.190 145.210 ;
        RECT 90.870 144.930 91.150 145.210 ;
        RECT 91.390 144.930 91.670 145.210 ;
        RECT 94.830 144.930 95.110 145.210 ;
        RECT 95.350 144.930 95.630 145.210 ;
        RECT 103.630 144.930 103.910 145.210 ;
        RECT 104.150 144.930 104.430 145.210 ;
        RECT 107.590 144.930 107.870 145.210 ;
        RECT 108.110 144.930 108.390 145.210 ;
        RECT 120.030 144.050 120.310 144.330 ;
        RECT 120.550 144.050 120.830 144.330 ;
        RECT 15.270 143.170 15.550 143.450 ;
        RECT 15.790 143.170 16.070 143.450 ;
        RECT 19.230 143.170 19.510 143.450 ;
        RECT 19.750 143.170 20.030 143.450 ;
        RECT 28.030 143.170 28.310 143.450 ;
        RECT 28.550 143.170 28.830 143.450 ;
        RECT 31.990 143.170 32.270 143.450 ;
        RECT 32.510 143.170 32.790 143.450 ;
        RECT 40.470 143.170 40.750 143.450 ;
        RECT 40.990 143.170 41.270 143.450 ;
        RECT 44.430 143.170 44.710 143.450 ;
        RECT 44.950 143.170 45.230 143.450 ;
        RECT 53.230 143.170 53.510 143.450 ;
        RECT 53.750 143.170 54.030 143.450 ;
        RECT 57.190 143.170 57.470 143.450 ;
        RECT 57.710 143.170 57.990 143.450 ;
        RECT 65.670 143.170 65.950 143.450 ;
        RECT 66.190 143.170 66.470 143.450 ;
        RECT 69.630 143.170 69.910 143.450 ;
        RECT 70.150 143.170 70.430 143.450 ;
        RECT 78.430 143.170 78.710 143.450 ;
        RECT 78.950 143.170 79.230 143.450 ;
        RECT 82.390 143.170 82.670 143.450 ;
        RECT 82.910 143.170 83.190 143.450 ;
        RECT 90.870 143.170 91.150 143.450 ;
        RECT 91.390 143.170 91.670 143.450 ;
        RECT 94.830 143.170 95.110 143.450 ;
        RECT 95.350 143.170 95.630 143.450 ;
        RECT 103.630 143.170 103.910 143.450 ;
        RECT 104.150 143.170 104.430 143.450 ;
        RECT 107.590 143.170 107.870 143.450 ;
        RECT 108.110 143.170 108.390 143.450 ;
        RECT 116.070 143.170 116.350 143.450 ;
        RECT 116.590 143.170 116.870 143.450 ;
        RECT 19.230 142.290 19.510 142.570 ;
        RECT 19.750 142.290 20.030 142.570 ;
        RECT 28.030 142.290 28.310 142.570 ;
        RECT 28.550 142.290 28.830 142.570 ;
        RECT 44.430 142.290 44.710 142.570 ;
        RECT 44.950 142.290 45.230 142.570 ;
        RECT 53.230 142.290 53.510 142.570 ;
        RECT 53.750 142.290 54.030 142.570 ;
        RECT 69.630 142.290 69.910 142.570 ;
        RECT 70.150 142.290 70.430 142.570 ;
        RECT 78.430 142.290 78.710 142.570 ;
        RECT 78.950 142.290 79.230 142.570 ;
        RECT 94.830 142.290 95.110 142.570 ;
        RECT 95.350 142.290 95.630 142.570 ;
        RECT 103.630 142.290 103.910 142.570 ;
        RECT 104.150 142.290 104.430 142.570 ;
        RECT 15.270 141.410 15.550 141.690 ;
        RECT 15.790 141.410 16.070 141.690 ;
        RECT 31.990 141.410 32.270 141.690 ;
        RECT 32.510 141.410 32.790 141.690 ;
        RECT 40.470 141.410 40.750 141.690 ;
        RECT 40.990 141.410 41.270 141.690 ;
        RECT 57.190 141.410 57.470 141.690 ;
        RECT 57.710 141.410 57.990 141.690 ;
        RECT 65.670 141.410 65.950 141.690 ;
        RECT 66.190 141.410 66.470 141.690 ;
        RECT 82.390 141.410 82.670 141.690 ;
        RECT 82.910 141.410 83.190 141.690 ;
        RECT 90.870 141.410 91.150 141.690 ;
        RECT 91.390 141.410 91.670 141.690 ;
        RECT 107.590 141.410 107.870 141.690 ;
        RECT 108.110 141.410 108.390 141.690 ;
        RECT 113.910 140.970 114.190 141.250 ;
        RECT 114.430 140.970 114.710 141.250 ;
        RECT 15.270 140.530 15.550 140.810 ;
        RECT 15.790 140.530 16.070 140.810 ;
        RECT 31.990 140.530 32.270 140.810 ;
        RECT 32.510 140.530 32.790 140.810 ;
        RECT 40.470 140.530 40.750 140.810 ;
        RECT 40.990 140.530 41.270 140.810 ;
        RECT 57.190 140.530 57.470 140.810 ;
        RECT 57.710 140.530 57.990 140.810 ;
        RECT 65.670 140.530 65.950 140.810 ;
        RECT 66.190 140.530 66.470 140.810 ;
        RECT 82.390 140.530 82.670 140.810 ;
        RECT 82.910 140.530 83.190 140.810 ;
        RECT 90.870 140.530 91.150 140.810 ;
        RECT 91.390 140.530 91.670 140.810 ;
        RECT 107.590 140.530 107.870 140.810 ;
        RECT 108.110 140.530 108.390 140.810 ;
        RECT 15.270 137.890 15.550 138.170 ;
        RECT 15.790 137.890 16.070 138.170 ;
        RECT 31.990 137.890 32.270 138.170 ;
        RECT 32.510 137.890 32.790 138.170 ;
        RECT 19.230 137.010 19.510 137.290 ;
        RECT 19.750 137.010 20.030 137.290 ;
        RECT 28.030 137.010 28.310 137.290 ;
        RECT 28.550 137.010 28.830 137.290 ;
        RECT 40.470 137.890 40.750 138.170 ;
        RECT 40.990 137.890 41.270 138.170 ;
        RECT 57.190 137.890 57.470 138.170 ;
        RECT 57.710 137.890 57.990 138.170 ;
        RECT 44.430 137.010 44.710 137.290 ;
        RECT 44.950 137.010 45.230 137.290 ;
        RECT 53.230 137.010 53.510 137.290 ;
        RECT 53.750 137.010 54.030 137.290 ;
        RECT 65.670 137.890 65.950 138.170 ;
        RECT 66.190 137.890 66.470 138.170 ;
        RECT 82.390 137.890 82.670 138.170 ;
        RECT 82.910 137.890 83.190 138.170 ;
        RECT 69.630 137.010 69.910 137.290 ;
        RECT 70.150 137.010 70.430 137.290 ;
        RECT 78.430 137.010 78.710 137.290 ;
        RECT 78.950 137.010 79.230 137.290 ;
        RECT 90.870 137.890 91.150 138.170 ;
        RECT 91.390 137.890 91.670 138.170 ;
        RECT 107.590 137.890 107.870 138.170 ;
        RECT 108.110 137.890 108.390 138.170 ;
        RECT 94.830 137.010 95.110 137.290 ;
        RECT 95.350 137.010 95.630 137.290 ;
        RECT 103.630 137.010 103.910 137.290 ;
        RECT 104.150 137.010 104.430 137.290 ;
        RECT 120.030 137.010 120.310 137.290 ;
        RECT 120.550 137.010 120.830 137.290 ;
        RECT 116.070 136.130 116.350 136.410 ;
        RECT 116.590 136.130 116.870 136.410 ;
        RECT 15.270 135.250 15.550 135.530 ;
        RECT 15.790 135.250 16.070 135.530 ;
        RECT 19.230 135.250 19.510 135.530 ;
        RECT 19.750 135.250 20.030 135.530 ;
        RECT 28.030 135.250 28.310 135.530 ;
        RECT 28.550 135.250 28.830 135.530 ;
        RECT 31.990 135.250 32.270 135.530 ;
        RECT 32.510 135.250 32.790 135.530 ;
        RECT 40.470 135.250 40.750 135.530 ;
        RECT 40.990 135.250 41.270 135.530 ;
        RECT 44.430 135.250 44.710 135.530 ;
        RECT 44.950 135.250 45.230 135.530 ;
        RECT 53.230 135.250 53.510 135.530 ;
        RECT 53.750 135.250 54.030 135.530 ;
        RECT 57.190 135.250 57.470 135.530 ;
        RECT 57.710 135.250 57.990 135.530 ;
        RECT 65.670 135.250 65.950 135.530 ;
        RECT 66.190 135.250 66.470 135.530 ;
        RECT 69.630 135.250 69.910 135.530 ;
        RECT 70.150 135.250 70.430 135.530 ;
        RECT 78.430 135.250 78.710 135.530 ;
        RECT 78.950 135.250 79.230 135.530 ;
        RECT 82.390 135.250 82.670 135.530 ;
        RECT 82.910 135.250 83.190 135.530 ;
        RECT 90.870 135.250 91.150 135.530 ;
        RECT 91.390 135.250 91.670 135.530 ;
        RECT 94.830 135.250 95.110 135.530 ;
        RECT 95.350 135.250 95.630 135.530 ;
        RECT 103.630 135.250 103.910 135.530 ;
        RECT 104.150 135.250 104.430 135.530 ;
        RECT 107.590 135.250 107.870 135.530 ;
        RECT 108.110 135.250 108.390 135.530 ;
        RECT 116.070 135.250 116.350 135.530 ;
        RECT 116.590 135.250 116.870 135.530 ;
        RECT 120.030 135.250 120.310 135.530 ;
        RECT 120.550 135.250 120.830 135.530 ;
        RECT 15.270 134.370 15.550 134.650 ;
        RECT 15.790 134.370 16.070 134.650 ;
        RECT 19.230 134.370 19.510 134.650 ;
        RECT 19.750 134.370 20.030 134.650 ;
        RECT 28.030 134.370 28.310 134.650 ;
        RECT 28.550 134.370 28.830 134.650 ;
        RECT 31.990 134.370 32.270 134.650 ;
        RECT 32.510 134.370 32.790 134.650 ;
        RECT 40.470 134.370 40.750 134.650 ;
        RECT 40.990 134.370 41.270 134.650 ;
        RECT 44.430 134.370 44.710 134.650 ;
        RECT 44.950 134.370 45.230 134.650 ;
        RECT 53.230 134.370 53.510 134.650 ;
        RECT 53.750 134.370 54.030 134.650 ;
        RECT 57.190 134.370 57.470 134.650 ;
        RECT 57.710 134.370 57.990 134.650 ;
        RECT 65.670 134.370 65.950 134.650 ;
        RECT 66.190 134.370 66.470 134.650 ;
        RECT 69.630 134.370 69.910 134.650 ;
        RECT 70.150 134.370 70.430 134.650 ;
        RECT 78.430 134.370 78.710 134.650 ;
        RECT 78.950 134.370 79.230 134.650 ;
        RECT 82.390 134.370 82.670 134.650 ;
        RECT 82.910 134.370 83.190 134.650 ;
        RECT 90.870 134.370 91.150 134.650 ;
        RECT 91.390 134.370 91.670 134.650 ;
        RECT 94.830 134.370 95.110 134.650 ;
        RECT 95.350 134.370 95.630 134.650 ;
        RECT 103.630 134.370 103.910 134.650 ;
        RECT 104.150 134.370 104.430 134.650 ;
        RECT 107.590 134.370 107.870 134.650 ;
        RECT 108.110 134.370 108.390 134.650 ;
        RECT 116.070 134.370 116.350 134.650 ;
        RECT 116.590 134.370 116.870 134.650 ;
        RECT 120.030 134.370 120.310 134.650 ;
        RECT 120.550 134.370 120.830 134.650 ;
        RECT 93.790 130.640 94.070 130.920 ;
        RECT 93.790 130.120 94.070 130.400 ;
        RECT 79.990 129.710 80.270 129.990 ;
        RECT 79.990 129.190 80.270 129.470 ;
        RECT 68.590 128.780 68.870 129.060 ;
        RECT 68.590 128.260 68.870 128.540 ;
        RECT 54.790 127.850 55.070 128.130 ;
        RECT 54.790 127.330 55.070 127.610 ;
        RECT 43.390 126.920 43.670 127.200 ;
        RECT 43.390 126.400 43.670 126.680 ;
        RECT 29.590 125.990 29.870 126.270 ;
        RECT 29.590 125.470 29.870 125.750 ;
        RECT 18.190 125.060 18.470 125.340 ;
        RECT 18.190 124.540 18.470 124.820 ;
        RECT 42.605 124.130 42.885 124.410 ;
        RECT 42.605 123.610 42.885 123.890 ;
        RECT 30.370 123.200 30.650 123.480 ;
        RECT 30.370 122.680 30.650 122.960 ;
        RECT 17.405 122.270 17.685 122.550 ;
        RECT 17.405 121.750 17.685 122.030 ;
        RECT 92.290 121.340 92.570 121.620 ;
        RECT 92.290 120.820 92.570 121.100 ;
        RECT 81.485 120.410 81.765 120.690 ;
        RECT 81.485 119.890 81.765 120.170 ;
        RECT 67.090 119.480 67.370 119.760 ;
        RECT 67.090 118.960 67.370 119.240 ;
        RECT 56.285 118.550 56.565 118.830 ;
        RECT 56.285 118.030 56.565 118.310 ;
        RECT 41.890 117.620 42.170 117.900 ;
        RECT 41.890 117.100 42.170 117.380 ;
        RECT 31.085 116.690 31.365 116.970 ;
        RECT 31.085 116.170 31.365 116.450 ;
        RECT 16.690 115.760 16.970 116.040 ;
        RECT 16.690 115.240 16.970 115.520 ;
        RECT 38.440 114.830 38.720 115.110 ;
        RECT 38.440 114.310 38.720 114.590 ;
        RECT 33.960 113.900 34.240 114.180 ;
        RECT 33.960 113.380 34.240 113.660 ;
        RECT 13.240 112.970 13.520 113.250 ;
        RECT 13.240 112.450 13.520 112.730 ;
        RECT 113.880 113.100 114.160 113.380 ;
        RECT 113.880 112.580 114.160 112.860 ;
        RECT 115.260 113.100 115.540 113.380 ;
        RECT 115.260 112.580 115.540 112.860 ;
        RECT 55.200 110.850 55.480 111.130 ;
        RECT 55.720 110.850 56.000 111.130 ;
        RECT 113.910 110.850 114.190 111.130 ;
        RECT 114.430 110.850 114.710 111.130 ;
        RECT 55.170 107.090 55.450 107.370 ;
        RECT 55.170 106.570 55.450 106.850 ;
        RECT 80.840 108.990 81.120 109.270 ;
        RECT 81.360 108.990 81.640 109.270 ;
        RECT 115.290 108.990 115.570 109.270 ;
        RECT 115.810 108.990 116.090 109.270 ;
        RECT 80.810 107.090 81.090 107.370 ;
        RECT 80.810 106.570 81.090 106.850 ;
        RECT 22.830 105.510 23.110 105.790 ;
        RECT 22.830 104.990 23.110 105.270 ;
        RECT 113.150 105.510 113.430 105.790 ;
        RECT 113.150 104.990 113.430 105.270 ;
        RECT 21.510 102.490 21.790 102.770 ;
        RECT 21.510 101.970 21.790 102.250 ;
        RECT 25.470 102.490 25.750 102.770 ;
        RECT 25.470 101.970 25.750 102.250 ;
        RECT 42.630 102.490 42.910 102.770 ;
        RECT 42.630 101.970 42.910 102.250 ;
        RECT 46.590 102.490 46.870 102.770 ;
        RECT 46.590 101.970 46.870 102.250 ;
        RECT 89.390 102.490 89.670 102.770 ;
        RECT 89.390 101.970 89.670 102.250 ;
        RECT 93.350 102.490 93.630 102.770 ;
        RECT 93.350 101.970 93.630 102.250 ;
        RECT 110.510 102.490 110.790 102.770 ;
        RECT 110.510 101.970 110.790 102.250 ;
        RECT 114.470 102.490 114.750 102.770 ;
        RECT 114.470 101.970 114.750 102.250 ;
        RECT 18.870 99.470 19.150 99.750 ;
        RECT 18.870 98.950 19.150 99.230 ;
        RECT 20.190 99.470 20.470 99.750 ;
        RECT 20.190 98.950 20.470 99.230 ;
        RECT 26.790 99.470 27.070 99.750 ;
        RECT 26.790 98.950 27.070 99.230 ;
        RECT 28.110 99.470 28.390 99.750 ;
        RECT 28.110 98.950 28.390 99.230 ;
        RECT 39.990 99.470 40.270 99.750 ;
        RECT 39.990 98.950 40.270 99.230 ;
        RECT 41.310 99.470 41.590 99.750 ;
        RECT 41.310 98.950 41.590 99.230 ;
        RECT 47.910 99.470 48.190 99.750 ;
        RECT 47.910 98.950 48.190 99.230 ;
        RECT 49.230 99.470 49.510 99.750 ;
        RECT 49.230 98.950 49.510 99.230 ;
        RECT 86.750 99.470 87.030 99.750 ;
        RECT 86.750 98.950 87.030 99.230 ;
        RECT 88.070 99.470 88.350 99.750 ;
        RECT 88.070 98.950 88.350 99.230 ;
        RECT 94.670 99.470 94.950 99.750 ;
        RECT 94.670 98.950 94.950 99.230 ;
        RECT 95.990 99.470 96.270 99.750 ;
        RECT 95.990 98.950 96.270 99.230 ;
        RECT 107.870 99.470 108.150 99.750 ;
        RECT 107.870 98.950 108.150 99.230 ;
        RECT 109.190 99.470 109.470 99.750 ;
        RECT 109.190 98.950 109.470 99.230 ;
        RECT 115.790 99.470 116.070 99.750 ;
        RECT 115.790 98.950 116.070 99.230 ;
        RECT 117.110 99.470 117.390 99.750 ;
        RECT 117.110 98.950 117.390 99.230 ;
        RECT 12.270 97.500 12.550 97.780 ;
        RECT 12.270 96.980 12.550 97.260 ;
        RECT 123.710 97.500 123.990 97.780 ;
        RECT 123.710 96.980 123.990 97.260 ;
        RECT 24.150 96.450 24.430 96.730 ;
        RECT 24.150 95.930 24.430 96.210 ;
        RECT 43.950 96.450 44.230 96.730 ;
        RECT 43.950 95.930 44.230 96.210 ;
        RECT 92.030 96.450 92.310 96.730 ;
        RECT 92.030 95.930 92.310 96.210 ;
        RECT 111.830 96.450 112.110 96.730 ;
        RECT 111.830 95.930 112.110 96.210 ;
        RECT 13.590 93.430 13.870 93.710 ;
        RECT 13.590 92.910 13.870 93.190 ;
        RECT 14.910 93.430 15.190 93.710 ;
        RECT 14.910 92.910 15.190 93.190 ;
        RECT 16.230 93.430 16.510 93.710 ;
        RECT 16.230 92.910 16.510 93.190 ;
        RECT 17.550 93.430 17.830 93.710 ;
        RECT 17.550 92.910 17.830 93.190 ;
        RECT 29.430 93.430 29.710 93.710 ;
        RECT 29.430 92.910 29.710 93.190 ;
        RECT 30.750 93.430 31.030 93.710 ;
        RECT 30.750 92.910 31.030 93.190 ;
        RECT 32.070 93.430 32.350 93.710 ;
        RECT 32.070 92.910 32.350 93.190 ;
        RECT 33.390 93.430 33.670 93.710 ;
        RECT 33.390 92.910 33.670 93.190 ;
        RECT 34.710 93.430 34.990 93.710 ;
        RECT 34.710 92.910 34.990 93.190 ;
        RECT 36.030 93.430 36.310 93.710 ;
        RECT 36.030 92.910 36.310 93.190 ;
        RECT 37.350 93.430 37.630 93.710 ;
        RECT 37.350 92.910 37.630 93.190 ;
        RECT 38.670 93.430 38.950 93.710 ;
        RECT 38.670 92.910 38.950 93.190 ;
        RECT 50.550 93.430 50.830 93.710 ;
        RECT 50.550 92.910 50.830 93.190 ;
        RECT 51.870 93.430 52.150 93.710 ;
        RECT 51.870 92.910 52.150 93.190 ;
        RECT 53.190 93.430 53.470 93.710 ;
        RECT 53.190 92.910 53.470 93.190 ;
        RECT 54.510 93.430 54.790 93.710 ;
        RECT 54.510 92.910 54.790 93.190 ;
        RECT 81.470 93.430 81.750 93.710 ;
        RECT 81.470 92.910 81.750 93.190 ;
        RECT 82.790 93.430 83.070 93.710 ;
        RECT 82.790 92.910 83.070 93.190 ;
        RECT 84.110 93.430 84.390 93.710 ;
        RECT 84.110 92.910 84.390 93.190 ;
        RECT 85.430 93.430 85.710 93.710 ;
        RECT 85.430 92.910 85.710 93.190 ;
        RECT 97.310 93.430 97.590 93.710 ;
        RECT 97.310 92.910 97.590 93.190 ;
        RECT 98.630 93.430 98.910 93.710 ;
        RECT 98.630 92.910 98.910 93.190 ;
        RECT 99.950 93.430 100.230 93.710 ;
        RECT 99.950 92.910 100.230 93.190 ;
        RECT 101.270 93.430 101.550 93.710 ;
        RECT 101.270 92.910 101.550 93.190 ;
        RECT 102.590 93.430 102.870 93.710 ;
        RECT 102.590 92.910 102.870 93.190 ;
        RECT 103.910 93.430 104.190 93.710 ;
        RECT 103.910 92.910 104.190 93.190 ;
        RECT 105.230 93.430 105.510 93.710 ;
        RECT 105.230 92.910 105.510 93.190 ;
        RECT 106.550 93.430 106.830 93.710 ;
        RECT 106.550 92.910 106.830 93.190 ;
        RECT 118.430 93.430 118.710 93.710 ;
        RECT 118.430 92.910 118.710 93.190 ;
        RECT 119.750 93.430 120.030 93.710 ;
        RECT 119.750 92.910 120.030 93.190 ;
        RECT 121.070 93.430 121.350 93.710 ;
        RECT 121.070 92.910 121.350 93.190 ;
        RECT 122.390 93.430 122.670 93.710 ;
        RECT 122.390 92.910 122.670 93.190 ;
        RECT 45.270 90.410 45.550 90.690 ;
        RECT 45.270 89.890 45.550 90.170 ;
        RECT 90.710 90.410 90.990 90.690 ;
        RECT 90.710 89.890 90.990 90.170 ;
        RECT 22.830 88.510 23.110 88.790 ;
        RECT 22.830 87.990 23.110 88.270 ;
        RECT 113.150 88.510 113.430 88.790 ;
        RECT 113.150 87.990 113.430 88.270 ;
        RECT 21.510 85.490 21.790 85.770 ;
        RECT 21.510 84.970 21.790 85.250 ;
        RECT 25.470 85.490 25.750 85.770 ;
        RECT 25.470 84.970 25.750 85.250 ;
        RECT 42.630 85.490 42.910 85.770 ;
        RECT 42.630 84.970 42.910 85.250 ;
        RECT 46.590 85.490 46.870 85.770 ;
        RECT 46.590 84.970 46.870 85.250 ;
        RECT 89.390 85.490 89.670 85.770 ;
        RECT 89.390 84.970 89.670 85.250 ;
        RECT 93.350 85.490 93.630 85.770 ;
        RECT 93.350 84.970 93.630 85.250 ;
        RECT 110.510 85.490 110.790 85.770 ;
        RECT 110.510 84.970 110.790 85.250 ;
        RECT 114.470 85.490 114.750 85.770 ;
        RECT 114.470 84.970 114.750 85.250 ;
        RECT 18.870 82.470 19.150 82.750 ;
        RECT 18.870 81.950 19.150 82.230 ;
        RECT 20.190 82.470 20.470 82.750 ;
        RECT 20.190 81.950 20.470 82.230 ;
        RECT 26.790 82.470 27.070 82.750 ;
        RECT 26.790 81.950 27.070 82.230 ;
        RECT 28.110 82.470 28.390 82.750 ;
        RECT 28.110 81.950 28.390 82.230 ;
        RECT 39.990 82.470 40.270 82.750 ;
        RECT 39.990 81.950 40.270 82.230 ;
        RECT 41.310 82.470 41.590 82.750 ;
        RECT 41.310 81.950 41.590 82.230 ;
        RECT 47.910 82.470 48.190 82.750 ;
        RECT 47.910 81.950 48.190 82.230 ;
        RECT 49.230 82.470 49.510 82.750 ;
        RECT 49.230 81.950 49.510 82.230 ;
        RECT 86.750 82.470 87.030 82.750 ;
        RECT 86.750 81.950 87.030 82.230 ;
        RECT 88.070 82.470 88.350 82.750 ;
        RECT 88.070 81.950 88.350 82.230 ;
        RECT 94.670 82.470 94.950 82.750 ;
        RECT 94.670 81.950 94.950 82.230 ;
        RECT 95.990 82.470 96.270 82.750 ;
        RECT 95.990 81.950 96.270 82.230 ;
        RECT 107.870 82.470 108.150 82.750 ;
        RECT 107.870 81.950 108.150 82.230 ;
        RECT 109.190 82.470 109.470 82.750 ;
        RECT 109.190 81.950 109.470 82.230 ;
        RECT 115.790 82.470 116.070 82.750 ;
        RECT 115.790 81.950 116.070 82.230 ;
        RECT 117.110 82.470 117.390 82.750 ;
        RECT 117.110 81.950 117.390 82.230 ;
        RECT 12.270 80.500 12.550 80.780 ;
        RECT 12.270 79.980 12.550 80.260 ;
        RECT 123.710 80.500 123.990 80.780 ;
        RECT 123.710 79.980 123.990 80.260 ;
        RECT 24.150 79.450 24.430 79.730 ;
        RECT 24.150 78.930 24.430 79.210 ;
        RECT 43.950 79.450 44.230 79.730 ;
        RECT 43.950 78.930 44.230 79.210 ;
        RECT 92.030 79.450 92.310 79.730 ;
        RECT 92.030 78.930 92.310 79.210 ;
        RECT 111.830 79.450 112.110 79.730 ;
        RECT 111.830 78.930 112.110 79.210 ;
        RECT 13.590 76.430 13.870 76.710 ;
        RECT 13.590 75.910 13.870 76.190 ;
        RECT 14.910 76.430 15.190 76.710 ;
        RECT 14.910 75.910 15.190 76.190 ;
        RECT 16.230 76.430 16.510 76.710 ;
        RECT 16.230 75.910 16.510 76.190 ;
        RECT 17.550 76.430 17.830 76.710 ;
        RECT 17.550 75.910 17.830 76.190 ;
        RECT 29.430 76.430 29.710 76.710 ;
        RECT 29.430 75.910 29.710 76.190 ;
        RECT 30.750 76.430 31.030 76.710 ;
        RECT 30.750 75.910 31.030 76.190 ;
        RECT 32.070 76.430 32.350 76.710 ;
        RECT 32.070 75.910 32.350 76.190 ;
        RECT 33.390 76.430 33.670 76.710 ;
        RECT 33.390 75.910 33.670 76.190 ;
        RECT 34.710 76.430 34.990 76.710 ;
        RECT 34.710 75.910 34.990 76.190 ;
        RECT 36.030 76.430 36.310 76.710 ;
        RECT 36.030 75.910 36.310 76.190 ;
        RECT 37.350 76.430 37.630 76.710 ;
        RECT 37.350 75.910 37.630 76.190 ;
        RECT 38.670 76.430 38.950 76.710 ;
        RECT 38.670 75.910 38.950 76.190 ;
        RECT 50.550 76.430 50.830 76.710 ;
        RECT 50.550 75.910 50.830 76.190 ;
        RECT 51.870 76.430 52.150 76.710 ;
        RECT 51.870 75.910 52.150 76.190 ;
        RECT 53.190 76.430 53.470 76.710 ;
        RECT 53.190 75.910 53.470 76.190 ;
        RECT 54.510 76.430 54.790 76.710 ;
        RECT 54.510 75.910 54.790 76.190 ;
        RECT 81.470 76.430 81.750 76.710 ;
        RECT 81.470 75.910 81.750 76.190 ;
        RECT 82.790 76.430 83.070 76.710 ;
        RECT 82.790 75.910 83.070 76.190 ;
        RECT 84.110 76.430 84.390 76.710 ;
        RECT 84.110 75.910 84.390 76.190 ;
        RECT 85.430 76.430 85.710 76.710 ;
        RECT 85.430 75.910 85.710 76.190 ;
        RECT 97.310 76.430 97.590 76.710 ;
        RECT 97.310 75.910 97.590 76.190 ;
        RECT 98.630 76.430 98.910 76.710 ;
        RECT 98.630 75.910 98.910 76.190 ;
        RECT 99.950 76.430 100.230 76.710 ;
        RECT 99.950 75.910 100.230 76.190 ;
        RECT 101.270 76.430 101.550 76.710 ;
        RECT 101.270 75.910 101.550 76.190 ;
        RECT 102.590 76.430 102.870 76.710 ;
        RECT 102.590 75.910 102.870 76.190 ;
        RECT 103.910 76.430 104.190 76.710 ;
        RECT 103.910 75.910 104.190 76.190 ;
        RECT 105.230 76.430 105.510 76.710 ;
        RECT 105.230 75.910 105.510 76.190 ;
        RECT 106.550 76.430 106.830 76.710 ;
        RECT 106.550 75.910 106.830 76.190 ;
        RECT 118.430 76.430 118.710 76.710 ;
        RECT 118.430 75.910 118.710 76.190 ;
        RECT 119.750 76.430 120.030 76.710 ;
        RECT 119.750 75.910 120.030 76.190 ;
        RECT 121.070 76.430 121.350 76.710 ;
        RECT 121.070 75.910 121.350 76.190 ;
        RECT 122.390 76.430 122.670 76.710 ;
        RECT 122.390 75.910 122.670 76.190 ;
        RECT 45.270 73.410 45.550 73.690 ;
        RECT 45.270 72.890 45.550 73.170 ;
        RECT 90.710 73.410 90.990 73.690 ;
        RECT 90.710 72.890 90.990 73.170 ;
        RECT 22.830 71.510 23.110 71.790 ;
        RECT 22.830 70.990 23.110 71.270 ;
        RECT 113.150 71.510 113.430 71.790 ;
        RECT 113.150 70.990 113.430 71.270 ;
        RECT 21.510 68.490 21.790 68.770 ;
        RECT 21.510 67.970 21.790 68.250 ;
        RECT 25.470 68.490 25.750 68.770 ;
        RECT 25.470 67.970 25.750 68.250 ;
        RECT 42.630 68.490 42.910 68.770 ;
        RECT 42.630 67.970 42.910 68.250 ;
        RECT 46.590 68.490 46.870 68.770 ;
        RECT 46.590 67.970 46.870 68.250 ;
        RECT 89.390 68.490 89.670 68.770 ;
        RECT 89.390 67.970 89.670 68.250 ;
        RECT 93.350 68.490 93.630 68.770 ;
        RECT 93.350 67.970 93.630 68.250 ;
        RECT 110.510 68.490 110.790 68.770 ;
        RECT 110.510 67.970 110.790 68.250 ;
        RECT 114.470 68.490 114.750 68.770 ;
        RECT 114.470 67.970 114.750 68.250 ;
        RECT 18.870 65.470 19.150 65.750 ;
        RECT 18.870 64.950 19.150 65.230 ;
        RECT 20.190 65.470 20.470 65.750 ;
        RECT 20.190 64.950 20.470 65.230 ;
        RECT 26.790 65.470 27.070 65.750 ;
        RECT 26.790 64.950 27.070 65.230 ;
        RECT 28.110 65.470 28.390 65.750 ;
        RECT 28.110 64.950 28.390 65.230 ;
        RECT 39.990 65.470 40.270 65.750 ;
        RECT 39.990 64.950 40.270 65.230 ;
        RECT 41.310 65.470 41.590 65.750 ;
        RECT 41.310 64.950 41.590 65.230 ;
        RECT 47.910 65.470 48.190 65.750 ;
        RECT 47.910 64.950 48.190 65.230 ;
        RECT 49.230 65.470 49.510 65.750 ;
        RECT 49.230 64.950 49.510 65.230 ;
        RECT 86.750 65.470 87.030 65.750 ;
        RECT 86.750 64.950 87.030 65.230 ;
        RECT 88.070 65.470 88.350 65.750 ;
        RECT 88.070 64.950 88.350 65.230 ;
        RECT 94.670 65.470 94.950 65.750 ;
        RECT 94.670 64.950 94.950 65.230 ;
        RECT 95.990 65.470 96.270 65.750 ;
        RECT 95.990 64.950 96.270 65.230 ;
        RECT 107.870 65.470 108.150 65.750 ;
        RECT 107.870 64.950 108.150 65.230 ;
        RECT 109.190 65.470 109.470 65.750 ;
        RECT 109.190 64.950 109.470 65.230 ;
        RECT 115.790 65.470 116.070 65.750 ;
        RECT 115.790 64.950 116.070 65.230 ;
        RECT 117.110 65.470 117.390 65.750 ;
        RECT 117.110 64.950 117.390 65.230 ;
        RECT 12.270 63.500 12.550 63.780 ;
        RECT 12.270 62.980 12.550 63.260 ;
        RECT 123.710 63.500 123.990 63.780 ;
        RECT 123.710 62.980 123.990 63.260 ;
        RECT 24.150 62.450 24.430 62.730 ;
        RECT 24.150 61.930 24.430 62.210 ;
        RECT 43.950 62.450 44.230 62.730 ;
        RECT 43.950 61.930 44.230 62.210 ;
        RECT 92.030 62.450 92.310 62.730 ;
        RECT 92.030 61.930 92.310 62.210 ;
        RECT 111.830 62.450 112.110 62.730 ;
        RECT 111.830 61.930 112.110 62.210 ;
        RECT 13.590 59.430 13.870 59.710 ;
        RECT 13.590 58.910 13.870 59.190 ;
        RECT 14.910 59.430 15.190 59.710 ;
        RECT 14.910 58.910 15.190 59.190 ;
        RECT 16.230 59.430 16.510 59.710 ;
        RECT 16.230 58.910 16.510 59.190 ;
        RECT 17.550 59.430 17.830 59.710 ;
        RECT 17.550 58.910 17.830 59.190 ;
        RECT 29.430 59.430 29.710 59.710 ;
        RECT 29.430 58.910 29.710 59.190 ;
        RECT 30.750 59.430 31.030 59.710 ;
        RECT 30.750 58.910 31.030 59.190 ;
        RECT 32.070 59.430 32.350 59.710 ;
        RECT 32.070 58.910 32.350 59.190 ;
        RECT 33.390 59.430 33.670 59.710 ;
        RECT 33.390 58.910 33.670 59.190 ;
        RECT 34.710 59.430 34.990 59.710 ;
        RECT 34.710 58.910 34.990 59.190 ;
        RECT 36.030 59.430 36.310 59.710 ;
        RECT 36.030 58.910 36.310 59.190 ;
        RECT 37.350 59.430 37.630 59.710 ;
        RECT 37.350 58.910 37.630 59.190 ;
        RECT 38.670 59.430 38.950 59.710 ;
        RECT 38.670 58.910 38.950 59.190 ;
        RECT 50.550 59.430 50.830 59.710 ;
        RECT 50.550 58.910 50.830 59.190 ;
        RECT 51.870 59.430 52.150 59.710 ;
        RECT 51.870 58.910 52.150 59.190 ;
        RECT 53.190 59.430 53.470 59.710 ;
        RECT 53.190 58.910 53.470 59.190 ;
        RECT 54.510 59.430 54.790 59.710 ;
        RECT 54.510 58.910 54.790 59.190 ;
        RECT 81.470 59.430 81.750 59.710 ;
        RECT 81.470 58.910 81.750 59.190 ;
        RECT 82.790 59.430 83.070 59.710 ;
        RECT 82.790 58.910 83.070 59.190 ;
        RECT 84.110 59.430 84.390 59.710 ;
        RECT 84.110 58.910 84.390 59.190 ;
        RECT 85.430 59.430 85.710 59.710 ;
        RECT 85.430 58.910 85.710 59.190 ;
        RECT 97.310 59.430 97.590 59.710 ;
        RECT 97.310 58.910 97.590 59.190 ;
        RECT 98.630 59.430 98.910 59.710 ;
        RECT 98.630 58.910 98.910 59.190 ;
        RECT 99.950 59.430 100.230 59.710 ;
        RECT 99.950 58.910 100.230 59.190 ;
        RECT 101.270 59.430 101.550 59.710 ;
        RECT 101.270 58.910 101.550 59.190 ;
        RECT 102.590 59.430 102.870 59.710 ;
        RECT 102.590 58.910 102.870 59.190 ;
        RECT 103.910 59.430 104.190 59.710 ;
        RECT 103.910 58.910 104.190 59.190 ;
        RECT 105.230 59.430 105.510 59.710 ;
        RECT 105.230 58.910 105.510 59.190 ;
        RECT 106.550 59.430 106.830 59.710 ;
        RECT 106.550 58.910 106.830 59.190 ;
        RECT 118.430 59.430 118.710 59.710 ;
        RECT 118.430 58.910 118.710 59.190 ;
        RECT 119.750 59.430 120.030 59.710 ;
        RECT 119.750 58.910 120.030 59.190 ;
        RECT 121.070 59.430 121.350 59.710 ;
        RECT 121.070 58.910 121.350 59.190 ;
        RECT 122.390 59.430 122.670 59.710 ;
        RECT 122.390 58.910 122.670 59.190 ;
        RECT 45.270 56.410 45.550 56.690 ;
        RECT 45.270 55.890 45.550 56.170 ;
        RECT 90.710 56.410 90.990 56.690 ;
        RECT 90.710 55.890 90.990 56.170 ;
        RECT 22.830 54.510 23.110 54.790 ;
        RECT 22.830 53.990 23.110 54.270 ;
        RECT 113.150 54.510 113.430 54.790 ;
        RECT 113.150 53.990 113.430 54.270 ;
        RECT 21.510 51.490 21.790 51.770 ;
        RECT 21.510 50.970 21.790 51.250 ;
        RECT 25.470 51.490 25.750 51.770 ;
        RECT 25.470 50.970 25.750 51.250 ;
        RECT 42.630 51.490 42.910 51.770 ;
        RECT 42.630 50.970 42.910 51.250 ;
        RECT 46.590 51.490 46.870 51.770 ;
        RECT 46.590 50.970 46.870 51.250 ;
        RECT 89.390 51.490 89.670 51.770 ;
        RECT 89.390 50.970 89.670 51.250 ;
        RECT 93.350 51.490 93.630 51.770 ;
        RECT 93.350 50.970 93.630 51.250 ;
        RECT 110.510 51.490 110.790 51.770 ;
        RECT 110.510 50.970 110.790 51.250 ;
        RECT 114.470 51.490 114.750 51.770 ;
        RECT 114.470 50.970 114.750 51.250 ;
        RECT 18.870 48.470 19.150 48.750 ;
        RECT 18.870 47.950 19.150 48.230 ;
        RECT 20.190 48.470 20.470 48.750 ;
        RECT 20.190 47.950 20.470 48.230 ;
        RECT 26.790 48.470 27.070 48.750 ;
        RECT 26.790 47.950 27.070 48.230 ;
        RECT 28.110 48.470 28.390 48.750 ;
        RECT 28.110 47.950 28.390 48.230 ;
        RECT 39.990 48.470 40.270 48.750 ;
        RECT 39.990 47.950 40.270 48.230 ;
        RECT 41.310 48.470 41.590 48.750 ;
        RECT 41.310 47.950 41.590 48.230 ;
        RECT 47.910 48.470 48.190 48.750 ;
        RECT 47.910 47.950 48.190 48.230 ;
        RECT 49.230 48.470 49.510 48.750 ;
        RECT 49.230 47.950 49.510 48.230 ;
        RECT 86.750 48.470 87.030 48.750 ;
        RECT 86.750 47.950 87.030 48.230 ;
        RECT 88.070 48.470 88.350 48.750 ;
        RECT 88.070 47.950 88.350 48.230 ;
        RECT 94.670 48.470 94.950 48.750 ;
        RECT 94.670 47.950 94.950 48.230 ;
        RECT 95.990 48.470 96.270 48.750 ;
        RECT 95.990 47.950 96.270 48.230 ;
        RECT 107.870 48.470 108.150 48.750 ;
        RECT 107.870 47.950 108.150 48.230 ;
        RECT 109.190 48.470 109.470 48.750 ;
        RECT 109.190 47.950 109.470 48.230 ;
        RECT 115.790 48.470 116.070 48.750 ;
        RECT 115.790 47.950 116.070 48.230 ;
        RECT 117.110 48.470 117.390 48.750 ;
        RECT 117.110 47.950 117.390 48.230 ;
        RECT 12.270 46.500 12.550 46.780 ;
        RECT 12.270 45.980 12.550 46.260 ;
        RECT 123.710 46.500 123.990 46.780 ;
        RECT 123.710 45.980 123.990 46.260 ;
        RECT 24.150 45.450 24.430 45.730 ;
        RECT 24.150 44.930 24.430 45.210 ;
        RECT 43.950 45.450 44.230 45.730 ;
        RECT 43.950 44.930 44.230 45.210 ;
        RECT 92.030 45.450 92.310 45.730 ;
        RECT 92.030 44.930 92.310 45.210 ;
        RECT 111.830 45.450 112.110 45.730 ;
        RECT 111.830 44.930 112.110 45.210 ;
        RECT 13.590 42.430 13.870 42.710 ;
        RECT 13.590 41.910 13.870 42.190 ;
        RECT 14.910 42.430 15.190 42.710 ;
        RECT 14.910 41.910 15.190 42.190 ;
        RECT 16.230 42.430 16.510 42.710 ;
        RECT 16.230 41.910 16.510 42.190 ;
        RECT 17.550 42.430 17.830 42.710 ;
        RECT 17.550 41.910 17.830 42.190 ;
        RECT 29.430 42.430 29.710 42.710 ;
        RECT 29.430 41.910 29.710 42.190 ;
        RECT 30.750 42.430 31.030 42.710 ;
        RECT 30.750 41.910 31.030 42.190 ;
        RECT 32.070 42.430 32.350 42.710 ;
        RECT 32.070 41.910 32.350 42.190 ;
        RECT 33.390 42.430 33.670 42.710 ;
        RECT 33.390 41.910 33.670 42.190 ;
        RECT 34.710 42.430 34.990 42.710 ;
        RECT 34.710 41.910 34.990 42.190 ;
        RECT 36.030 42.430 36.310 42.710 ;
        RECT 36.030 41.910 36.310 42.190 ;
        RECT 37.350 42.430 37.630 42.710 ;
        RECT 37.350 41.910 37.630 42.190 ;
        RECT 38.670 42.430 38.950 42.710 ;
        RECT 38.670 41.910 38.950 42.190 ;
        RECT 50.550 42.430 50.830 42.710 ;
        RECT 50.550 41.910 50.830 42.190 ;
        RECT 51.870 42.430 52.150 42.710 ;
        RECT 51.870 41.910 52.150 42.190 ;
        RECT 53.190 42.430 53.470 42.710 ;
        RECT 53.190 41.910 53.470 42.190 ;
        RECT 54.510 42.430 54.790 42.710 ;
        RECT 54.510 41.910 54.790 42.190 ;
        RECT 81.470 42.430 81.750 42.710 ;
        RECT 81.470 41.910 81.750 42.190 ;
        RECT 82.790 42.430 83.070 42.710 ;
        RECT 82.790 41.910 83.070 42.190 ;
        RECT 84.110 42.430 84.390 42.710 ;
        RECT 84.110 41.910 84.390 42.190 ;
        RECT 85.430 42.430 85.710 42.710 ;
        RECT 85.430 41.910 85.710 42.190 ;
        RECT 97.310 42.430 97.590 42.710 ;
        RECT 97.310 41.910 97.590 42.190 ;
        RECT 98.630 42.430 98.910 42.710 ;
        RECT 98.630 41.910 98.910 42.190 ;
        RECT 99.950 42.430 100.230 42.710 ;
        RECT 99.950 41.910 100.230 42.190 ;
        RECT 101.270 42.430 101.550 42.710 ;
        RECT 101.270 41.910 101.550 42.190 ;
        RECT 102.590 42.430 102.870 42.710 ;
        RECT 102.590 41.910 102.870 42.190 ;
        RECT 103.910 42.430 104.190 42.710 ;
        RECT 103.910 41.910 104.190 42.190 ;
        RECT 105.230 42.430 105.510 42.710 ;
        RECT 105.230 41.910 105.510 42.190 ;
        RECT 106.550 42.430 106.830 42.710 ;
        RECT 106.550 41.910 106.830 42.190 ;
        RECT 118.430 42.430 118.710 42.710 ;
        RECT 118.430 41.910 118.710 42.190 ;
        RECT 119.750 42.430 120.030 42.710 ;
        RECT 119.750 41.910 120.030 42.190 ;
        RECT 121.070 42.430 121.350 42.710 ;
        RECT 121.070 41.910 121.350 42.190 ;
        RECT 122.390 42.430 122.670 42.710 ;
        RECT 122.390 41.910 122.670 42.190 ;
        RECT 45.270 39.410 45.550 39.690 ;
        RECT 45.270 38.890 45.550 39.170 ;
        RECT 90.710 39.410 90.990 39.690 ;
        RECT 90.710 38.890 90.990 39.170 ;
        RECT 44.550 36.280 45.630 36.600 ;
        RECT 11.790 35.480 12.870 35.800 ;
        RECT 44.550 34.680 45.630 35.000 ;
        RECT 11.790 33.880 12.870 34.200 ;
        RECT 44.550 33.080 45.630 33.400 ;
        RECT 90.630 36.280 91.710 36.600 ;
        RECT 123.390 35.480 124.470 35.800 ;
        RECT 90.630 34.680 91.710 35.000 ;
        RECT 123.390 33.880 124.470 34.200 ;
        RECT 90.630 33.080 91.710 33.400 ;
        RECT 11.790 32.280 12.870 32.600 ;
        RECT 123.390 32.280 124.470 32.600 ;
        RECT 44.550 31.480 45.630 31.800 ;
        RECT 11.790 30.680 12.870 31.000 ;
        RECT 44.550 29.880 45.630 30.200 ;
        RECT 11.790 29.080 12.870 29.400 ;
        RECT 90.630 31.480 91.710 31.800 ;
        RECT 123.390 30.680 124.470 31.000 ;
        RECT 90.630 29.880 91.710 30.200 ;
        RECT 52.330 29.380 52.610 29.660 ;
        RECT 52.850 29.380 53.130 29.660 ;
        RECT 56.290 29.380 56.570 29.660 ;
        RECT 56.810 29.380 57.090 29.660 ;
        RECT 79.170 29.380 79.450 29.660 ;
        RECT 79.690 29.380 79.970 29.660 ;
        RECT 83.130 29.380 83.410 29.660 ;
        RECT 83.650 29.380 83.930 29.660 ;
        RECT 44.550 28.280 45.630 28.600 ;
        RECT 52.330 28.500 52.610 28.780 ;
        RECT 52.850 28.500 53.130 28.780 ;
        RECT 56.290 28.500 56.570 28.780 ;
        RECT 56.810 28.500 57.090 28.780 ;
        RECT 79.170 28.500 79.450 28.780 ;
        RECT 79.690 28.500 79.970 28.780 ;
        RECT 83.130 28.500 83.410 28.780 ;
        RECT 83.650 28.500 83.930 28.780 ;
        RECT 123.390 29.080 124.470 29.400 ;
        RECT 90.630 28.280 91.710 28.600 ;
        RECT 11.790 27.480 12.870 27.800 ;
        RECT 58.890 27.620 59.170 27.900 ;
        RECT 59.410 27.620 59.690 27.900 ;
        RECT 76.570 27.620 76.850 27.900 ;
        RECT 77.090 27.620 77.370 27.900 ;
        RECT 123.390 27.480 124.470 27.800 ;
        RECT 44.550 26.680 45.630 27.000 ;
        RECT 52.330 26.740 52.610 27.020 ;
        RECT 52.850 26.740 53.130 27.020 ;
        RECT 56.290 26.740 56.570 27.020 ;
        RECT 56.810 26.740 57.090 27.020 ;
        RECT 79.170 26.740 79.450 27.020 ;
        RECT 79.690 26.740 79.970 27.020 ;
        RECT 83.130 26.740 83.410 27.020 ;
        RECT 83.650 26.740 83.930 27.020 ;
        RECT 11.790 25.880 12.870 26.200 ;
        RECT 90.630 26.680 91.710 27.000 ;
        RECT 52.330 25.860 52.610 26.140 ;
        RECT 52.850 25.860 53.130 26.140 ;
        RECT 56.290 25.860 56.570 26.140 ;
        RECT 56.810 25.860 57.090 26.140 ;
        RECT 71.970 25.860 72.250 26.140 ;
        RECT 72.490 25.860 72.770 26.140 ;
        RECT 79.170 25.860 79.450 26.140 ;
        RECT 79.690 25.860 79.970 26.140 ;
        RECT 83.130 25.860 83.410 26.140 ;
        RECT 83.650 25.860 83.930 26.140 ;
        RECT 44.550 25.080 45.630 25.400 ;
        RECT 11.790 24.280 12.870 24.600 ;
        RECT 52.330 24.980 52.610 25.260 ;
        RECT 52.850 24.980 53.130 25.260 ;
        RECT 56.290 24.980 56.570 25.260 ;
        RECT 56.810 24.980 57.090 25.260 ;
        RECT 44.550 23.480 45.630 23.800 ;
        RECT 52.330 23.220 52.610 23.500 ;
        RECT 52.850 23.220 53.130 23.500 ;
        RECT 56.290 23.220 56.570 23.500 ;
        RECT 56.810 23.220 57.090 23.500 ;
        RECT 11.790 22.680 12.870 23.000 ;
        RECT 52.330 22.340 52.610 22.620 ;
        RECT 52.850 22.340 53.130 22.620 ;
        RECT 44.550 21.880 45.630 22.200 ;
        RECT 11.790 21.080 12.870 21.400 ;
        RECT 50.170 21.460 50.450 21.740 ;
        RECT 50.690 21.460 50.970 21.740 ;
        RECT 44.550 20.280 45.630 20.600 ;
        RECT 56.290 20.580 56.570 20.860 ;
        RECT 56.810 20.580 57.090 20.860 ;
        RECT 11.790 19.480 12.870 19.800 ;
        RECT 44.550 18.680 45.630 19.000 ;
        RECT 50.170 18.380 50.450 18.660 ;
        RECT 50.690 18.380 50.970 18.660 ;
        RECT 11.790 17.880 12.870 18.200 ;
        RECT 44.550 17.080 45.630 17.400 ;
        RECT 11.790 16.280 12.870 16.600 ;
        RECT 44.550 15.480 45.630 15.800 ;
        RECT 11.790 14.680 12.870 15.000 ;
        RECT 44.550 13.880 45.630 14.200 ;
        RECT 11.790 13.080 12.870 13.400 ;
        RECT 52.330 17.940 52.610 18.220 ;
        RECT 52.850 17.940 53.130 18.220 ;
        RECT 56.290 17.940 56.570 18.220 ;
        RECT 56.810 17.940 57.090 18.220 ;
        RECT 123.390 25.880 124.470 26.200 ;
        RECT 79.170 24.980 79.450 25.260 ;
        RECT 79.690 24.980 79.970 25.260 ;
        RECT 83.130 24.980 83.410 25.260 ;
        RECT 83.650 24.980 83.930 25.260 ;
        RECT 90.630 25.080 91.710 25.400 ;
        RECT 123.390 24.280 124.470 24.600 ;
        RECT 79.170 23.220 79.450 23.500 ;
        RECT 79.690 23.220 79.970 23.500 ;
        RECT 83.130 23.220 83.410 23.500 ;
        RECT 83.650 23.220 83.930 23.500 ;
        RECT 90.630 23.480 91.710 23.800 ;
        RECT 123.390 22.680 124.470 23.000 ;
        RECT 83.130 22.340 83.410 22.620 ;
        RECT 83.650 22.340 83.930 22.620 ;
        RECT 63.330 18.820 63.610 19.100 ;
        RECT 63.850 18.820 64.130 19.100 ;
        RECT 71.970 18.820 72.250 19.100 ;
        RECT 72.490 18.820 72.770 19.100 ;
        RECT 90.630 21.880 91.710 22.200 ;
        RECT 85.290 21.460 85.570 21.740 ;
        RECT 85.810 21.460 86.090 21.740 ;
        RECT 79.170 20.580 79.450 20.860 ;
        RECT 79.690 20.580 79.970 20.860 ;
        RECT 123.390 21.080 124.470 21.400 ;
        RECT 90.630 20.280 91.710 20.600 ;
        RECT 79.170 17.940 79.450 18.220 ;
        RECT 79.690 17.940 79.970 18.220 ;
        RECT 83.130 17.940 83.410 18.220 ;
        RECT 83.650 17.940 83.930 18.220 ;
        RECT 52.330 15.300 52.610 15.580 ;
        RECT 52.850 15.300 53.130 15.580 ;
        RECT 56.290 15.300 56.570 15.580 ;
        RECT 56.810 15.300 57.090 15.580 ;
        RECT 79.170 15.300 79.450 15.580 ;
        RECT 79.690 15.300 79.970 15.580 ;
        RECT 83.130 15.300 83.410 15.580 ;
        RECT 83.650 15.300 83.930 15.580 ;
        RECT 52.330 14.420 52.610 14.700 ;
        RECT 52.850 14.420 53.130 14.700 ;
        RECT 56.290 14.420 56.570 14.700 ;
        RECT 56.810 14.420 57.090 14.700 ;
        RECT 63.330 14.420 63.610 14.700 ;
        RECT 63.850 14.420 64.130 14.700 ;
        RECT 72.130 14.420 72.410 14.700 ;
        RECT 72.650 14.420 72.930 14.700 ;
        RECT 79.170 14.420 79.450 14.700 ;
        RECT 79.690 14.420 79.970 14.700 ;
        RECT 83.130 14.420 83.410 14.700 ;
        RECT 83.650 14.420 83.930 14.700 ;
        RECT 52.330 13.540 52.610 13.820 ;
        RECT 52.850 13.540 53.130 13.820 ;
        RECT 56.290 13.540 56.570 13.820 ;
        RECT 56.810 13.540 57.090 13.820 ;
        RECT 45.850 13.070 46.130 13.350 ;
        RECT 46.370 13.070 46.650 13.350 ;
        RECT 56.290 10.220 56.570 10.500 ;
        RECT 56.810 10.220 57.090 10.500 ;
        RECT 56.290 9.700 56.570 9.980 ;
        RECT 56.810 9.700 57.090 9.980 ;
        RECT 52.330 6.620 52.610 6.900 ;
        RECT 52.850 6.620 53.130 6.900 ;
        RECT 52.330 6.100 52.610 6.380 ;
        RECT 52.850 6.100 53.130 6.380 ;
        RECT 58.890 3.950 59.170 4.230 ;
        RECT 59.410 3.950 59.690 4.230 ;
        RECT 79.170 13.540 79.450 13.820 ;
        RECT 79.690 13.540 79.970 13.820 ;
        RECT 83.130 13.540 83.410 13.820 ;
        RECT 83.650 13.540 83.930 13.820 ;
        RECT 123.390 19.480 124.470 19.800 ;
        RECT 85.290 18.380 85.570 18.660 ;
        RECT 85.810 18.380 86.090 18.660 ;
        RECT 90.630 18.680 91.710 19.000 ;
        RECT 123.390 17.880 124.470 18.200 ;
        RECT 90.630 17.080 91.710 17.400 ;
        RECT 123.390 16.280 124.470 16.600 ;
        RECT 90.630 15.480 91.710 15.800 ;
        RECT 123.390 14.680 124.470 15.000 ;
        RECT 90.630 13.880 91.710 14.200 ;
        RECT 89.610 13.070 89.890 13.350 ;
        RECT 90.130 13.070 90.410 13.350 ;
        RECT 123.390 13.080 124.470 13.400 ;
        RECT 79.170 10.220 79.450 10.500 ;
        RECT 79.690 10.220 79.970 10.500 ;
        RECT 79.170 9.700 79.450 9.980 ;
        RECT 79.690 9.700 79.970 9.980 ;
        RECT 83.130 6.620 83.410 6.900 ;
        RECT 83.650 6.620 83.930 6.900 ;
        RECT 83.130 6.100 83.410 6.380 ;
        RECT 83.650 6.100 83.930 6.380 ;
        RECT 76.570 3.950 76.850 4.230 ;
        RECT 77.090 3.950 77.370 4.230 ;
        RECT 72.515 2.925 73.065 3.475 ;
        RECT 63.495 1.515 64.045 2.065 ;
      LAYER met3 ;
        RECT 29.710 224.615 30.090 224.625 ;
        RECT 57.470 224.615 57.905 224.685 ;
        RECT 29.710 224.315 57.905 224.615 ;
        RECT 59.150 224.360 60.010 224.690 ;
        RECT 61.605 224.440 61.955 224.485 ;
        RECT 86.865 224.440 87.195 224.455 ;
        RECT 29.710 224.305 30.090 224.315 ;
        RECT 57.470 224.275 57.905 224.315 ;
        RECT 61.090 224.140 87.195 224.440 ;
        RECT 61.605 224.135 61.955 224.140 ;
        RECT 86.865 224.125 87.195 224.140 ;
        RECT 88.590 224.250 88.970 224.260 ;
        RECT 108.035 224.250 108.365 224.265 ;
        RECT 88.590 223.950 108.365 224.250 ;
        RECT 88.590 223.940 88.970 223.950 ;
        RECT 108.035 223.935 108.365 223.950 ;
        RECT 34.890 223.780 35.270 223.790 ;
        RECT 35.985 223.780 36.335 223.805 ;
        RECT 34.890 223.480 36.335 223.780 ;
        RECT 34.890 223.470 35.270 223.480 ;
        RECT 35.985 223.455 36.335 223.480 ;
        RECT 40.835 223.750 41.165 223.765 ;
        RECT 70.190 223.750 70.570 223.760 ;
        RECT 40.835 223.450 70.570 223.750 ;
        RECT 40.835 223.435 41.165 223.450 ;
        RECT 70.190 223.440 70.570 223.450 ;
        RECT 84.910 223.550 85.290 223.560 ;
        RECT 91.235 223.550 91.565 223.565 ;
        RECT 84.910 223.250 91.565 223.550 ;
        RECT 84.910 223.240 85.290 223.250 ;
        RECT 91.235 223.235 91.565 223.250 ;
        RECT 111.315 223.005 111.645 223.335 ;
        RECT 114.470 223.320 114.810 223.470 ;
        RECT 15.735 222.950 16.065 222.965 ;
        RECT 55.810 222.950 56.190 222.960 ;
        RECT 15.735 222.650 56.190 222.950 ;
        RECT 15.735 222.635 16.065 222.650 ;
        RECT 55.810 222.640 56.190 222.650 ;
        RECT 57.535 222.950 57.865 222.965 ;
        RECT 73.870 222.950 74.250 222.960 ;
        RECT 57.535 222.650 74.250 222.950 ;
        RECT 57.535 222.635 57.865 222.650 ;
        RECT 73.870 222.640 74.250 222.650 ;
        RECT 81.260 222.950 81.580 222.990 ;
        RECT 82.635 222.950 82.965 222.965 ;
        RECT 81.260 222.650 82.965 222.950 ;
        RECT 81.260 222.610 81.580 222.650 ;
        RECT 82.635 222.635 82.965 222.650 ;
        RECT 32.335 222.250 32.665 222.265 ;
        RECT 64.310 222.250 64.690 222.260 ;
        RECT 32.335 221.950 64.690 222.250 ;
        RECT 32.335 221.935 32.665 221.950 ;
        RECT 64.310 221.940 64.690 221.950 ;
        RECT 66.035 222.250 66.365 222.265 ;
        RECT 77.550 222.250 77.930 222.260 ;
        RECT 66.035 221.950 77.930 222.250 ;
        RECT 66.035 221.935 66.365 221.950 ;
        RECT 77.550 221.940 77.930 221.950 ;
        RECT 79.400 222.040 79.750 222.065 ;
        RECT 111.330 222.040 111.630 223.005 ;
        RECT 79.400 221.740 111.630 222.040 ;
        RECT 114.470 222.980 135.030 223.320 ;
        RECT 114.470 221.810 114.810 222.980 ;
        RECT 79.400 221.715 79.750 221.740 ;
        RECT 113.950 221.470 115.670 221.810 ;
        RECT 15.310 199.070 16.230 220.930 ;
        RECT 13.205 157.120 13.555 197.975 ;
        RECT 19.270 197.630 20.190 220.930 ;
        RECT 22.050 197.400 22.970 198.550 ;
        RECT 25.090 197.400 26.010 198.550 ;
        RECT 28.070 197.630 28.990 220.930 ;
        RECT 22.050 197.120 26.010 197.400 ;
        RECT 22.050 195.620 26.050 197.120 ;
        RECT 31.055 195.670 31.395 196.230 ;
        RECT 22.050 195.500 26.010 195.620 ;
        RECT 19.170 193.160 20.090 194.950 ;
        RECT 22.050 193.160 22.970 195.500 ;
        RECT 25.090 193.160 26.010 195.500 ;
        RECT 30.730 195.130 31.395 195.670 ;
        RECT 27.970 193.160 28.890 194.950 ;
        RECT 19.170 192.240 28.890 193.160 ;
        RECT 13.205 156.780 14.130 157.120 ;
        RECT 13.205 146.375 13.555 156.780 ;
        RECT 13.210 112.390 13.550 146.375 ;
        RECT 15.210 134.070 16.130 191.590 ;
        RECT 16.660 115.180 17.000 157.850 ;
        RECT 17.375 121.690 17.715 162.250 ;
        RECT 18.160 124.480 18.500 166.650 ;
        RECT 19.170 134.070 20.090 192.240 ;
        RECT 22.050 153.700 22.970 192.240 ;
        RECT 25.090 153.700 26.010 192.240 ;
        RECT 27.970 134.070 28.890 192.240 ;
        RECT 29.560 125.410 29.900 166.650 ;
        RECT 30.345 161.330 30.685 162.250 ;
        RECT 30.340 122.620 30.680 161.330 ;
        RECT 31.055 157.850 31.395 195.130 ;
        RECT 32.030 191.590 32.950 220.930 ;
        RECT 34.330 195.595 34.670 197.970 ;
        RECT 38.830 195.595 39.170 197.870 ;
        RECT 34.305 195.205 34.695 195.595 ;
        RECT 38.805 195.205 39.195 195.595 ;
        RECT 31.930 190.440 32.950 191.590 ;
        RECT 40.510 191.390 41.430 220.930 ;
        RECT 44.470 197.630 45.390 220.930 ;
        RECT 47.250 197.120 48.170 198.550 ;
        RECT 50.290 197.120 51.210 198.550 ;
        RECT 53.270 197.630 54.190 220.930 ;
        RECT 31.055 156.930 31.400 157.850 ;
        RECT 31.055 116.110 31.395 156.930 ;
        RECT 31.930 134.070 32.850 190.440 ;
        RECT 40.410 189.940 41.430 191.390 ;
        RECT 33.930 156.780 34.850 157.120 ;
        RECT 38.410 156.780 39.330 157.120 ;
        RECT 33.930 113.320 34.270 156.780 ;
        RECT 38.410 114.250 38.750 156.780 ;
        RECT 40.410 134.070 41.330 189.940 ;
        RECT 41.860 117.040 42.200 196.430 ;
        RECT 47.250 195.620 51.350 197.120 ;
        RECT 44.370 193.060 45.290 194.950 ;
        RECT 47.250 193.060 48.170 195.620 ;
        RECT 50.290 193.060 51.210 195.620 ;
        RECT 53.170 193.060 54.090 194.950 ;
        RECT 44.370 192.140 54.090 193.060 ;
        RECT 42.575 123.550 42.915 162.250 ;
        RECT 43.360 126.340 43.700 166.650 ;
        RECT 44.370 134.070 45.290 192.140 ;
        RECT 47.250 153.700 48.170 192.140 ;
        RECT 50.290 153.700 51.210 192.140 ;
        RECT 53.170 134.070 54.090 192.140 ;
        RECT 54.760 127.270 55.100 166.650 ;
        RECT 55.545 161.330 55.885 162.250 ;
        RECT 56.255 157.850 56.595 195.630 ;
        RECT 57.230 191.690 58.150 220.930 ;
        RECT 59.630 195.495 59.970 198.070 ;
        RECT 63.930 195.495 64.270 198.070 ;
        RECT 59.605 195.105 59.995 195.495 ;
        RECT 63.905 195.105 64.295 195.495 ;
        RECT 57.130 190.540 58.150 191.690 ;
        RECT 65.710 191.350 66.630 220.930 ;
        RECT 69.670 197.630 70.590 220.930 ;
        RECT 72.450 197.300 73.370 198.550 ;
        RECT 75.490 197.300 76.410 198.550 ;
        RECT 78.470 197.630 79.390 220.930 ;
        RECT 56.255 156.930 56.600 157.850 ;
        RECT 56.255 117.970 56.595 156.930 ;
        RECT 57.130 134.070 58.050 190.540 ;
        RECT 65.610 190.240 66.630 191.350 ;
        RECT 59.130 156.780 60.050 157.120 ;
        RECT 63.610 156.780 64.530 157.120 ;
        RECT 65.610 134.070 66.530 190.240 ;
        RECT 67.060 118.900 67.400 195.930 ;
        RECT 72.450 195.500 76.410 197.300 ;
        RECT 81.455 195.595 81.795 196.330 ;
        RECT 69.570 193.260 70.490 194.950 ;
        RECT 72.450 193.260 73.370 195.500 ;
        RECT 75.490 193.260 76.410 195.500 ;
        RECT 81.405 195.205 81.795 195.595 ;
        RECT 78.370 193.260 79.290 194.950 ;
        RECT 69.570 192.340 79.290 193.260 ;
        RECT 67.775 161.330 68.115 162.250 ;
        RECT 68.560 128.200 68.900 166.650 ;
        RECT 69.570 134.070 70.490 192.340 ;
        RECT 72.450 153.700 73.370 192.340 ;
        RECT 75.490 153.700 76.410 192.340 ;
        RECT 78.370 134.070 79.290 192.340 ;
        RECT 79.960 129.130 80.300 166.650 ;
        RECT 80.745 161.330 81.085 162.250 ;
        RECT 81.455 157.850 81.795 195.205 ;
        RECT 82.430 191.490 83.350 220.930 ;
        RECT 84.730 195.230 85.070 198.070 ;
        RECT 89.130 195.495 89.470 198.070 ;
        RECT 89.105 195.105 89.495 195.495 ;
        RECT 90.910 191.690 91.830 220.930 ;
        RECT 94.870 197.630 95.790 220.930 ;
        RECT 97.650 197.120 98.570 198.550 ;
        RECT 100.690 197.120 101.610 198.550 ;
        RECT 103.670 197.630 104.590 220.930 ;
        RECT 107.630 199.070 108.550 220.930 ;
        RECT 115.330 207.900 115.670 221.470 ;
        RECT 113.950 207.560 115.670 207.900 ;
        RECT 113.310 204.040 115.030 204.380 ;
        RECT 82.330 190.440 83.350 191.490 ;
        RECT 81.455 156.930 81.800 157.850 ;
        RECT 81.455 119.830 81.795 156.930 ;
        RECT 82.330 134.070 83.250 190.440 ;
        RECT 90.810 189.240 91.830 191.690 ;
        RECT 84.330 156.780 85.250 157.120 ;
        RECT 88.810 156.780 89.730 157.120 ;
        RECT 90.810 134.070 91.730 189.240 ;
        RECT 92.260 120.760 92.600 196.030 ;
        RECT 97.650 195.620 101.610 197.120 ;
        RECT 109.930 196.770 110.270 197.970 ;
        RECT 106.655 196.430 110.270 196.770 ;
        RECT 94.770 193.360 95.690 194.950 ;
        RECT 97.650 193.360 98.570 195.620 ;
        RECT 100.690 193.360 101.610 195.620 ;
        RECT 94.770 192.440 101.610 193.360 ;
        RECT 92.975 161.330 93.315 162.250 ;
        RECT 93.760 130.060 94.100 166.650 ;
        RECT 94.770 134.070 95.690 192.440 ;
        RECT 97.650 153.700 98.570 192.440 ;
        RECT 100.690 153.700 101.610 192.440 ;
        RECT 102.550 150.985 102.890 196.070 ;
        RECT 102.525 150.595 102.915 150.985 ;
        RECT 103.570 134.070 104.490 194.950 ;
        RECT 105.160 165.730 105.500 166.650 ;
        RECT 105.945 161.330 106.285 162.250 ;
        RECT 106.655 157.850 106.995 196.430 ;
        RECT 111.830 192.170 112.170 199.470 ;
        RECT 113.310 197.970 113.650 204.040 ;
        RECT 116.110 200.860 117.030 221.810 ;
        RECT 116.010 199.070 117.030 200.860 ;
        RECT 113.310 197.630 115.030 197.970 ;
        RECT 114.230 196.730 114.570 197.630 ;
        RECT 111.830 191.830 113.200 192.170 ;
        RECT 106.655 156.930 107.000 157.850 ;
        RECT 107.530 134.070 108.450 191.590 ;
        RECT 112.860 179.145 113.200 191.830 ;
        RECT 112.835 178.755 113.225 179.145 ;
        RECT 114.650 163.820 115.570 164.160 ;
        RECT 109.530 156.780 110.450 157.120 ;
        RECT 113.850 140.940 114.770 141.280 ;
        RECT 113.850 112.520 114.190 140.940 ;
        RECT 115.230 112.520 115.570 163.820 ;
        RECT 116.010 134.070 116.930 199.070 ;
        RECT 120.070 197.630 120.990 221.810 ;
        RECT 134.690 220.930 135.030 222.980 ;
        RECT 132.440 220.590 155.200 220.930 ;
        RECT 130.730 196.095 131.070 215.370 ;
        RECT 130.705 195.705 131.095 196.095 ;
        RECT 119.970 161.960 120.890 194.950 ;
        RECT 140.035 190.650 141.035 206.905 ;
        RECT 143.995 195.590 144.995 206.905 ;
        RECT 147.530 197.095 147.870 198.300 ;
        RECT 147.505 196.705 147.895 197.095 ;
        RECT 143.995 193.795 146.300 195.590 ;
        RECT 144.530 193.790 146.300 193.795 ;
        RECT 144.690 183.500 146.190 193.790 ;
        RECT 134.880 163.100 154.740 181.500 ;
        RECT 119.970 161.620 121.690 161.960 ;
        RECT 119.970 146.120 120.890 161.620 ;
        RECT 121.350 161.520 121.690 161.620 ;
        RECT 121.350 161.180 123.050 161.520 ;
        RECT 119.970 145.780 121.690 146.120 ;
        RECT 119.970 134.070 120.890 145.780 ;
        RECT 121.350 145.680 121.690 145.780 ;
        RECT 121.350 145.340 123.050 145.680 ;
        RECT 134.880 143.500 154.740 161.900 ;
        RECT 134.880 123.900 154.740 142.300 ;
        RECT 55.140 110.820 124.440 111.160 ;
        RECT 55.140 108.960 124.440 109.300 ;
        RECT 55.140 106.510 55.480 107.430 ;
        RECT 12.240 38.170 12.580 106.510 ;
        RECT 12.900 106.170 55.480 106.510 ;
        RECT 12.900 89.510 13.240 106.170 ;
        RECT 13.560 89.830 13.900 105.850 ;
        RECT 14.220 89.510 14.560 106.170 ;
        RECT 14.880 89.830 15.220 105.850 ;
        RECT 15.540 89.510 15.880 106.170 ;
        RECT 16.200 89.830 16.540 105.850 ;
        RECT 16.860 89.510 17.200 106.170 ;
        RECT 17.520 89.830 17.860 105.850 ;
        RECT 18.180 89.510 18.520 106.170 ;
        RECT 18.840 89.830 19.180 105.850 ;
        RECT 19.500 89.510 19.840 106.170 ;
        RECT 20.160 89.830 20.500 105.850 ;
        RECT 20.820 89.510 21.160 106.170 ;
        RECT 21.480 89.830 21.820 105.850 ;
        RECT 22.140 89.510 22.480 106.170 ;
        RECT 22.800 89.830 23.140 105.850 ;
        RECT 23.460 89.510 23.800 106.170 ;
        RECT 24.120 89.830 24.460 105.850 ;
        RECT 24.780 89.510 25.120 106.170 ;
        RECT 25.440 89.830 25.780 105.850 ;
        RECT 26.100 89.510 26.440 106.170 ;
        RECT 26.760 89.830 27.100 105.850 ;
        RECT 27.420 89.510 27.760 106.170 ;
        RECT 28.080 89.830 28.420 105.850 ;
        RECT 28.740 89.510 29.080 106.170 ;
        RECT 29.400 89.830 29.740 105.850 ;
        RECT 30.060 89.510 30.400 106.170 ;
        RECT 30.720 89.830 31.060 105.850 ;
        RECT 31.380 89.510 31.720 106.170 ;
        RECT 32.040 89.830 32.380 105.850 ;
        RECT 32.700 89.510 33.040 106.170 ;
        RECT 33.360 89.830 33.700 105.850 ;
        RECT 34.020 89.510 34.360 106.170 ;
        RECT 34.680 89.830 35.020 105.850 ;
        RECT 35.340 89.510 35.680 106.170 ;
        RECT 36.000 89.830 36.340 105.850 ;
        RECT 36.660 89.510 37.000 106.170 ;
        RECT 37.320 89.830 37.660 105.850 ;
        RECT 37.980 89.510 38.320 106.170 ;
        RECT 38.640 89.830 38.980 105.850 ;
        RECT 39.300 89.510 39.640 106.170 ;
        RECT 39.960 89.830 40.300 105.850 ;
        RECT 40.620 89.510 40.960 106.170 ;
        RECT 41.280 89.830 41.620 105.850 ;
        RECT 41.940 89.510 42.280 106.170 ;
        RECT 42.600 89.830 42.940 105.850 ;
        RECT 43.260 89.510 43.600 106.170 ;
        RECT 43.920 89.830 44.260 105.850 ;
        RECT 44.580 89.510 44.920 106.170 ;
        RECT 45.240 89.830 45.580 105.850 ;
        RECT 45.900 89.510 46.240 106.170 ;
        RECT 46.560 89.830 46.900 105.850 ;
        RECT 47.220 89.510 47.560 106.170 ;
        RECT 47.880 89.830 48.220 105.850 ;
        RECT 48.540 89.510 48.880 106.170 ;
        RECT 49.200 89.830 49.540 105.850 ;
        RECT 49.860 89.510 50.200 106.170 ;
        RECT 50.520 89.830 50.860 105.850 ;
        RECT 51.180 89.510 51.520 106.170 ;
        RECT 51.840 89.830 52.180 105.850 ;
        RECT 52.500 89.510 52.840 106.170 ;
        RECT 53.160 89.830 53.500 105.850 ;
        RECT 53.820 89.510 54.160 106.170 ;
        RECT 54.480 89.830 54.820 105.850 ;
        RECT 55.140 89.510 55.480 106.170 ;
        RECT 12.900 89.170 55.480 89.510 ;
        RECT 12.900 72.510 13.240 89.170 ;
        RECT 13.560 72.830 13.900 88.850 ;
        RECT 14.220 72.510 14.560 89.170 ;
        RECT 14.880 72.830 15.220 88.850 ;
        RECT 15.540 72.510 15.880 89.170 ;
        RECT 16.200 72.830 16.540 88.850 ;
        RECT 16.860 72.510 17.200 89.170 ;
        RECT 17.520 72.830 17.860 88.850 ;
        RECT 18.180 72.510 18.520 89.170 ;
        RECT 18.840 72.830 19.180 88.850 ;
        RECT 19.500 72.510 19.840 89.170 ;
        RECT 20.160 72.830 20.500 88.850 ;
        RECT 20.820 72.510 21.160 89.170 ;
        RECT 21.480 72.830 21.820 88.850 ;
        RECT 22.140 72.510 22.480 89.170 ;
        RECT 22.800 72.830 23.140 88.850 ;
        RECT 23.460 72.510 23.800 89.170 ;
        RECT 24.120 72.830 24.460 88.850 ;
        RECT 24.780 72.510 25.120 89.170 ;
        RECT 25.440 72.830 25.780 88.850 ;
        RECT 26.100 72.510 26.440 89.170 ;
        RECT 26.760 72.830 27.100 88.850 ;
        RECT 27.420 72.510 27.760 89.170 ;
        RECT 28.080 72.830 28.420 88.850 ;
        RECT 28.740 72.510 29.080 89.170 ;
        RECT 29.400 72.830 29.740 88.850 ;
        RECT 30.060 72.510 30.400 89.170 ;
        RECT 30.720 72.830 31.060 88.850 ;
        RECT 31.380 72.510 31.720 89.170 ;
        RECT 32.040 72.830 32.380 88.850 ;
        RECT 32.700 72.510 33.040 89.170 ;
        RECT 33.360 72.830 33.700 88.850 ;
        RECT 34.020 72.510 34.360 89.170 ;
        RECT 34.680 72.830 35.020 88.850 ;
        RECT 35.340 72.510 35.680 89.170 ;
        RECT 36.000 72.830 36.340 88.850 ;
        RECT 36.660 72.510 37.000 89.170 ;
        RECT 37.320 72.830 37.660 88.850 ;
        RECT 37.980 72.510 38.320 89.170 ;
        RECT 38.640 72.830 38.980 88.850 ;
        RECT 39.300 72.510 39.640 89.170 ;
        RECT 39.960 72.830 40.300 88.850 ;
        RECT 40.620 72.510 40.960 89.170 ;
        RECT 41.280 72.830 41.620 88.850 ;
        RECT 41.940 72.510 42.280 89.170 ;
        RECT 42.600 72.830 42.940 88.850 ;
        RECT 43.260 72.510 43.600 89.170 ;
        RECT 43.920 72.830 44.260 88.850 ;
        RECT 44.580 72.510 44.920 89.170 ;
        RECT 45.240 72.830 45.580 88.850 ;
        RECT 45.900 72.510 46.240 89.170 ;
        RECT 46.560 72.830 46.900 88.850 ;
        RECT 47.220 72.510 47.560 89.170 ;
        RECT 47.880 72.830 48.220 88.850 ;
        RECT 48.540 72.510 48.880 89.170 ;
        RECT 49.200 72.830 49.540 88.850 ;
        RECT 49.860 72.510 50.200 89.170 ;
        RECT 50.520 72.830 50.860 88.850 ;
        RECT 51.180 72.510 51.520 89.170 ;
        RECT 51.840 72.830 52.180 88.850 ;
        RECT 52.500 72.510 52.840 89.170 ;
        RECT 53.160 72.830 53.500 88.850 ;
        RECT 53.820 72.510 54.160 89.170 ;
        RECT 54.480 72.830 54.820 88.850 ;
        RECT 55.140 72.510 55.480 89.170 ;
        RECT 12.900 72.170 55.480 72.510 ;
        RECT 12.900 55.510 13.240 72.170 ;
        RECT 13.560 55.830 13.900 71.850 ;
        RECT 14.220 55.510 14.560 72.170 ;
        RECT 14.880 55.830 15.220 71.850 ;
        RECT 15.540 55.510 15.880 72.170 ;
        RECT 16.200 55.830 16.540 71.850 ;
        RECT 16.860 55.510 17.200 72.170 ;
        RECT 17.520 55.830 17.860 71.850 ;
        RECT 18.180 55.510 18.520 72.170 ;
        RECT 18.840 55.830 19.180 71.850 ;
        RECT 19.500 55.510 19.840 72.170 ;
        RECT 20.160 55.830 20.500 71.850 ;
        RECT 20.820 55.510 21.160 72.170 ;
        RECT 21.480 55.830 21.820 71.850 ;
        RECT 22.140 55.510 22.480 72.170 ;
        RECT 22.800 55.830 23.140 71.850 ;
        RECT 23.460 55.510 23.800 72.170 ;
        RECT 24.120 55.830 24.460 71.850 ;
        RECT 24.780 55.510 25.120 72.170 ;
        RECT 25.440 55.830 25.780 71.850 ;
        RECT 26.100 55.510 26.440 72.170 ;
        RECT 26.760 55.830 27.100 71.850 ;
        RECT 27.420 55.510 27.760 72.170 ;
        RECT 28.080 55.830 28.420 71.850 ;
        RECT 28.740 55.510 29.080 72.170 ;
        RECT 29.400 55.830 29.740 71.850 ;
        RECT 30.060 55.510 30.400 72.170 ;
        RECT 30.720 55.830 31.060 71.850 ;
        RECT 31.380 55.510 31.720 72.170 ;
        RECT 32.040 55.830 32.380 71.850 ;
        RECT 32.700 55.510 33.040 72.170 ;
        RECT 33.360 55.830 33.700 71.850 ;
        RECT 34.020 55.510 34.360 72.170 ;
        RECT 34.680 55.830 35.020 71.850 ;
        RECT 35.340 55.510 35.680 72.170 ;
        RECT 36.000 55.830 36.340 71.850 ;
        RECT 36.660 55.510 37.000 72.170 ;
        RECT 37.320 55.830 37.660 71.850 ;
        RECT 37.980 55.510 38.320 72.170 ;
        RECT 38.640 55.830 38.980 71.850 ;
        RECT 39.300 55.510 39.640 72.170 ;
        RECT 39.960 55.830 40.300 71.850 ;
        RECT 40.620 55.510 40.960 72.170 ;
        RECT 41.280 55.830 41.620 71.850 ;
        RECT 41.940 55.510 42.280 72.170 ;
        RECT 42.600 55.830 42.940 71.850 ;
        RECT 43.260 55.510 43.600 72.170 ;
        RECT 43.920 55.830 44.260 71.850 ;
        RECT 44.580 55.510 44.920 72.170 ;
        RECT 45.240 55.830 45.580 71.850 ;
        RECT 45.900 55.510 46.240 72.170 ;
        RECT 46.560 55.830 46.900 71.850 ;
        RECT 47.220 55.510 47.560 72.170 ;
        RECT 47.880 55.830 48.220 71.850 ;
        RECT 48.540 55.510 48.880 72.170 ;
        RECT 49.200 55.830 49.540 71.850 ;
        RECT 49.860 55.510 50.200 72.170 ;
        RECT 50.520 55.830 50.860 71.850 ;
        RECT 51.180 55.510 51.520 72.170 ;
        RECT 51.840 55.830 52.180 71.850 ;
        RECT 52.500 55.510 52.840 72.170 ;
        RECT 53.160 55.830 53.500 71.850 ;
        RECT 53.820 55.510 54.160 72.170 ;
        RECT 54.480 55.830 54.820 71.850 ;
        RECT 55.140 55.510 55.480 72.170 ;
        RECT 12.900 55.170 55.480 55.510 ;
        RECT 12.900 38.510 13.240 55.170 ;
        RECT 13.560 38.830 13.900 54.850 ;
        RECT 14.220 38.510 14.560 55.170 ;
        RECT 14.880 38.830 15.220 54.850 ;
        RECT 15.540 38.510 15.880 55.170 ;
        RECT 16.200 38.830 16.540 54.850 ;
        RECT 16.860 38.510 17.200 55.170 ;
        RECT 17.520 38.830 17.860 54.850 ;
        RECT 18.180 38.510 18.520 55.170 ;
        RECT 18.840 38.830 19.180 54.850 ;
        RECT 19.500 38.510 19.840 55.170 ;
        RECT 20.160 38.830 20.500 54.850 ;
        RECT 20.820 38.510 21.160 55.170 ;
        RECT 21.480 38.830 21.820 54.850 ;
        RECT 22.140 38.510 22.480 55.170 ;
        RECT 22.800 38.830 23.140 54.850 ;
        RECT 23.460 38.510 23.800 55.170 ;
        RECT 24.120 38.830 24.460 54.850 ;
        RECT 24.780 38.510 25.120 55.170 ;
        RECT 25.440 38.830 25.780 54.850 ;
        RECT 26.100 38.510 26.440 55.170 ;
        RECT 26.760 38.830 27.100 54.850 ;
        RECT 27.420 38.510 27.760 55.170 ;
        RECT 28.080 38.830 28.420 54.850 ;
        RECT 28.740 38.510 29.080 55.170 ;
        RECT 29.400 38.830 29.740 54.850 ;
        RECT 30.060 38.510 30.400 55.170 ;
        RECT 30.720 38.830 31.060 54.850 ;
        RECT 31.380 38.510 31.720 55.170 ;
        RECT 32.040 38.830 32.380 54.850 ;
        RECT 32.700 38.510 33.040 55.170 ;
        RECT 33.360 38.830 33.700 54.850 ;
        RECT 34.020 38.510 34.360 55.170 ;
        RECT 34.680 38.830 35.020 54.850 ;
        RECT 35.340 38.510 35.680 55.170 ;
        RECT 36.000 38.830 36.340 54.850 ;
        RECT 36.660 38.510 37.000 55.170 ;
        RECT 37.320 38.830 37.660 54.850 ;
        RECT 37.980 38.510 38.320 55.170 ;
        RECT 38.640 38.830 38.980 54.850 ;
        RECT 39.300 38.510 39.640 55.170 ;
        RECT 39.960 38.830 40.300 54.850 ;
        RECT 40.620 38.510 40.960 55.170 ;
        RECT 41.280 38.830 41.620 54.850 ;
        RECT 41.940 38.510 42.280 55.170 ;
        RECT 42.600 38.830 42.940 54.850 ;
        RECT 43.260 38.510 43.600 55.170 ;
        RECT 43.920 38.830 44.260 54.850 ;
        RECT 44.580 38.510 44.920 55.170 ;
        RECT 45.240 38.830 45.580 54.850 ;
        RECT 45.900 38.510 46.240 55.170 ;
        RECT 46.560 38.830 46.900 54.850 ;
        RECT 47.220 38.510 47.560 55.170 ;
        RECT 47.880 38.830 48.220 54.850 ;
        RECT 48.540 38.510 48.880 55.170 ;
        RECT 49.200 38.830 49.540 54.850 ;
        RECT 49.860 38.510 50.200 55.170 ;
        RECT 50.520 38.830 50.860 54.850 ;
        RECT 51.180 38.510 51.520 55.170 ;
        RECT 51.840 38.830 52.180 54.850 ;
        RECT 52.500 38.510 52.840 55.170 ;
        RECT 53.160 38.830 53.500 54.850 ;
        RECT 53.820 38.510 54.160 55.170 ;
        RECT 54.480 38.830 54.820 54.850 ;
        RECT 55.140 38.510 55.480 55.170 ;
        RECT 80.780 106.510 81.120 107.430 ;
        RECT 80.780 106.170 123.360 106.510 ;
        RECT 80.780 89.510 81.120 106.170 ;
        RECT 81.440 89.830 81.780 105.850 ;
        RECT 82.100 89.510 82.440 106.170 ;
        RECT 82.760 89.830 83.100 105.850 ;
        RECT 83.420 89.510 83.760 106.170 ;
        RECT 84.080 89.830 84.420 105.850 ;
        RECT 84.740 89.510 85.080 106.170 ;
        RECT 85.400 89.830 85.740 105.850 ;
        RECT 86.060 89.510 86.400 106.170 ;
        RECT 86.720 89.830 87.060 105.850 ;
        RECT 87.380 89.510 87.720 106.170 ;
        RECT 88.040 89.830 88.380 105.850 ;
        RECT 88.700 89.510 89.040 106.170 ;
        RECT 89.360 89.830 89.700 105.850 ;
        RECT 90.020 89.510 90.360 106.170 ;
        RECT 90.680 89.830 91.020 105.850 ;
        RECT 91.340 89.510 91.680 106.170 ;
        RECT 92.000 89.830 92.340 105.850 ;
        RECT 92.660 89.510 93.000 106.170 ;
        RECT 93.320 89.830 93.660 105.850 ;
        RECT 93.980 89.510 94.320 106.170 ;
        RECT 94.640 89.830 94.980 105.850 ;
        RECT 95.300 89.510 95.640 106.170 ;
        RECT 95.960 89.830 96.300 105.850 ;
        RECT 96.620 89.510 96.960 106.170 ;
        RECT 97.280 89.830 97.620 105.850 ;
        RECT 97.940 89.510 98.280 106.170 ;
        RECT 98.600 89.830 98.940 105.850 ;
        RECT 99.260 89.510 99.600 106.170 ;
        RECT 99.920 89.830 100.260 105.850 ;
        RECT 100.580 89.510 100.920 106.170 ;
        RECT 101.240 89.830 101.580 105.850 ;
        RECT 101.900 89.510 102.240 106.170 ;
        RECT 102.560 89.830 102.900 105.850 ;
        RECT 103.220 89.510 103.560 106.170 ;
        RECT 103.880 89.830 104.220 105.850 ;
        RECT 104.540 89.510 104.880 106.170 ;
        RECT 105.200 89.830 105.540 105.850 ;
        RECT 105.860 89.510 106.200 106.170 ;
        RECT 106.520 89.830 106.860 105.850 ;
        RECT 107.180 89.510 107.520 106.170 ;
        RECT 107.840 89.830 108.180 105.850 ;
        RECT 108.500 89.510 108.840 106.170 ;
        RECT 109.160 89.830 109.500 105.850 ;
        RECT 109.820 89.510 110.160 106.170 ;
        RECT 110.480 89.830 110.820 105.850 ;
        RECT 111.140 89.510 111.480 106.170 ;
        RECT 111.800 89.830 112.140 105.850 ;
        RECT 112.460 89.510 112.800 106.170 ;
        RECT 113.120 89.830 113.460 105.850 ;
        RECT 113.780 89.510 114.120 106.170 ;
        RECT 114.440 89.830 114.780 105.850 ;
        RECT 115.100 89.510 115.440 106.170 ;
        RECT 115.760 89.830 116.100 105.850 ;
        RECT 116.420 89.510 116.760 106.170 ;
        RECT 117.080 89.830 117.420 105.850 ;
        RECT 117.740 89.510 118.080 106.170 ;
        RECT 118.400 89.830 118.740 105.850 ;
        RECT 119.060 89.510 119.400 106.170 ;
        RECT 119.720 89.830 120.060 105.850 ;
        RECT 120.380 89.510 120.720 106.170 ;
        RECT 121.040 89.830 121.380 105.850 ;
        RECT 121.700 89.510 122.040 106.170 ;
        RECT 122.360 89.830 122.700 105.850 ;
        RECT 123.020 89.510 123.360 106.170 ;
        RECT 80.780 89.170 123.360 89.510 ;
        RECT 80.780 72.510 81.120 89.170 ;
        RECT 81.440 72.830 81.780 88.850 ;
        RECT 82.100 72.510 82.440 89.170 ;
        RECT 82.760 72.830 83.100 88.850 ;
        RECT 83.420 72.510 83.760 89.170 ;
        RECT 84.080 72.830 84.420 88.850 ;
        RECT 84.740 72.510 85.080 89.170 ;
        RECT 85.400 72.830 85.740 88.850 ;
        RECT 86.060 72.510 86.400 89.170 ;
        RECT 86.720 72.830 87.060 88.850 ;
        RECT 87.380 72.510 87.720 89.170 ;
        RECT 88.040 72.830 88.380 88.850 ;
        RECT 88.700 72.510 89.040 89.170 ;
        RECT 89.360 72.830 89.700 88.850 ;
        RECT 90.020 72.510 90.360 89.170 ;
        RECT 90.680 72.830 91.020 88.850 ;
        RECT 91.340 72.510 91.680 89.170 ;
        RECT 92.000 72.830 92.340 88.850 ;
        RECT 92.660 72.510 93.000 89.170 ;
        RECT 93.320 72.830 93.660 88.850 ;
        RECT 93.980 72.510 94.320 89.170 ;
        RECT 94.640 72.830 94.980 88.850 ;
        RECT 95.300 72.510 95.640 89.170 ;
        RECT 95.960 72.830 96.300 88.850 ;
        RECT 96.620 72.510 96.960 89.170 ;
        RECT 97.280 72.830 97.620 88.850 ;
        RECT 97.940 72.510 98.280 89.170 ;
        RECT 98.600 72.830 98.940 88.850 ;
        RECT 99.260 72.510 99.600 89.170 ;
        RECT 99.920 72.830 100.260 88.850 ;
        RECT 100.580 72.510 100.920 89.170 ;
        RECT 101.240 72.830 101.580 88.850 ;
        RECT 101.900 72.510 102.240 89.170 ;
        RECT 102.560 72.830 102.900 88.850 ;
        RECT 103.220 72.510 103.560 89.170 ;
        RECT 103.880 72.830 104.220 88.850 ;
        RECT 104.540 72.510 104.880 89.170 ;
        RECT 105.200 72.830 105.540 88.850 ;
        RECT 105.860 72.510 106.200 89.170 ;
        RECT 106.520 72.830 106.860 88.850 ;
        RECT 107.180 72.510 107.520 89.170 ;
        RECT 107.840 72.830 108.180 88.850 ;
        RECT 108.500 72.510 108.840 89.170 ;
        RECT 109.160 72.830 109.500 88.850 ;
        RECT 109.820 72.510 110.160 89.170 ;
        RECT 110.480 72.830 110.820 88.850 ;
        RECT 111.140 72.510 111.480 89.170 ;
        RECT 111.800 72.830 112.140 88.850 ;
        RECT 112.460 72.510 112.800 89.170 ;
        RECT 113.120 72.830 113.460 88.850 ;
        RECT 113.780 72.510 114.120 89.170 ;
        RECT 114.440 72.830 114.780 88.850 ;
        RECT 115.100 72.510 115.440 89.170 ;
        RECT 115.760 72.830 116.100 88.850 ;
        RECT 116.420 72.510 116.760 89.170 ;
        RECT 117.080 72.830 117.420 88.850 ;
        RECT 117.740 72.510 118.080 89.170 ;
        RECT 118.400 72.830 118.740 88.850 ;
        RECT 119.060 72.510 119.400 89.170 ;
        RECT 119.720 72.830 120.060 88.850 ;
        RECT 120.380 72.510 120.720 89.170 ;
        RECT 121.040 72.830 121.380 88.850 ;
        RECT 121.700 72.510 122.040 89.170 ;
        RECT 122.360 72.830 122.700 88.850 ;
        RECT 123.020 72.510 123.360 89.170 ;
        RECT 80.780 72.170 123.360 72.510 ;
        RECT 80.780 55.510 81.120 72.170 ;
        RECT 81.440 55.830 81.780 71.850 ;
        RECT 82.100 55.510 82.440 72.170 ;
        RECT 82.760 55.830 83.100 71.850 ;
        RECT 83.420 55.510 83.760 72.170 ;
        RECT 84.080 55.830 84.420 71.850 ;
        RECT 84.740 55.510 85.080 72.170 ;
        RECT 85.400 55.830 85.740 71.850 ;
        RECT 86.060 55.510 86.400 72.170 ;
        RECT 86.720 55.830 87.060 71.850 ;
        RECT 87.380 55.510 87.720 72.170 ;
        RECT 88.040 55.830 88.380 71.850 ;
        RECT 88.700 55.510 89.040 72.170 ;
        RECT 89.360 55.830 89.700 71.850 ;
        RECT 90.020 55.510 90.360 72.170 ;
        RECT 90.680 55.830 91.020 71.850 ;
        RECT 91.340 55.510 91.680 72.170 ;
        RECT 92.000 55.830 92.340 71.850 ;
        RECT 92.660 55.510 93.000 72.170 ;
        RECT 93.320 55.830 93.660 71.850 ;
        RECT 93.980 55.510 94.320 72.170 ;
        RECT 94.640 55.830 94.980 71.850 ;
        RECT 95.300 55.510 95.640 72.170 ;
        RECT 95.960 55.830 96.300 71.850 ;
        RECT 96.620 55.510 96.960 72.170 ;
        RECT 97.280 55.830 97.620 71.850 ;
        RECT 97.940 55.510 98.280 72.170 ;
        RECT 98.600 55.830 98.940 71.850 ;
        RECT 99.260 55.510 99.600 72.170 ;
        RECT 99.920 55.830 100.260 71.850 ;
        RECT 100.580 55.510 100.920 72.170 ;
        RECT 101.240 55.830 101.580 71.850 ;
        RECT 101.900 55.510 102.240 72.170 ;
        RECT 102.560 55.830 102.900 71.850 ;
        RECT 103.220 55.510 103.560 72.170 ;
        RECT 103.880 55.830 104.220 71.850 ;
        RECT 104.540 55.510 104.880 72.170 ;
        RECT 105.200 55.830 105.540 71.850 ;
        RECT 105.860 55.510 106.200 72.170 ;
        RECT 106.520 55.830 106.860 71.850 ;
        RECT 107.180 55.510 107.520 72.170 ;
        RECT 107.840 55.830 108.180 71.850 ;
        RECT 108.500 55.510 108.840 72.170 ;
        RECT 109.160 55.830 109.500 71.850 ;
        RECT 109.820 55.510 110.160 72.170 ;
        RECT 110.480 55.830 110.820 71.850 ;
        RECT 111.140 55.510 111.480 72.170 ;
        RECT 111.800 55.830 112.140 71.850 ;
        RECT 112.460 55.510 112.800 72.170 ;
        RECT 113.120 55.830 113.460 71.850 ;
        RECT 113.780 55.510 114.120 72.170 ;
        RECT 114.440 55.830 114.780 71.850 ;
        RECT 115.100 55.510 115.440 72.170 ;
        RECT 115.760 55.830 116.100 71.850 ;
        RECT 116.420 55.510 116.760 72.170 ;
        RECT 117.080 55.830 117.420 71.850 ;
        RECT 117.740 55.510 118.080 72.170 ;
        RECT 118.400 55.830 118.740 71.850 ;
        RECT 119.060 55.510 119.400 72.170 ;
        RECT 119.720 55.830 120.060 71.850 ;
        RECT 120.380 55.510 120.720 72.170 ;
        RECT 121.040 55.830 121.380 71.850 ;
        RECT 121.700 55.510 122.040 72.170 ;
        RECT 122.360 55.830 122.700 71.850 ;
        RECT 123.020 55.510 123.360 72.170 ;
        RECT 80.780 55.170 123.360 55.510 ;
        RECT 80.780 38.510 81.120 55.170 ;
        RECT 81.440 38.830 81.780 54.850 ;
        RECT 82.100 38.510 82.440 55.170 ;
        RECT 82.760 38.830 83.100 54.850 ;
        RECT 83.420 38.510 83.760 55.170 ;
        RECT 84.080 38.830 84.420 54.850 ;
        RECT 84.740 38.510 85.080 55.170 ;
        RECT 85.400 38.830 85.740 54.850 ;
        RECT 86.060 38.510 86.400 55.170 ;
        RECT 86.720 38.830 87.060 54.850 ;
        RECT 87.380 38.510 87.720 55.170 ;
        RECT 88.040 38.830 88.380 54.850 ;
        RECT 88.700 38.510 89.040 55.170 ;
        RECT 89.360 38.830 89.700 54.850 ;
        RECT 90.020 38.510 90.360 55.170 ;
        RECT 90.680 38.830 91.020 54.850 ;
        RECT 91.340 38.510 91.680 55.170 ;
        RECT 92.000 38.830 92.340 54.850 ;
        RECT 92.660 38.510 93.000 55.170 ;
        RECT 93.320 38.830 93.660 54.850 ;
        RECT 93.980 38.510 94.320 55.170 ;
        RECT 94.640 38.830 94.980 54.850 ;
        RECT 95.300 38.510 95.640 55.170 ;
        RECT 95.960 38.830 96.300 54.850 ;
        RECT 96.620 38.510 96.960 55.170 ;
        RECT 97.280 38.830 97.620 54.850 ;
        RECT 97.940 38.510 98.280 55.170 ;
        RECT 98.600 38.830 98.940 54.850 ;
        RECT 99.260 38.510 99.600 55.170 ;
        RECT 99.920 38.830 100.260 54.850 ;
        RECT 100.580 38.510 100.920 55.170 ;
        RECT 101.240 38.830 101.580 54.850 ;
        RECT 101.900 38.510 102.240 55.170 ;
        RECT 102.560 38.830 102.900 54.850 ;
        RECT 103.220 38.510 103.560 55.170 ;
        RECT 103.880 38.830 104.220 54.850 ;
        RECT 104.540 38.510 104.880 55.170 ;
        RECT 105.200 38.830 105.540 54.850 ;
        RECT 105.860 38.510 106.200 55.170 ;
        RECT 106.520 38.830 106.860 54.850 ;
        RECT 107.180 38.510 107.520 55.170 ;
        RECT 107.840 38.830 108.180 54.850 ;
        RECT 108.500 38.510 108.840 55.170 ;
        RECT 109.160 38.830 109.500 54.850 ;
        RECT 109.820 38.510 110.160 55.170 ;
        RECT 110.480 38.830 110.820 54.850 ;
        RECT 111.140 38.510 111.480 55.170 ;
        RECT 111.800 38.830 112.140 54.850 ;
        RECT 112.460 38.510 112.800 55.170 ;
        RECT 113.120 38.830 113.460 54.850 ;
        RECT 113.780 38.510 114.120 55.170 ;
        RECT 114.440 38.830 114.780 54.850 ;
        RECT 115.100 38.510 115.440 55.170 ;
        RECT 115.760 38.830 116.100 54.850 ;
        RECT 116.420 38.510 116.760 55.170 ;
        RECT 117.080 38.830 117.420 54.850 ;
        RECT 117.740 38.510 118.080 55.170 ;
        RECT 118.400 38.830 118.740 54.850 ;
        RECT 119.060 38.510 119.400 55.170 ;
        RECT 119.720 38.830 120.060 54.850 ;
        RECT 120.380 38.510 120.720 55.170 ;
        RECT 121.040 38.830 121.380 54.850 ;
        RECT 121.700 38.510 122.040 55.170 ;
        RECT 122.360 38.830 122.700 54.850 ;
        RECT 123.020 38.510 123.360 55.170 ;
        RECT 12.900 38.170 62.970 38.510 ;
        RECT 11.070 36.580 46.710 36.640 ;
        RECT 11.070 36.240 47.350 36.580 ;
        RECT 11.070 35.440 45.990 35.840 ;
        RECT 11.070 34.240 11.430 35.440 ;
        RECT 46.350 35.040 46.710 36.240 ;
        RECT 11.790 34.640 46.710 35.040 ;
        RECT 11.070 33.840 45.270 34.240 ;
        RECT 45.630 33.840 45.990 34.240 ;
        RECT 11.070 32.640 11.430 33.840 ;
        RECT 46.350 33.440 46.710 34.640 ;
        RECT 11.790 33.040 12.510 33.440 ;
        RECT 12.870 33.040 46.710 33.440 ;
        RECT 11.070 32.580 46.710 32.640 ;
        RECT 10.430 32.240 46.710 32.580 ;
        RECT 10.430 27.780 10.770 32.240 ;
        RECT 11.070 31.780 46.710 31.840 ;
        RECT 47.010 31.780 47.350 36.240 ;
        RECT 11.070 31.440 47.350 31.780 ;
        RECT 11.070 30.640 45.990 31.040 ;
        RECT 11.070 29.440 11.430 30.640 ;
        RECT 46.350 30.240 46.710 31.440 ;
        RECT 11.790 29.840 46.710 30.240 ;
        RECT 11.070 29.040 45.270 29.440 ;
        RECT 45.630 29.040 45.990 29.440 ;
        RECT 11.070 27.840 11.430 29.040 ;
        RECT 46.350 28.640 46.710 29.840 ;
        RECT 11.790 28.240 12.510 28.640 ;
        RECT 12.870 28.240 46.710 28.640 ;
        RECT 11.070 27.780 46.710 27.840 ;
        RECT 10.430 27.440 46.710 27.780 ;
        RECT 10.430 22.980 10.770 27.440 ;
        RECT 11.070 26.980 46.710 27.040 ;
        RECT 47.010 26.980 47.350 31.440 ;
        RECT 11.070 26.640 47.350 26.980 ;
        RECT 11.070 25.840 45.990 26.240 ;
        RECT 11.070 24.640 11.430 25.840 ;
        RECT 46.350 25.440 46.710 26.640 ;
        RECT 11.790 25.040 46.710 25.440 ;
        RECT 11.070 24.240 45.270 24.640 ;
        RECT 45.630 24.240 45.990 24.640 ;
        RECT 11.070 23.040 11.430 24.240 ;
        RECT 46.350 23.840 46.710 25.040 ;
        RECT 11.790 23.440 12.510 23.840 ;
        RECT 12.870 23.440 46.710 23.840 ;
        RECT 11.070 22.980 46.710 23.040 ;
        RECT 10.430 22.640 46.710 22.980 ;
        RECT 10.430 18.180 10.770 22.640 ;
        RECT 11.070 22.180 46.710 22.240 ;
        RECT 47.010 22.180 47.350 26.640 ;
        RECT 11.070 21.840 47.350 22.180 ;
        RECT 11.070 21.040 45.990 21.440 ;
        RECT 11.070 19.840 11.430 21.040 ;
        RECT 46.350 20.640 46.710 21.840 ;
        RECT 11.790 20.240 46.710 20.640 ;
        RECT 11.070 19.440 45.270 19.840 ;
        RECT 45.630 19.440 45.990 19.840 ;
        RECT 11.070 18.240 11.430 19.440 ;
        RECT 46.350 19.040 46.710 20.240 ;
        RECT 11.790 18.640 12.510 19.040 ;
        RECT 12.870 18.640 46.710 19.040 ;
        RECT 47.010 21.770 47.350 21.840 ;
        RECT 47.010 21.430 51.030 21.770 ;
        RECT 11.070 18.180 46.710 18.240 ;
        RECT 10.430 17.840 46.710 18.180 ;
        RECT 10.430 13.380 10.770 17.840 ;
        RECT 11.070 17.380 46.710 17.440 ;
        RECT 47.010 17.380 47.350 21.430 ;
        RECT 50.110 18.350 51.810 18.690 ;
        RECT 51.470 18.250 51.810 18.350 ;
        RECT 52.270 18.250 53.190 37.240 ;
        RECT 51.470 17.910 53.190 18.250 ;
        RECT 11.070 17.040 47.350 17.380 ;
        RECT 11.070 16.240 45.990 16.640 ;
        RECT 11.070 15.040 11.430 16.240 ;
        RECT 46.350 15.840 46.710 17.040 ;
        RECT 11.790 15.440 46.710 15.840 ;
        RECT 11.070 14.640 45.270 15.040 ;
        RECT 45.630 14.640 45.990 15.040 ;
        RECT 11.070 13.440 11.430 14.640 ;
        RECT 46.350 14.240 46.710 15.440 ;
        RECT 11.790 13.840 12.510 14.240 ;
        RECT 12.870 13.840 46.710 14.240 ;
        RECT 11.070 13.380 46.710 13.440 ;
        RECT 10.430 13.040 46.710 13.380 ;
        RECT 52.270 6.040 53.190 17.910 ;
        RECT 56.230 9.640 57.150 37.240 ;
        RECT 58.830 27.590 59.750 27.930 ;
        RECT 59.120 4.260 59.460 27.590 ;
        RECT 62.630 19.130 62.970 38.170 ;
        RECT 73.290 38.170 123.360 38.510 ;
        RECT 123.680 38.170 124.020 106.510 ;
        RECT 134.880 104.300 154.740 122.700 ;
        RECT 134.880 84.700 154.740 103.100 ;
        RECT 134.880 65.100 154.740 83.500 ;
        RECT 134.880 45.500 154.740 63.900 ;
        RECT 64.650 25.830 72.830 26.170 ;
        RECT 64.650 19.130 64.990 25.830 ;
        RECT 73.290 19.130 73.630 38.170 ;
        RECT 76.510 27.590 77.430 27.930 ;
        RECT 62.630 18.790 64.990 19.130 ;
        RECT 71.910 18.790 73.630 19.130 ;
        RECT 63.270 14.390 64.190 14.730 ;
        RECT 72.070 14.390 72.990 14.730 ;
        RECT 76.800 4.260 77.140 27.590 ;
        RECT 79.110 9.640 80.030 37.240 ;
        RECT 83.070 18.250 83.990 37.240 ;
        RECT 89.550 36.580 125.190 36.640 ;
        RECT 88.910 36.240 125.190 36.580 ;
        RECT 88.910 31.780 89.250 36.240 ;
        RECT 89.550 35.040 89.910 36.240 ;
        RECT 90.270 35.440 125.190 35.840 ;
        RECT 89.550 34.640 124.470 35.040 ;
        RECT 89.550 33.440 89.910 34.640 ;
        RECT 124.830 34.240 125.190 35.440 ;
        RECT 90.270 33.840 90.630 34.240 ;
        RECT 90.990 33.840 125.190 34.240 ;
        RECT 89.550 33.040 123.390 33.440 ;
        RECT 123.750 33.040 124.470 33.440 ;
        RECT 124.830 32.640 125.190 33.840 ;
        RECT 89.550 32.580 125.190 32.640 ;
        RECT 89.550 32.240 125.830 32.580 ;
        RECT 89.550 31.780 125.190 31.840 ;
        RECT 88.910 31.440 125.190 31.780 ;
        RECT 88.910 26.980 89.250 31.440 ;
        RECT 89.550 30.240 89.910 31.440 ;
        RECT 90.270 30.640 125.190 31.040 ;
        RECT 89.550 29.840 124.470 30.240 ;
        RECT 89.550 28.640 89.910 29.840 ;
        RECT 124.830 29.440 125.190 30.640 ;
        RECT 90.270 29.040 90.630 29.440 ;
        RECT 90.990 29.040 125.190 29.440 ;
        RECT 89.550 28.240 123.390 28.640 ;
        RECT 123.750 28.240 124.470 28.640 ;
        RECT 124.830 27.840 125.190 29.040 ;
        RECT 89.550 27.780 125.190 27.840 ;
        RECT 125.490 27.780 125.830 32.240 ;
        RECT 89.550 27.440 125.830 27.780 ;
        RECT 89.550 26.980 125.190 27.040 ;
        RECT 88.910 26.640 125.190 26.980 ;
        RECT 88.910 22.180 89.250 26.640 ;
        RECT 89.550 25.440 89.910 26.640 ;
        RECT 90.270 25.840 125.190 26.240 ;
        RECT 89.550 25.040 124.470 25.440 ;
        RECT 89.550 23.840 89.910 25.040 ;
        RECT 124.830 24.640 125.190 25.840 ;
        RECT 90.270 24.240 90.630 24.640 ;
        RECT 90.990 24.240 125.190 24.640 ;
        RECT 89.550 23.440 123.390 23.840 ;
        RECT 123.750 23.440 124.470 23.840 ;
        RECT 124.830 23.040 125.190 24.240 ;
        RECT 89.550 22.980 125.190 23.040 ;
        RECT 125.490 22.980 125.830 27.440 ;
        RECT 134.880 25.900 154.740 44.300 ;
        RECT 89.550 22.640 125.830 22.980 ;
        RECT 89.550 22.180 125.190 22.240 ;
        RECT 88.910 21.840 125.190 22.180 ;
        RECT 88.910 21.770 89.250 21.840 ;
        RECT 85.230 21.430 89.250 21.770 ;
        RECT 84.450 18.350 86.150 18.690 ;
        RECT 84.450 18.250 84.790 18.350 ;
        RECT 83.070 17.910 84.790 18.250 ;
        RECT 83.070 6.040 83.990 17.910 ;
        RECT 88.910 17.380 89.250 21.430 ;
        RECT 89.550 20.640 89.910 21.840 ;
        RECT 90.270 21.040 125.190 21.440 ;
        RECT 89.550 20.240 124.470 20.640 ;
        RECT 89.550 19.040 89.910 20.240 ;
        RECT 124.830 19.840 125.190 21.040 ;
        RECT 90.270 19.440 90.630 19.840 ;
        RECT 90.990 19.440 125.190 19.840 ;
        RECT 89.550 18.640 123.390 19.040 ;
        RECT 123.750 18.640 124.470 19.040 ;
        RECT 124.830 18.240 125.190 19.440 ;
        RECT 89.550 18.180 125.190 18.240 ;
        RECT 125.490 18.180 125.830 22.640 ;
        RECT 89.550 17.840 125.830 18.180 ;
        RECT 89.550 17.380 125.190 17.440 ;
        RECT 88.910 17.040 125.190 17.380 ;
        RECT 89.550 15.840 89.910 17.040 ;
        RECT 90.270 16.240 125.190 16.640 ;
        RECT 89.550 15.440 124.470 15.840 ;
        RECT 89.550 14.240 89.910 15.440 ;
        RECT 124.830 15.040 125.190 16.240 ;
        RECT 90.270 14.640 90.630 15.040 ;
        RECT 90.990 14.640 125.190 15.040 ;
        RECT 89.550 13.840 123.390 14.240 ;
        RECT 123.750 13.840 124.470 14.240 ;
        RECT 124.830 13.440 125.190 14.640 ;
        RECT 89.550 13.380 125.190 13.440 ;
        RECT 125.490 13.380 125.830 17.840 ;
        RECT 89.550 13.040 125.830 13.380 ;
        RECT 134.880 6.300 154.740 24.700 ;
        RECT 58.830 3.920 59.750 4.260 ;
        RECT 76.510 3.920 77.430 4.260 ;
        RECT 156.565 3.500 157.155 3.525 ;
        RECT 72.490 2.900 157.160 3.500 ;
        RECT 156.565 2.875 157.155 2.900 ;
        RECT 63.470 2.085 135.080 2.090 ;
        RECT 63.470 1.495 135.105 2.085 ;
        RECT 63.470 1.490 135.080 1.495 ;
      LAYER via3 ;
        RECT 29.740 224.305 30.060 224.625 ;
        RECT 59.180 224.365 59.500 224.685 ;
        RECT 88.620 223.940 88.940 224.260 ;
        RECT 34.920 223.470 35.240 223.790 ;
        RECT 70.220 223.440 70.540 223.760 ;
        RECT 84.940 223.240 85.260 223.560 ;
        RECT 55.840 222.640 56.160 222.960 ;
        RECT 73.900 222.640 74.220 222.960 ;
        RECT 81.260 222.640 81.580 222.960 ;
        RECT 64.340 221.940 64.660 222.260 ;
        RECT 77.580 221.940 77.900 222.260 ;
        RECT 23.255 195.625 24.745 197.115 ;
        RECT 15.210 190.640 16.130 191.560 ;
        RECT 31.930 190.640 32.850 191.560 ;
        RECT 40.410 190.440 41.330 191.360 ;
        RECT 48.455 195.625 49.945 197.115 ;
        RECT 57.130 190.740 58.050 191.660 ;
        RECT 65.610 189.140 66.530 190.060 ;
        RECT 73.650 195.620 75.150 197.120 ;
        RECT 82.330 190.540 83.250 191.460 ;
        RECT 90.810 190.740 91.730 191.660 ;
        RECT 98.755 195.625 100.245 197.115 ;
        RECT 107.530 190.640 108.450 191.560 ;
        RECT 154.830 220.590 155.170 220.930 ;
        RECT 116.010 190.840 116.930 191.760 ;
        RECT 147.530 197.930 147.870 198.270 ;
        RECT 144.695 193.915 146.185 195.405 ;
        RECT 140.035 190.680 141.035 191.680 ;
        RECT 144.690 183.530 146.190 185.030 ;
        RECT 134.980 163.240 135.300 181.360 ;
        RECT 134.980 143.640 135.300 161.760 ;
        RECT 134.980 124.040 135.300 142.160 ;
        RECT 44.550 36.280 45.630 36.600 ;
        RECT 11.790 35.480 12.870 35.800 ;
        RECT 44.550 34.680 45.630 35.000 ;
        RECT 11.790 33.880 12.870 34.200 ;
        RECT 44.550 33.080 45.630 33.400 ;
        RECT 11.790 32.280 12.870 32.600 ;
        RECT 44.550 31.480 45.630 31.800 ;
        RECT 11.790 30.680 12.870 31.000 ;
        RECT 44.550 29.880 45.630 30.200 ;
        RECT 11.790 29.080 12.870 29.400 ;
        RECT 44.550 28.280 45.630 28.600 ;
        RECT 11.790 27.480 12.870 27.800 ;
        RECT 44.550 26.680 45.630 27.000 ;
        RECT 11.790 25.880 12.870 26.200 ;
        RECT 44.550 25.080 45.630 25.400 ;
        RECT 11.790 24.280 12.870 24.600 ;
        RECT 44.550 23.480 45.630 23.800 ;
        RECT 11.790 22.680 12.870 23.000 ;
        RECT 44.550 21.880 45.630 22.200 ;
        RECT 11.790 21.080 12.870 21.400 ;
        RECT 44.550 20.280 45.630 20.600 ;
        RECT 11.790 19.480 12.870 19.800 ;
        RECT 44.550 18.680 45.630 19.000 ;
        RECT 11.790 17.880 12.870 18.200 ;
        RECT 44.550 17.080 45.630 17.400 ;
        RECT 11.790 16.280 12.870 16.600 ;
        RECT 44.550 15.480 45.630 15.800 ;
        RECT 11.790 14.680 12.870 15.000 ;
        RECT 44.550 13.880 45.630 14.200 ;
        RECT 11.790 13.080 12.870 13.400 ;
        RECT 134.980 104.440 135.300 122.560 ;
        RECT 134.980 84.840 135.300 102.960 ;
        RECT 134.980 65.240 135.300 83.360 ;
        RECT 134.980 45.640 135.300 63.760 ;
        RECT 90.630 36.280 91.710 36.600 ;
        RECT 123.390 35.480 124.470 35.800 ;
        RECT 90.630 34.680 91.710 35.000 ;
        RECT 123.390 33.880 124.470 34.200 ;
        RECT 90.630 33.080 91.710 33.400 ;
        RECT 123.390 32.280 124.470 32.600 ;
        RECT 90.630 31.480 91.710 31.800 ;
        RECT 123.390 30.680 124.470 31.000 ;
        RECT 90.630 29.880 91.710 30.200 ;
        RECT 123.390 29.080 124.470 29.400 ;
        RECT 90.630 28.280 91.710 28.600 ;
        RECT 123.390 27.480 124.470 27.800 ;
        RECT 90.630 26.680 91.710 27.000 ;
        RECT 123.390 25.880 124.470 26.200 ;
        RECT 90.630 25.080 91.710 25.400 ;
        RECT 123.390 24.280 124.470 24.600 ;
        RECT 90.630 23.480 91.710 23.800 ;
        RECT 123.390 22.680 124.470 23.000 ;
        RECT 134.980 26.040 135.300 44.160 ;
        RECT 90.630 21.880 91.710 22.200 ;
        RECT 123.390 21.080 124.470 21.400 ;
        RECT 90.630 20.280 91.710 20.600 ;
        RECT 123.390 19.480 124.470 19.800 ;
        RECT 90.630 18.680 91.710 19.000 ;
        RECT 123.390 17.880 124.470 18.200 ;
        RECT 90.630 17.080 91.710 17.400 ;
        RECT 123.390 16.280 124.470 16.600 ;
        RECT 90.630 15.480 91.710 15.800 ;
        RECT 123.390 14.680 124.470 15.000 ;
        RECT 90.630 13.880 91.710 14.200 ;
        RECT 123.390 13.080 124.470 13.400 ;
        RECT 134.980 6.440 135.300 24.560 ;
        RECT 156.565 2.905 157.155 3.495 ;
        RECT 134.485 1.495 135.075 2.085 ;
      LAYER met4 ;
        RECT 147.810 224.760 147.870 225.070 ;
        RECT 7.670 224.460 7.970 224.610 ;
        RECT 11.350 224.460 11.650 224.610 ;
        RECT 15.030 224.460 15.330 224.620 ;
        RECT 18.710 224.460 19.010 224.640 ;
        RECT 29.750 224.630 30.050 224.760 ;
        RECT 59.190 224.690 59.490 224.760 ;
        RECT 22.390 224.460 22.690 224.620 ;
        RECT 26.070 224.460 26.370 224.630 ;
        RECT 3.990 224.160 28.995 224.460 ;
        RECT 29.735 224.300 30.065 224.630 ;
        RECT 33.430 224.460 33.730 224.630 ;
        RECT 37.110 224.460 37.410 224.610 ;
        RECT 40.790 224.460 41.090 224.620 ;
        RECT 44.470 224.460 44.770 224.610 ;
        RECT 48.150 224.460 48.450 224.610 ;
        RECT 51.830 224.460 52.130 224.610 ;
        RECT 55.510 224.460 55.810 224.640 ;
        RECT 33.050 224.160 57.225 224.460 ;
        RECT 59.175 224.360 59.505 224.690 ;
        RECT 28.695 223.780 34.100 223.860 ;
        RECT 34.915 223.780 35.245 223.795 ;
        RECT 28.695 223.560 35.245 223.780 ;
        RECT 62.870 223.650 63.170 224.760 ;
        RECT 66.550 224.365 66.850 224.760 ;
        RECT 64.335 224.035 66.865 224.365 ;
        RECT 33.030 223.480 35.245 223.560 ;
        RECT 34.915 223.465 35.245 223.480 ;
        RECT 55.850 223.350 63.170 223.650 ;
        RECT 55.850 222.965 56.150 223.350 ;
        RECT 55.835 222.635 56.165 222.965 ;
        RECT 64.350 222.265 64.650 224.035 ;
        RECT 70.230 223.765 70.530 224.760 ;
        RECT 70.215 223.435 70.545 223.765 ;
        RECT 73.910 222.965 74.210 224.760 ;
        RECT 73.895 222.635 74.225 222.965 ;
        RECT 77.590 222.265 77.890 224.760 ;
        RECT 81.270 222.965 81.570 224.760 ;
        RECT 84.950 223.565 85.250 224.760 ;
        RECT 88.630 224.265 88.930 224.760 ;
        RECT 147.510 224.500 147.870 224.760 ;
        RECT 88.615 223.935 88.945 224.265 ;
        RECT 84.935 223.235 85.265 223.565 ;
        RECT 81.255 222.635 81.585 222.965 ;
        RECT 64.335 221.935 64.665 222.265 ;
        RECT 77.575 221.935 77.905 222.265 ;
        RECT 147.530 198.275 147.870 224.500 ;
        RECT 154.830 224.760 154.870 225.270 ;
        RECT 154.830 220.935 155.170 224.760 ;
        RECT 154.825 220.585 155.175 220.935 ;
        RECT 147.525 197.925 147.875 198.275 ;
        RECT 73.645 197.120 75.155 197.125 ;
        RECT 2.500 195.620 121.250 197.120 ;
        RECT 73.645 195.615 75.155 195.620 ;
        RECT 119.750 195.410 121.250 195.620 ;
        RECT 119.750 193.910 154.640 195.410 ;
        RECT 7.450 190.410 156.000 191.910 ;
        RECT 65.610 190.065 66.530 190.410 ;
        RECT 65.605 189.135 66.535 190.065 ;
        RECT 11.070 36.240 46.710 36.640 ;
        RECT 11.070 35.440 45.990 35.840 ;
        RECT 11.070 34.240 11.430 35.440 ;
        RECT 46.350 35.040 46.710 36.240 ;
        RECT 11.790 34.640 46.710 35.040 ;
        RECT 11.070 33.840 45.990 34.240 ;
        RECT 11.070 32.640 11.430 33.840 ;
        RECT 46.350 33.440 46.710 34.640 ;
        RECT 11.790 33.040 46.710 33.440 ;
        RECT 89.550 36.240 125.190 36.640 ;
        RECT 89.550 35.040 89.910 36.240 ;
        RECT 90.270 35.440 125.190 35.840 ;
        RECT 89.550 34.640 124.470 35.040 ;
        RECT 89.550 33.440 89.910 34.640 ;
        RECT 124.830 34.240 125.190 35.440 ;
        RECT 90.270 33.840 125.190 34.240 ;
        RECT 89.550 33.040 124.470 33.440 ;
        RECT 124.830 32.640 125.190 33.840 ;
        RECT 11.070 32.240 46.710 32.640 ;
        RECT 89.550 32.240 125.190 32.640 ;
        RECT 11.070 31.440 46.710 31.840 ;
        RECT 11.070 30.640 45.990 31.040 ;
        RECT 11.070 29.440 11.430 30.640 ;
        RECT 46.350 30.240 46.710 31.440 ;
        RECT 11.790 29.840 46.710 30.240 ;
        RECT 11.070 29.040 45.990 29.440 ;
        RECT 11.070 27.840 11.430 29.040 ;
        RECT 46.350 28.640 46.710 29.840 ;
        RECT 11.790 28.240 46.710 28.640 ;
        RECT 89.550 31.440 125.190 31.840 ;
        RECT 89.550 30.240 89.910 31.440 ;
        RECT 90.270 30.640 125.190 31.040 ;
        RECT 89.550 29.840 124.470 30.240 ;
        RECT 89.550 28.640 89.910 29.840 ;
        RECT 124.830 29.440 125.190 30.640 ;
        RECT 90.270 29.040 125.190 29.440 ;
        RECT 89.550 28.240 124.470 28.640 ;
        RECT 124.830 27.840 125.190 29.040 ;
        RECT 11.070 27.440 46.710 27.840 ;
        RECT 89.550 27.440 125.190 27.840 ;
        RECT 11.070 26.640 46.710 27.040 ;
        RECT 11.070 25.840 45.990 26.240 ;
        RECT 11.070 24.640 11.430 25.840 ;
        RECT 46.350 25.440 46.710 26.640 ;
        RECT 11.790 25.040 46.710 25.440 ;
        RECT 11.070 24.240 45.990 24.640 ;
        RECT 11.070 23.040 11.430 24.240 ;
        RECT 46.350 23.840 46.710 25.040 ;
        RECT 11.790 23.440 46.710 23.840 ;
        RECT 89.550 26.640 125.190 27.040 ;
        RECT 89.550 25.440 89.910 26.640 ;
        RECT 90.270 25.840 125.190 26.240 ;
        RECT 89.550 25.040 124.470 25.440 ;
        RECT 89.550 23.840 89.910 25.040 ;
        RECT 124.830 24.640 125.190 25.840 ;
        RECT 90.270 24.240 125.190 24.640 ;
        RECT 89.550 23.440 124.470 23.840 ;
        RECT 124.830 23.040 125.190 24.240 ;
        RECT 11.070 22.640 46.710 23.040 ;
        RECT 89.550 22.640 125.190 23.040 ;
        RECT 11.070 21.840 46.710 22.240 ;
        RECT 11.070 21.040 45.990 21.440 ;
        RECT 11.070 19.840 11.430 21.040 ;
        RECT 46.350 20.640 46.710 21.840 ;
        RECT 11.790 20.240 46.710 20.640 ;
        RECT 11.070 19.440 45.990 19.840 ;
        RECT 11.070 18.240 11.430 19.440 ;
        RECT 46.350 19.040 46.710 20.240 ;
        RECT 11.790 18.640 46.710 19.040 ;
        RECT 89.550 21.840 125.190 22.240 ;
        RECT 89.550 20.640 89.910 21.840 ;
        RECT 90.270 21.040 125.190 21.440 ;
        RECT 89.550 20.240 124.470 20.640 ;
        RECT 89.550 19.040 89.910 20.240 ;
        RECT 124.830 19.840 125.190 21.040 ;
        RECT 90.270 19.440 125.190 19.840 ;
        RECT 89.550 18.640 124.470 19.040 ;
        RECT 124.830 18.240 125.190 19.440 ;
        RECT 11.070 17.840 46.710 18.240 ;
        RECT 89.550 17.840 125.190 18.240 ;
        RECT 11.070 17.040 46.710 17.440 ;
        RECT 11.070 16.240 45.990 16.640 ;
        RECT 11.070 15.040 11.430 16.240 ;
        RECT 46.350 15.840 46.710 17.040 ;
        RECT 11.790 15.440 46.710 15.840 ;
        RECT 11.070 14.640 45.990 15.040 ;
        RECT 11.070 13.440 11.430 14.640 ;
        RECT 46.350 14.240 46.710 15.440 ;
        RECT 11.790 13.840 46.710 14.240 ;
        RECT 89.550 17.040 125.190 17.440 ;
        RECT 89.550 15.840 89.910 17.040 ;
        RECT 90.270 16.240 125.190 16.640 ;
        RECT 89.550 15.440 124.470 15.840 ;
        RECT 89.550 14.240 89.910 15.440 ;
        RECT 124.830 15.040 125.190 16.240 ;
        RECT 90.270 14.640 125.190 15.040 ;
        RECT 89.550 13.840 124.470 14.240 ;
        RECT 124.830 13.440 125.190 14.640 ;
        RECT 11.070 13.040 46.710 13.440 ;
        RECT 89.550 13.040 125.190 13.440 ;
        RECT 134.880 5.700 135.400 190.410 ;
        RECT 144.685 183.525 146.195 185.035 ;
        RECT 144.690 181.990 146.190 183.525 ;
        RECT 145.280 181.105 145.800 181.990 ;
        RECT 136.735 163.495 154.345 181.105 ;
        RECT 145.280 161.505 145.800 163.495 ;
        RECT 136.735 143.895 154.345 161.505 ;
        RECT 145.280 141.905 145.800 143.895 ;
        RECT 136.735 124.295 154.345 141.905 ;
        RECT 145.280 122.305 145.800 124.295 ;
        RECT 136.735 104.695 154.345 122.305 ;
        RECT 145.280 102.705 145.800 104.695 ;
        RECT 136.735 85.095 154.345 102.705 ;
        RECT 145.280 83.105 145.800 85.095 ;
        RECT 136.735 65.495 154.345 83.105 ;
        RECT 145.280 63.505 145.800 65.495 ;
        RECT 136.735 45.895 154.345 63.505 ;
        RECT 145.280 43.905 145.800 45.895 ;
        RECT 136.735 26.295 154.345 43.905 ;
        RECT 145.280 24.305 145.800 26.295 ;
        RECT 136.735 6.695 154.345 24.305 ;
        RECT 145.280 5.700 145.800 6.695 ;
        RECT 134.480 1.000 135.080 2.090 ;
        RECT 156.560 1.000 157.160 3.500 ;
  END
END tt_um_TT06_SAR_wulffern
END LIBRARY

