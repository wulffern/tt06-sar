* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[1] uio_oe[2]
*+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[1] uio_out[2] uio_out[3]
*+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7] uio_oe[0] ui_in[0]
*+ uo_out[6] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3] uio_out[0]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=243.9396 ps=1.2855k w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=247.698 ps=1.29678k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VPWR tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X51 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X52 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X56 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X58 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X63 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X65 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X66 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X72 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X74 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X76 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X77 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X78 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X79 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_SAR8B_CV_0.XA6.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X88 VPWR SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X90 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X95 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X96 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X97 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X98 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X99 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R8 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X100 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X101 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X106 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X107 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X108 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X114 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X115 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X116 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X118 VGND SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X119 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R10 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X120 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X121 SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X122 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X124 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X125 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X130 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X131 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X132 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X134 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X135 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X136 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X137 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X146 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X147 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X148 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X149 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X150 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X155 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X158 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R13 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X160 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X163 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X166 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X167 SUNSAR_SAR8B_CV_0.XA4.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R14 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X169 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X174 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X175 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X176 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X177 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R15 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X178 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X181 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X182 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X185 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X186 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X188 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X193 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X194 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X195 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X198 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X199 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R16 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X201 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X205 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X206 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R17 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X207 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X212 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X213 VGND SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R18 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X214 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X216 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X221 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R19 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X223 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X225 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X228 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X229 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X230 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X232 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X233 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X235 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X236 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X237 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X239 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X246 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X253 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X255 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X263 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X266 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X268 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X270 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X275 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X276 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X278 uio_oe[0] tt_um_TT06_SAR_done_0.x4.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X280 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X282 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X284 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.XA5.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R23 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X286 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X292 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X294 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2a.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X300 uio_out[0] tt_um_TT06_SAR_done_0.x3.MN0.S VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X307 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X308 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X309 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X310 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X311 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X312 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X313 VPWR SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X314 VGND SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X316 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X318 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R24 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R25 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X321 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X322 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X324 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X328 SUNSAR_SAR8B_CV_0.XB2.XA3.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R26 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X333 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X337 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X338 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X341 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R27 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X342 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X344 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X346 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X347 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X348 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X349 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R28 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X351 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X352 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X359 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X360 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R29 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X364 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X365 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X366 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X368 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R30 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X370 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X371 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X372 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R31 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X373 SUNSAR_SAR8B_CV_0.XA3.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X374 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X375 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X376 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R32 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X377 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X378 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X379 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X381 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X382 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X384 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X385 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R33 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X386 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X387 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X389 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X390 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X391 SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X393 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R34 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X394 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X395 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X400 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X402 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X404 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X407 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X410 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R35 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R36 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X413 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X414 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X416 SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X417 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X418 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X419 SUNSAR_SAR8B_CV_0.XA20.XA10.A tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X420 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X421 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X422 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X423 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X424 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X425 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X426 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X427 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X428 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R37 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X429 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X433 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X434 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X435 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X436 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X437 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R38 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X440 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X441 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X442 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X443 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X447 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X449 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X450 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X452 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X453 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X454 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X455 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X457 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X458 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X459 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X462 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X463 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R41 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X464 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R42 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X465 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X468 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X470 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X471 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X472 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X473 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X474 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R43 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X477 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X478 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X479 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X480 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X481 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X482 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X486 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 VGND SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X489 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X491 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X492 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X493 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X494 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X496 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X498 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X499 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X500 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R44 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X501 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X502 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X503 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X505 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X506 SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X508 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X510 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X511 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X512 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X513 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X514 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X515 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R46 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X516 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X517 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X519 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X520 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X521 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X522 SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X525 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X526 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X527 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X528 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X530 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X532 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R47 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X533 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2a.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X536 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X537 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X540 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X541 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R48 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X544 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X545 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X548 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R49 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X553 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X554 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X557 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X558 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X560 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X561 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X562 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X564 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X565 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X567 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X568 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X570 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X571 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X572 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X573 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X574 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X575 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_CAPT8B_CV_0.XA2.MP0.G SUNSAR_CAPT8B_CV_0.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X578 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X579 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X580 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X581 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X582 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X583 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X584 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X587 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X588 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X589 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X590 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X591 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X592 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X593 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X594 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X595 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R51 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X596 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X598 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X601 SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X602 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R52 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X603 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X604 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X605 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X606 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X609 VGND SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X610 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X613 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X614 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X616 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X618 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X619 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X621 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X624 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X626 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X631 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X637 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X640 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R53 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X642 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X644 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R54 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X645 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X647 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X648 SUNSAR_SAR8B_CV_0.XA7.XA6.MP0.D SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X649 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X650 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X652 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X653 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R55 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X654 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X656 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X657 VGND SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X658 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X661 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X663 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X664 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X665 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X666 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R57 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X667 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X669 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2a.A VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X670 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X674 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X675 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X676 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X680 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X681 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X682 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X683 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X684 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X685 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X686 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X687 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X688 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X690 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R58 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X691 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X693 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X694 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X695 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X696 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X697 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X699 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X700 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X701 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X704 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X705 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X706 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X707 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X709 VGND tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X710 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X713 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X714 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X715 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X716 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R60 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X717 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X718 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X719 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X720 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X721 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X722 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R61 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X726 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X727 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X728 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X729 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X730 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X731 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X732 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X734 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X735 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X738 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X740 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X741 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R62 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X742 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X745 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X746 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X747 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X749 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X751 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X752 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X753 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R65 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X754 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X755 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 SUNSAR_SAR8B_CV_0.XA2.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X759 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X760 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X762 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X763 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X765 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X766 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X767 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X768 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X770 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X771 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X773 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X774 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X777 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X778 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X779 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X780 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X782 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R67 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X783 VGND SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X786 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X787 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R68 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X788 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X790 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X791 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X792 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X793 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X798 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X800 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X802 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X809 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X810 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X813 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X814 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X816 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X817 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X818 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X819 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X821 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X822 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X823 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X824 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X825 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X828 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X829 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X830 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X831 SUNSAR_SAR8B_CV_0.XA0.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X832 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X833 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X834 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X835 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X836 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X837 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X838 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X839 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X842 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X843 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X844 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X845 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R70 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X847 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X848 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X849 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X850 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X852 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X853 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X854 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X855 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X858 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X859 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X862 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X864 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X867 SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X868 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X872 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X873 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X874 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X875 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X876 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X878 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X879 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VGND SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X883 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X884 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X886 VGND SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X887 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VPWR SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X890 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X892 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R71 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X893 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X894 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X895 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X896 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2a.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X897 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X899 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X901 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R72 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X902 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X903 VGND SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X905 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R73 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X906 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X909 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X910 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R74 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X911 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X912 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X913 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X914 tt_um_TT06_SAR_done_0.x4.MN0.G tt_um_TT06_SAR_done_0.x4.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X915 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X917 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R75 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X918 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X920 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X923 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X924 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X925 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X926 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X928 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X929 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R76 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X930 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X931 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X932 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X933 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X934 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X935 uio_out[0] tt_um_TT06_SAR_done_0.x3.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X936 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X937 SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X939 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X940 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X941 SUNSAR_SAR8B_CV_0.XA1.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X942 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R77 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X944 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X945 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X946 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X947 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R78 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X948 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X949 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X950 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X951 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X953 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X954 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X955 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X957 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XB1.XA3.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X959 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X961 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X962 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R79 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X963 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X964 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X965 VGND SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X967 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 TIE_L SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X970 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X971 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X972 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X974 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R80 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X975 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X976 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X978 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X980 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X982 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X984 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X985 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X986 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X987 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X988 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X993 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R81 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X994 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X995 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X997 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X999 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1000 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1001 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1002 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1004 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1005 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R82 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1008 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1013 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1014 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R83 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1016 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1018 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1019 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1020 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1021 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1022 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1025 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1033 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1034 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1035 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1036 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1037 SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1038 SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1039 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1040 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1041 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1042 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1043 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1044 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1045 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1046 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1047 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1048 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1049 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1050 VGND tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1051 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1052 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1053 SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1054 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 a_15210_29612# VPWR 0.397362f
C1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.CK 0.524159f
C2 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 1.77563f
C3 VPWR a_13842_37180# 0.473697f
C4 a_22770_29964# SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.134249f
C5 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_2768# 0.172147f
C6 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.596437f
C7 VPWR a_18882_32956# 0.436368f
C8 VPWR a_15230_40296# 0.455577f
C9 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO 0.144331f
C10 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VPWR 1.06875f
C11 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.432466f
C12 a_5130_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C13 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA2.Y 0.241356f
C14 VPWR a_23942_42760# 0.388156f
C15 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.16676f
C16 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.39041f
C17 VPWR a_18882_35420# 0.39968f
C18 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.324243f
C19 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN 0.143148f
C20 a_6282_28556# SUNSAR_SAR8B_CV_0.XA1.ENO 0.135353f
C21 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.246146f
C22 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S 0.106927f
C23 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.55251f
C24 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.ENO 0.503825f
C25 SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR 0.665006f
C26 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.07223f
C27 VPWR a_13862_40296# 0.457343f
C28 VPWR a_5150_40648# 0.492592f
C29 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR 0.104609f
C30 TIE_L1 uo_out[7] 0.206895f
C31 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D VPWR 0.137646f
C32 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y a_12710_42408# 0.100131f
C33 VPWR a_20250_36300# 0.395776f
C34 VPWR a_10170_36300# 0.398846f
C35 a_3762_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C36 a_10170_32076# VPWR 0.436368f
C37 VPWR a_10190_41880# 0.395781f
C38 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.649845f
C39 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C40 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.45828f
C41 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO 0.152052f
C42 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.SARN 13.6519f
C43 TIE_L1 TIE_L 0.257793f
C44 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C45 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.305131f
C46 VPWR a_3782_40648# 0.491225f
C47 TIE_L1 VPWR 0.114647f
C48 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43816# 0.127669f
C49 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35068# 0.127528f
C50 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VPWR 1.05322f
C51 a_15210_27500# VPWR 0.382397f
C52 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.104933f
C53 VPWR a_18882_36300# 0.399161f
C54 VPWR a_8802_36300# 0.399161f
C55 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C56 a_8802_32076# VPWR 0.436368f
C57 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA8.A 0.527529f
C58 VPWR a_8822_41880# 0.395781f
C59 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.744161f
C60 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.109613f
C61 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO 0.339883f
C62 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C63 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.449584f
C64 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.CKN 0.200119f
C65 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 1.77562f
C66 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.SARN 13.6523f
C67 VPWR a_10170_37180# 0.474068f
C68 a_9990_4566# VPWR 0.413433f
C69 VPWR a_15210_32956# 0.436368f
C70 SUNSAR_CAPT8B_CV_0.XA4.MP1.G SUNSAR_CAPT8B_CV_0.XA4.Y 0.206292f
C71 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.318734f
C72 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D VPWR 0.138148f
C73 a_13842_27500# VPWR 0.382189f
C74 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.791379f
C75 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D 0.112858f
C76 VPWR a_20270_42760# 0.391454f
C77 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.52234f
C78 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189112f
C79 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 2.59087f
C80 VPWR a_15210_35420# 0.39968f
C81 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C82 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CN1 0.466806f
C83 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.133602f
C84 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.101001f
C85 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 2.95303f
C86 VPWR a_8802_37180# 0.473729f
C87 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_3728# 0.172147f
C88 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VPWR 0.452478f
C89 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C90 VPWR a_13842_32956# 0.436368f
C91 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C92 VPWR a_10190_40296# 0.455675f
C93 VPWR tt_um_TT06_SAR_done_0.DONE 8.46867f
C94 SUNSAR_CAPT8B_CV_0.XG12.QN a_16382_43816# 0.129239f
C95 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VPWR 1.06875f
C96 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.432466f
C97 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.464697f
C98 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D 0.112858f
C99 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA6.CEO 0.381914f
C100 VPWR a_18902_42760# 0.391454f
C101 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C102 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 2.2622f
C103 VPWR a_13842_35420# 0.39968f
C104 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C105 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.449584f
C106 a_2610_28556# SUNSAR_SAR8B_CV_0.XA0.ENO 0.132757f
C107 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.CKN 0.41624f
C108 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.D<5> 0.102632f
C109 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.2165f
C110 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.ENO 0.438277f
C111 VPWR a_8822_40296# 0.457343f
C112 VPWR a_23942_41000# 0.390551f
C113 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VPWR 0.271482f
C114 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO 0.144331f
C115 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D VPWR 0.137646f
C116 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.12241f
C117 VPWR a_15210_36300# 0.398846f
C118 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 4.24508f
C119 VPWR a_5130_36300# 0.398846f
C120 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.375196f
C121 a_5130_32076# VPWR 0.436368f
C122 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.276413f
C123 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO 0.154232f
C124 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C125 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CN1 0.466806f
C126 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.133602f
C127 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 0.250503f
C128 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S 0.106927f
C129 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.309657f
C130 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C131 VPWR a_5150_41000# 0.388161f
C132 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VPWR 1.05322f
C133 a_10170_27500# VPWR 0.382397f
C134 VPWR a_13842_36300# 0.399161f
C135 VPWR a_3762_36300# 0.399161f
C136 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.241356f
C137 a_3762_32076# VPWR 0.436368f
C138 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA7.ENO 0.152518f
C139 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.63636f
C140 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO 0.3401f
C141 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.431984f
C142 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 2.95304f
C143 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.249907f
C144 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.SARN 3.57448f
C145 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.ENO 0.793076f
C146 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR 0.519052f
C147 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.11382f
C148 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.587991f
C149 VPWR a_10170_32956# 0.436368f
C150 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR 0.104609f
C151 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35068# 0.129098f
C152 VPWR a_3782_41000# 0.388256f
C153 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D VPWR 0.138148f
C154 a_8802_27500# VPWR 0.382189f
C155 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR 0.104609f
C156 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.393125f
C157 VPWR tt_um_TT06_SAR_done_0.x3.MN0.S 0.695784f
C158 VPWR a_15230_42760# 0.391454f
C159 VPWR a_10170_35420# 0.39968f
C160 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 3.07164f
C161 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CN1 0.466806f
C162 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.133602f
C163 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 1.77562f
C164 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_4688# 0.172147f
C165 a_16542_4918# VPWR 0.470354f
C166 VPWR a_8802_32956# 0.436368f
C167 VPWR a_5150_40296# 0.455605f
C168 VPWR a_20270_41000# 0.388156f
C169 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VPWR 0.271482f
C170 TIE_L2 uo_out[7] 0.100011f
C171 SUNSAR_CAPT8B_CV_0.XF11.QN a_12710_43816# 0.127669f
C172 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO 0.144331f
C173 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VPWR 1.06875f
C174 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C175 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 4.25322f
C176 VPWR a_23922_36652# 0.449853f
C177 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.284482f
C178 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.383512f
C179 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR 0.618979f
C180 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA6.ENO 0.150467f
C181 VPWR a_28727_40659# 0.39147f
C182 VPWR a_13862_42760# 0.391454f
C183 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.744161f
C184 VPWR a_8802_35420# 0.39968f
C185 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S 0.106927f
C186 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.86675f
C187 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.ENO 0.503825f
C188 VPWR a_3782_40296# 0.457343f
C189 VPWR a_18902_41000# 0.388256f
C190 VPWR a_23942_41352# 0.376408f
C191 a_23922_28556# VPWR 0.499441f
C192 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.12241f
C193 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA5.CEO 0.303978f
C194 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR 0.324111f
C195 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA8.A 0.527529f
C196 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.SARN 5.22744f
C197 ui_in[0] SUNSAR_SAR8B_CV_0.EN 0.969482f
C198 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARN 0.64474f
C199 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.649845f
C200 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.10225f
C201 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C202 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CN1 0.466806f
C203 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.133602f
C204 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.M3.G 0.224309f
C205 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN 0.538639f
C206 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.EN 2.96993f
C207 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.EN 1.15994f
C208 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR 0.519052f
C209 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C210 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43816# 0.129239f
C211 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.432466f
C212 a_5130_27500# VPWR 0.382397f
C213 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR 0.104609f
C214 clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.438597f
C215 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.CEO 0.13078f
C216 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR 2.30036f
C217 VPWR tt_um_TT06_SAR_done_0.x4.MN0.G 0.511762f
C218 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.137745f
C219 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.233892f
C220 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C221 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.227625f
C222 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.246063f
C223 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 1.77562f
C224 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.D<7> 0.187721f
C225 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.ENO 1.2771f
C226 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.545186f
C227 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VPWR 0.452478f
C228 VPWR a_5130_32956# 0.436368f
C229 VPWR a_23942_40648# 0.489579f
C230 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR 0.104609f
C231 a_3762_27500# VPWR 0.382189f
C232 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D 0.112858f
C233 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA3.CEO 0.303978f
C234 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR 2.31184f
C235 VPWR a_28727_41011# 0.468616f
C236 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA5.ENO 0.104122f
C237 VPWR a_10190_42760# 0.391454f
C238 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C239 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.162703f
C240 VPWR a_5130_35420# 0.39968f
C241 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CN1 0.466806f
C242 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.133602f
C243 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 0.305131f
C244 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 2.95308f
C245 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_5648# 0.172147f
C246 VPWR a_3762_32956# 0.436368f
C247 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C248 VPWR a_15230_41000# 0.388156f
C249 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35068# 0.127528f
C250 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.321724f
C251 a_20250_28556# VPWR 0.406628f
C252 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.791351f
C253 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C254 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D 0.112858f
C255 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.CEO 0.13078f
C256 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA4.CEO 0.352238f
C257 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR 2.31184f
C258 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA5.ENO 0.155821f
C259 VPWR a_8822_42760# 0.391454f
C260 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.155424f
C261 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.26537f
C262 VPWR a_3762_35420# 0.39968f
C263 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.40569f
C264 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.412143f
C265 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.118152f
C266 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1615f
C267 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.ENO 0.434116f
C268 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_2928# 0.105547f
C269 a_9990_4918# VPWR 0.468783f
C270 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.62595f
C271 VPWR a_13862_41000# 0.388256f
C272 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO 0.144331f
C273 a_18882_28556# VPWR 0.406628f
C274 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y a_7670_42408# 0.100131f
C275 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.310451f
C276 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR 2.31184f
C277 VPWR a_28727_41363# 0.440399f
C278 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.268769f
C279 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2165f
C280 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO 0.152052f
C281 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C282 a_21422_41000# SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.115667f
C283 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S 0.106927f
C284 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.170578f
C285 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2a.A 4.93712f
C286 VPWR a_20270_40648# 0.492579f
C287 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C288 ua[0] SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.247314f
C289 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.432466f
C290 a_20250_27852# VPWR 0.358413f
C291 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 3.09787f
C292 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA2.CEO 0.352238f
C293 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR 2.31184f
C294 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA4.ENO 0.150467f
C295 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C296 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.63636f
C297 VPWR SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.106794f
C298 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> 0.595738f
C299 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.CKN 0.200119f
C300 a_20270_41000# SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.156079f
C301 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 2.95307f
C302 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.166192f
C303 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.ENO 1.2771f
C304 VPWR a_23922_33132# 0.415713f
C305 VPWR a_18902_40648# 0.491225f
C306 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.267144f
C307 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VPWR 0.271482f
C308 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP 0.123668f
C309 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.12241f
C310 a_18882_27852# VPWR 0.358599f
C311 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR 0.104609f
C312 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.276413f
C313 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.375196f
C314 VPWR a_23942_40296# 0.453754f
C315 VPWR a_5150_42760# 0.391454f
C316 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.119314f
C317 VPWR SUNSAR_SAR8B_CV_0.XA7.XA10.Y 0.718455f
C318 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.658328f
C319 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.146458f
C320 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.227625f
C321 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA8.A 0.527529f
C322 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 1.77562f
C323 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.30523f
C324 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.166272f
C325 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_6608# 0.172147f
C326 a_16542_5270# VPWR 0.489055f
C327 VPWR a_10190_41000# 0.388175f
C328 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO 0.144331f
C329 a_15210_28556# VPWR 0.406628f
C330 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.791379f
C331 VPWR a_20250_34716# 0.396749f
C332 VPWR a_5150_41352# 0.394053f
C333 VPWR a_3782_42760# 0.391454f
C334 VPWR a_20270_41352# 0.394053f
C335 VPWR SUNSAR_SAR8B_CV_0.XA4.XA10.Y 0.725614f
C336 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S 0.101562f
C337 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.166192f
C338 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S 0.106927f
C339 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.245678f
C340 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.205884f
C341 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6519f
C342 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.ENO 0.491653f
C343 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_3888# 0.105547f
C344 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 2.66621f
C345 VPWR a_8822_41000# 0.388256f
C346 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR 0.104609f
C347 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.143554f
C348 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35068# 0.129098f
C349 a_13842_28556# VPWR 0.406628f
C350 ui_in[0] SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.172623f
C351 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.694484f
C352 VPWR a_18882_34716# 0.399819f
C353 VPWR a_3782_41352# 0.394053f
C354 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.204048f
C355 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA3.ENO 0.104122f
C356 VPWR a_18902_41352# 0.394053f
C357 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L 1.05246f
C358 VPWR SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.722887f
C359 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.119314f
C360 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C361 VPWR SUNSAR_SAR8B_CV_0.XA7.XA8.A 1.20972f
C362 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 0.635098f
C363 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C364 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C365 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.166272f
C366 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.238636f
C367 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 2.64055f
C368 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VPWR 0.271482f
C369 clk SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.210661f
C370 SUNSAR_SAR8B_CV_0.SARP ua[1] 1.01251f
C371 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.209352f
C372 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR 0.104609f
C373 VPWR a_23942_44344# 0.342053f
C374 SUNSAR_SAR8B_CV_0.XA7.XA11.Y a_21402_36828# 0.104051f
C375 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.284482f
C376 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.383512f
C377 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA3.ENO 0.155821f
C378 VPWR a_20270_40296# 0.455248f
C379 VPWR SUNSAR_SAR8B_CV_0.CK_SAMPLE 9.398339f
C380 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_34540# 0.103065f
C381 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.704356f
C382 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.101979f
C383 VPWR SUNSAR_SAR8B_CV_0.XA6.XA10.Y 0.725614f
C384 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.924613f
C385 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> 0.625035f
C386 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y 0.22339f
C387 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.227625f
C388 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.166192f
C389 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 1.77562f
C390 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.ENO 1.2771f
C391 a_9990_5270# VPWR 0.490626f
C392 SUNSAR_SAR8B_CV_0.XA20.XA2a.A SUNSAR_SAR8B_CV_0.XA20.XA2.CO 1.43919f
C393 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 2.64054f
C394 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.12241f
C395 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA1.CEO 0.303978f
C396 VPWR SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.635621f
C397 tt_um_TT06_SAR_done_0.x3.MN0.S tt_um_TT06_SAR_done_0.DONE 0.186749f
C398 VPWR a_18902_40296# 0.457343f
C399 VPWR SUNSAR_SAR8B_CV_0.EN 41.9219f
C400 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.119314f
C401 VPWR SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.722887f
C402 VPWR SUNSAR_SAR8B_CV_0.XA6.XA8.A 1.22023f
C403 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.M3.G 0.224309f
C404 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C405 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C406 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN 0.206912f
C407 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 2.95303f
C408 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR 0.808658f
C409 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 2.64055f
C410 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.419738f
C411 a_10170_28556# VPWR 0.406628f
C412 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.432466f
C413 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.200058f
C414 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.11641f
C415 VPWR a_15210_34716# 0.399819f
C416 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.CEO 0.13078f
C417 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA2.ENO 0.150467f
C418 VPWR a_15230_41352# 0.394053f
C419 VPWR a_23942_43112# 0.393308f
C420 VPWR SUNSAR_SAR8B_CV_0.XA2.XA10.Y 0.725614f
C421 a_13842_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C422 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C423 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.4271f
C424 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.101979f
C425 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C426 a_18902_41000# SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.15757f
C427 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.205884f
C428 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.251051f
C429 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.55251f
C430 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.ENO 0.11341f
C431 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_4848# 0.105547f
C432 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 2.64054f
C433 VPWR a_10190_43816# 0.391817f
C434 SUNSAR_CAPT8B_CV_0.XA4.MP1.G SUNSAR_CAPT8B_CV_0.XA3.Y 0.300065f
C435 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR 0.104609f
C436 a_8802_28556# VPWR 0.406628f
C437 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.EN 0.176398f
C438 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.143675f
C439 VPWR a_13842_34716# 0.399819f
C440 VPWR SUNSAR_SAR8B_CV_0.D<0> 5.48841f
C441 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.112859f
C442 VPWR a_13862_41352# 0.394053f
C443 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C444 VPWR SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.722887f
C445 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C446 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1615f
C447 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.930839f
C448 a_17750_41000# SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.114097f
C449 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S 0.106927f
C450 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.XA2.Y 0.306905f
C451 a_10170_28908# VPWR 0.395394f
C452 VPWR a_5150_44168# 0.340085f
C453 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.419738f
C454 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.7271f
C455 VPWR a_8822_43816# 0.391817f
C456 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.145738f
C457 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35068# 0.127528f
C458 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN 0.253395f
C459 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.144778f
C460 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.180903f
C461 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA0.CEO 0.352238f
C462 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S 0.106927f
C463 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.11263f
C464 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.63636f
C465 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.11536f
C466 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.101979f
C467 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> 0.625175f
C468 a_15210_28908# VPWR 0.395394f
C469 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 2.95305f
C470 a_8802_28908# VPWR 0.395394f
C471 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_2768# 0.172147f
C472 a_16542_5622# VPWR 0.472384f
C473 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C474 a_15210_27852# VPWR 0.358413f
C475 a_10170_28204# VPWR 0.361706f
C476 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.72582f
C477 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN 0.24816f
C478 VPWR a_5150_41880# 0.395781f
C479 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C480 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR 0.104609f
C481 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.139471f
C482 SUNSAR_SAR8B_CV_0.XA6.XA11.Y a_17730_36828# 0.10248f
C483 VPWR a_15230_44168# 0.340085f
C484 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S 0.106927f
C485 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.242472f
C486 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA1.ENO 0.104122f
C487 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA4.A 1.63909f
C488 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.55251f
C489 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.119314f
C490 a_10170_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C491 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C492 VPWR SUNSAR_SAR8B_CV_0.XA5.XA8.A 1.2202f
C493 a_13842_28908# VPWR 0.395394f
C494 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.227625f
C495 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C496 SUNSAR_SAR8B_CV_0.XA7.XA10.Y a_21402_36300# 0.13402f
C497 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA2.Y 1.77562f
C498 a_12690_36300# SUNSAR_SAR8B_CV_0.XA4.XA10.Y 0.13253f
C499 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.301485f
C500 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.738812f
C501 a_13842_27852# VPWR 0.358599f
C502 a_8802_28204# VPWR 0.36179f
C503 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 2.72889f
C504 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35420# 0.160931f
C505 VPWR a_3782_41880# 0.395781f
C506 a_18882_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C507 a_5130_28556# VPWR 0.406628f
C508 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.432466f
C509 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.791351f
C510 VPWR a_10170_34716# 0.399819f
C511 VPWR a_13862_44168# 0.3405f
C512 VPWR SUNSAR_SAR8B_CV_0.D<1> 5.18522f
C513 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.204048f
C514 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA1.ENO 0.155821f
C515 VPWR a_10190_41352# 0.394053f
C516 a_8802_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C517 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.ENO 0.328435f
C518 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.ENO 0.252047f
C519 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.93081f
C520 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.205884f
C521 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S 0.106927f
C522 a_16542_5974# VPWR 0.449888f
C523 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_5808# 0.105547f
C524 VPWR a_5150_43816# 0.391817f
C525 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN 0.248827f
C526 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VPWR 0.271482f
C527 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_20250_35420# 0.133834f
C528 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.143554f
C529 a_3762_28556# VPWR 0.406628f
C530 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.12241f
C531 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y a_2630_42408# 0.100131f
C532 a_10190_41880# SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 0.100592f
C533 VPWR a_8802_34716# 0.399819f
C534 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.276252f
C535 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.375025f
C536 VPWR a_8822_41352# 0.394053f
C537 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.SARN 13.6519f
C538 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C539 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.ENO 0.693521f
C540 VPWR SUNSAR_SAR8B_CV_0.XA4.XA8.A 1.22023f
C541 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.ENO 1.11884f
C542 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<2> 0.137975f
C543 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.440586f
C544 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.437693f
C545 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C546 a_16382_41000# SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.115667f
C547 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.308722f
C548 a_5130_28908# VPWR 0.395394f
C549 a_11322_36300# SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.13402f
C550 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.738798f
C551 VPWR a_20250_33836# 0.407174f
C552 VPWR a_3782_43816# 0.391817f
C553 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.118162f
C554 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR 0.104609f
C555 SUNSAR_SAR8B_CV_0.XA5.XA11.Y a_16362_36828# 0.104051f
C556 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.ENO 0.150467f
C557 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA4.A 1.63909f
C558 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.233892f
C559 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31666f
C560 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.297144f
C561 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.ENO 0.820808f
C562 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.ENO 1.18612f
C563 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> 0.625035f
C564 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.227625f
C565 a_15230_41000# SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.156079f
C566 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 1.77562f
C567 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.248979f
C568 a_3762_28908# VPWR 0.395394f
C569 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.153964f
C570 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_3728# 0.172147f
C571 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23942_42760# 0.101843f
C572 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR 0.808658f
C573 a_10170_27852# VPWR 0.358413f
C574 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C575 ua[0] SUNSAR_SAR8B_CV_0.SARN 1.02347f
C576 VPWR a_18882_33836# 0.409601f
C577 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.204048f
C578 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN 0.249322f
C579 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR 0.104609f
C580 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35068# 0.129098f
C581 a_15210_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C582 VPWR SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 1.20019f
C583 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C584 VPWR SUNSAR_SAR8B_CV_0.D<2> 5.20829f
C585 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 54.2165f
C586 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.111867f
C587 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.ENO 0.6934f
C588 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.ENO 1.03123f
C589 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C590 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.930839f
C591 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.506551f
C592 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 2.9531f
C593 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.CK 1.59176f
C594 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.740872f
C595 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22790_42760# 0.13379f
C596 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.301485f
C597 a_8802_27852# VPWR 0.358599f
C598 ua[1] SUNSAR_SAR8B_CV_0.SARN 0.806872f
C599 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.449584f
C600 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.393665f
C601 VPWR SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 11.7505f
C602 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VPWR 0.271482f
C603 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_18882_35420# 0.133834f
C604 a_20250_28908# VPWR 0.395394f
C605 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 3.86364f
C606 VPWR a_5130_34716# 0.399819f
C607 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S 0.106927f
C608 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.204048f
C609 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.ENO 0.820808f
C610 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.ENO 1.18612f
C611 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<3> 0.105016f
C612 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.437693f
C613 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.22339f
C614 VPWR SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.765792f
C615 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.205884f
C616 a_9990_5622# VPWR 0.470814f
C617 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C618 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.254583f
C619 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_6768# 0.105547f
C620 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN 0.267395f
C621 a_22790_41880# SUNSAR_CAPT8B_CV_0.XA4.Y 0.111538f
C622 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.241356f
C623 VPWR a_23942_43992# 0.388156f
C624 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.437693f
C625 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35420# 0.160931f
C626 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.106927f
C627 a_18882_28908# VPWR 0.395394f
C628 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.12241f
C629 VPWR a_3762_34716# 0.399819f
C630 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S 0.106927f
C631 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA4.A 1.63909f
C632 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.174995f
C633 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.182408f
C634 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.ENO 0.6934f
C635 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C636 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.ENO 1.03123f
C637 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C638 VPWR SUNSAR_SAR8B_CV_0.XA3.XA8.A 1.2202f
C639 SUNSAR_SAR8B_CV_0.XA6.XA10.Y a_17730_36300# 0.13253f
C640 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR 0.104609f
C641 VPWR a_15210_33836# 0.409601f
C642 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.449584f
C643 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.145738f
C644 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.106927f
C645 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.432466f
C646 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.649845f
C647 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.290432f
C648 VPWR SUNSAR_SAR8B_CV_0.D<3> 5.17056f
C649 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.102131f
C650 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.4471f
C651 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.63636f
C652 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.475004f
C653 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y 0.342913f
C654 VPWR SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.728421f
C655 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.291229f
C656 a_16542_2630# VPWR 0.448659f
C657 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.93081f
C658 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.ENO 0.820808f
C659 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.ENO 1.18612f
C660 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> 0.625175f
C661 VPWR a_20270_43816# 0.391817f
C662 a_9990_5974# VPWR 0.451043f
C663 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_4688# 0.172147f
C664 a_5130_27852# VPWR 0.358413f
C665 VPWR a_13842_33836# 0.409601f
C666 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.204048f
C667 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR 0.104609f
C668 VPWR SUNSAR_CAPT8B_CV_0.XI14.QN 0.901631f
C669 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN 0.248612f
C670 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.437693f
C671 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.744161f
C672 SUNSAR_SAR8B_CV_0.SARP VPWR 0.139564f
C673 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.146492f
C674 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK 3.91346f
C675 SUNSAR_SAR8B_CV_0.XA4.XA11.Y a_12690_36828# 0.10248f
C676 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.215804f
C677 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP 0.252966f
C678 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON a_20250_30316# 0.127528f
C679 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.EN 0.131572f
C680 VPWR SUNSAR_SAR8B_CV_0.XB1.TIE_L 7.37316f
C681 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 6.86675f
C682 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C683 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.ENO 1.03107f
C684 VPWR SUNSAR_SAR8B_CV_0.XA2.XA8.A 1.22023f
C685 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.ENO 0.6934f
C686 a_2610_31196# SUNSAR_SAR8B_CV_0.D<7> 0.11099f
C687 SUNSAR_SAR8B_CV_0.XA5.XA10.Y a_16362_36300# 0.13402f
C688 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.227625f
C689 VPWR a_18902_43816# 0.391817f
C690 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR 0.104609f
C691 a_7650_36300# SUNSAR_SAR8B_CV_0.XA2.XA10.Y 0.13253f
C692 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA6.ENO 0.291697f
C693 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.301485f
C694 a_23922_26796# VPWR 0.442318f
C695 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.153964f
C696 a_3762_27852# VPWR 0.358599f
C697 VPWR SUNSAR_CAPT8B_CV_0.XH13.QN 0.901622f
C698 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35068# 0.127528f
C699 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C700 VPWR a_23922_34892# 0.395601f
C701 a_13950_4390# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.15559f
C702 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA4.A 1.63909f
C703 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_22790_43640# 0.127669f
C704 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.D<7> 0.240612f
C705 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.D<7> 0.180455f
C706 a_13862_41000# SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.15757f
C707 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.205884f
C708 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C709 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN 0.248535f
C710 VPWR SUNSAR_CAPT8B_CV_0.XG12.QN 0.901622f
C711 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.143554f
C712 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.106927f
C713 a_20250_29612# VPWR 0.398044f
C714 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<0> 0.492001f
C715 VPWR SUNSAR_SAR8B_CV_0.D<4> 5.15123f
C716 a_12582_4390# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.15559f
C717 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON a_18882_30316# 0.129098f
C718 VPWR a_20250_36828# 0.392512f
C719 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.145483f
C720 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.930839f
C721 a_12710_41000# SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.114097f
C722 a_6282_36300# SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.13402f
C723 VPWR a_10170_33836# 0.409601f
C724 VPWR SUNSAR_CAPT8B_CV_0.XF11.QN 0.901622f
C725 VPWR a_20270_44168# 0.340085f
C726 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35420# 0.160931f
C727 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.106927f
C728 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.432466f
C729 VPWR SUNSAR_SAR8B_CV_0.XA7.ENO 4.77251f
C730 SUNSAR_SAR8B_CV_0.XA3.XA11.Y a_11322_36828# 0.104051f
C731 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S 0.106927f
C732 VPWR a_18882_36828# 0.395703f
C733 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> 1.08082f
C734 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C735 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.227625f
C736 VPWR a_15230_43816# 0.391817f
C737 SUNSAR_CAPT8B_CV_0.XI14.XA4.A a_20270_42760# 0.111734f
C738 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C739 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_5648# 0.172147f
C740 a_20250_26796# VPWR 0.441753f
C741 VPWR a_8802_33836# 0.409601f
C742 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VPWR 0.271482f
C743 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.241356f
C744 VPWR SUNSAR_CAPT8B_CV_0.XE10.QN 0.901622f
C745 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN 0.258218f
C746 VPWR a_18902_44168# 0.3405f
C747 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_15210_35420# 0.133834f
C748 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.12241f
C749 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 0.724217f
C750 VPWR SUNSAR_SAR8B_CV_0.XA6.ENO 5.54203f
C751 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.182595f
C752 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S 0.106927f
C753 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.102131f
C754 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA4.A 1.63909f
C755 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 27.1615f
C756 a_9990_2630# VPWR 0.447504f
C757 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.EN 0.176792f
C758 VPWR SUNSAR_SAR8B_CV_0.XA1.XA8.A 1.2202f
C759 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.201839f
C760 ua[1] ua[0] 3.85017f
C761 VPWR a_13862_43816# 0.391817f
C762 a_6302_41000# SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.115667f
C763 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.301485f
C764 a_18882_26796# VPWR 0.442908f
C765 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C766 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 1.62434f
C767 VPWR SUNSAR_CAPT8B_CV_0.XD09.QN 0.901622f
C768 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.393049f
C769 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.530644f
C770 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 4.0111f
C771 VPWR SUNSAR_SAR8B_CV_0.XA5.ENO 4.84607f
C772 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<1> 0.297507f
C773 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2165f
C774 VPWR SUNSAR_SAR8B_CV_0.D<5> 5.14531f
C775 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C776 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.204048f
C777 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA7.ENO 0.30776f
C778 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.42393f
C779 SUNSAR_SAR8B_CV_0.XB2.XA3.B ua[0] 0.241597f
C780 a_16542_2982# VPWR 0.490338f
C781 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.93081f
C782 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C783 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.205884f
C784 a_5150_41000# SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.156079f
C785 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN 0.263255f
C786 VPWR SUNSAR_CAPT8B_CV_0.XC08.QN 0.901622f
C787 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C788 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.106927f
C789 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.744161f
C790 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C791 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 0.722427f
C792 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.324105f
C793 VPWR SUNSAR_SAR8B_CV_0.XA4.ENO 5.52623f
C794 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.151329f
C795 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON a_15210_30316# 0.127528f
C796 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA6.ENO 0.128204f
C797 clk SUNSAR_CAPT8B_CV_0.XA4.Y 0.206733f
C798 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARN 0.591428f
C799 VPWR a_15210_36828# 0.395582f
C800 SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S ua[0] 0.100365f
C801 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.ENO 0.10132f
C802 VPWR SUNSAR_SAR8B_CV_0.XA0.XA8.A 1.22398f
C803 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<6> 0.199516f
C804 a_11342_41000# SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.115667f
C805 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.318734f
C806 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C807 VPWR a_5130_33836# 0.409601f
C808 a_20250_30316# VPWR 0.403745f
C809 VPWR SUNSAR_CAPT8B_CV_0.XB07.QN 0.901622f
C810 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C811 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_13842_35420# 0.133834f
C812 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.106927f
C813 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.649845f
C814 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.2199f
C815 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.227341f
C816 VPWR SUNSAR_SAR8B_CV_0.XA3.ENO 4.84607f
C817 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.CEO 0.138f
C818 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA4.A 1.63909f
C819 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.63636f
C820 VPWR a_13842_36828# 0.395703f
C821 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA1.ENO 0.34399f
C822 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> 1.20727f
C823 a_10190_41000# SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.156079f
C824 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN 0.112859f
C825 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.SARN 1.62434f
C826 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_2928# 0.105547f
C827 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_6608# 0.172147f
C828 a_15210_26796# VPWR 0.441753f
C829 SUNSAR_CAPT8B_CV_0.XH13.XA4.A a_18902_42760# 0.113305f
C830 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C831 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.204048f
C832 VPWR a_3762_33836# 0.409601f
C833 VPWR SUNSAR_CAPT8B_CV_0.XA2.MP0.G 0.667429f
C834 a_18882_30316# VPWR 0.403802f
C835 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C836 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35420# 0.160931f
C837 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.398331f
C838 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.SARN 0.103734f
C839 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 0.722417f
C840 VPWR SUNSAR_SAR8B_CV_0.XA2.ENO 5.52623f
C841 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.158152f
C842 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<2> 0.297715f
C843 SUNSAR_SAR8B_CV_0.XA2.XA11.Y a_7650_36828# 0.10248f
C844 VPWR SUNSAR_SAR8B_CV_0.D<6> 5.17441f
C845 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON a_13842_30316# 0.129098f
C846 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA6.ENO 0.363295f
C847 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6519f
C848 SUNSAR_SAR8B_CV_0.XB1.XA3.B ua[1] 0.241597f
C849 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.ENO 0.193518f
C850 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.D<0> 0.215251f
C851 tt_um_TT06_SAR_done_0.DONE SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.227625f
C852 uio_oe[0] uio_out[0] 1.55761f
C853 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN 0.11263f
C854 a_13842_26796# VPWR 0.442908f
C855 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.301485f
C856 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.M3.G 0.263588f
C857 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.25689f
C858 VPWR SUNSAR_SAR8B_CV_0.XA1.ENO 4.84607f
C859 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C860 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S 0.106927f
C861 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.107567f
C862 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.1501f
C863 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.204048f
C864 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.107674f
C865 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.232115f
C866 SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S ua[1] 0.100365f
C867 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.ENO 0.238862f
C868 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<7> 0.178111f
C869 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.106828f
C870 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN 0.112859f
C871 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.205884f
C872 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C873 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.94014f
C874 VPWR SUNSAR_SAR8B_CV_0.SARN 0.132799f
C875 a_22790_41000# SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.11811f
C876 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C877 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.106927f
C878 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.118161f
C879 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.79343f
C880 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C881 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 0.722427f
C882 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO 0.15234f
C883 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.220689f
C884 VPWR SUNSAR_SAR8B_CV_0.XA0.ENO 5.52718f
C885 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S 0.106927f
C886 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_3334# 0.120042f
C887 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA4.A 1.63909f
C888 VPWR a_10170_36828# 0.396003f
C889 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.174995f
C890 a_9990_2982# VPWR 0.491909f
C891 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<7> 2.50324f
C892 clk uio_out[0] 0.120689f
C893 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN 0.11263f
C894 VPWR a_23922_35948# 0.390687f
C895 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.105035f
C896 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.393063f
C897 a_15210_30316# VPWR 0.404384f
C898 a_15210_31196# VPWR 0.44007f
C899 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C900 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.106927f
C901 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.129613f
C902 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.227352f
C903 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO 0.340491f
C904 SUNSAR_SAR8B_CV_0.XA1.XA11.Y a_6282_36828# 0.104051f
C905 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<3> 0.297504f
C906 VPWR SUNSAR_SAR8B_CV_0.D<7> 3.61291f
C907 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.109137f
C908 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_3334# 0.113134f
C909 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA5.ENO 0.316693f
C910 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.233892f
C911 VPWR a_8802_36828# 0.396052f
C912 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.726497f
C913 a_16542_3334# VPWR 0.380282f
C914 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> 0.746324f
C915 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.419738f
C916 uo_out[0] uio_out[0] 0.201579f
C917 clk uio_oe[0] 0.260056f
C918 a_3782_41000# SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.15757f
C919 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_3888# 0.105547f
C920 a_10170_26796# VPWR 0.441753f
C921 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.241356f
C922 a_13842_31196# VPWR 0.44007f
C923 a_13842_30316# VPWR 0.404384f
C924 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.118226f
C925 VPWR a_20250_35068# 0.391458f
C926 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 0.722417f
C927 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.377598f
C928 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.CMP_OP 7.93512f
C929 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON a_10170_30316# 0.127528f
C930 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA4.ENO 0.126806f
C931 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.55251f
C932 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.D<1> 0.228326f
C933 a_5130_29612# VPWR 0.397362f
C934 uo_out[0] uio_oe[0] 0.670799f
C935 clk ui_in[0] 0.169609f
C936 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.318734f
C937 a_2630_41000# SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.114097f
C938 a_8802_26796# VPWR 0.442908f
C939 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.301485f
C940 VPWR SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.405511f
C941 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35420# 0.160931f
C942 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.527529f
C943 VPWR a_23942_42408# 0.3915f
C944 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.649845f
C945 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.13041f
C946 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.394834f
C947 VPWR a_18882_35068# 0.394528f
C948 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1615f
C949 VPWR a_23942_41880# 0.398828f
C950 a_13950_4742# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.156331f
C951 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_2982# 0.158066f
C952 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA4.A 1.63909f
C953 SUNSAR_CAPT8B_CV_0.XA5.XA2.A a_22790_42408# 0.10248f
C954 a_3762_29612# VPWR 0.397362f
C955 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.419738f
C956 a_8822_41000# SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.15757f
C957 uo_out[1] uio_oe[0] 0.432144f
C958 SUNSAR_CAPT8B_CV_0.XG12.XA4.A a_15230_42760# 0.111734f
C959 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C960 VPWR a_20250_35948# 0.414756f
C961 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 1.70987f
C962 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.183415f
C963 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C964 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_10170_35420# 0.133834f
C965 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.744161f
C966 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.118161f
C967 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.293159f
C968 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<4> 0.297602f
C969 a_12582_4742# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.156331f
C970 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON a_8802_30316# 0.129098f
C971 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA4.ENO 0.363295f
C972 VPWR a_5130_36828# 0.395767f
C973 a_7670_41000# SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.114097f
C974 uo_out[2] uio_oe[0] 0.267754f
C975 a_2610_36300# SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.13253f
C976 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.205975f
C977 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.107823f
C978 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.589705f
C979 VPWR a_18882_35948# 0.417826f
C980 a_10170_31196# VPWR 0.44007f
C981 a_10170_30316# VPWR 0.404384f
C982 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C983 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.205884f
C984 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 5.19722f
C985 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CP0 0.331282f
C986 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.638386f
C987 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.280191f
C988 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.CEO 0.432008f
C989 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.110962f
C990 VPWR SUNSAR_CAPT8B_CV_0.XA4.Y 1.18734f
C991 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.63636f
C992 VPWR a_3762_36828# 0.395857f
C993 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y a_21422_42408# 0.113479f
C994 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR 0.337652f
C995 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO 0.127551f
C996 uo_out[3] uio_oe[0] 0.212351f
C997 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN 0.36754f
C998 a_5130_26796# VPWR 0.441753f
C999 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_4848# 0.105547f
C1000 VPWR a_3782_44168# 0.3405f
C1001 a_8802_31196# VPWR 0.44007f
C1002 a_8802_30316# VPWR 0.404384f
C1003 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C1004 VPWR a_5130_37180# 0.474051f
C1005 VPWR a_20270_42408# 0.391292f
C1006 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.152045f
C1007 VPWR a_15210_35068# 0.394528f
C1008 SUNSAR_SAR8B_CV_0.XA0.XA11.Y a_2610_36828# 0.10248f
C1009 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.158152f
C1010 VPWR a_20270_41880# 0.395781f
C1011 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP 0.435464f
C1012 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.55251f
C1013 a_9990_3334# VPWR 0.380282f
C1014 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.175642f
C1015 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK 0.331207f
C1016 a_23922_29964# VPWR 0.429137f
C1017 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.D<2> 0.228332f
C1018 uo_out[5] uio_out[0] 0.109219f
C1019 uo_out[4] uio_oe[0] 0.550054f
C1020 uo_out[1] uo_out[0] 0.355472f
C1021 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18344f
C1022 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.318734f
C1023 a_3762_26796# VPWR 0.442908f
C1024 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.301485f
C1025 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 4.36162f
C1026 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.178114f
C1027 VPWR a_3762_37180# 0.473713f
C1028 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_8802_35420# 0.133834f
C1029 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C1030 VPWR a_18902_42408# 0.391292f
C1031 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA4.Y 0.504864f
C1032 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO 0.152052f
C1033 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.SARN 13.6519f
C1034 VPWR a_13842_35068# 0.394528f
C1035 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<5> 0.297941f
C1036 VPWR a_18902_41880# 0.395781f
C1037 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C1038 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_2982# 0.158066f
C1039 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.379175p
C1040 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA3.ENO 0.316693f
C1041 VPWR a_20270_43288# 0.394205f
C1042 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.714341f
C1043 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.55251f
C1044 VPWR ua[0] 0.51729f
C1045 uo_out[5] uio_oe[0] 1.55329f
C1046 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.EN 0.315968f
C1047 SUNSAR_CAPT8B_CV_0.XF11.XA4.A a_13862_42760# 0.113305f
C1048 VPWR a_15210_35948# 0.417826f
C1049 VPWR a_23922_34540# 0.502044f
C1050 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.241356f
C1051 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35420# 0.160931f
C1052 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA8.A 0.527529f
C1053 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO 0.339883f
C1054 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.220689f
C1055 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.702226f
C1056 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON a_5130_30316# 0.127528f
C1057 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C1058 a_22770_28556# SUNSAR_SAR8B_CV_0.XA20.XA1.CK 0.140127f
C1059 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA2.ENO 0.126806f
C1060 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.26479f
C1061 VPWR a_18902_43288# 0.394205f
C1062 VPWR SUNSAR_SAR8B_CV_0.XA7.CEO 1.1111f
C1063 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.372599f
C1064 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.108751f
C1065 VPWR ua[1] 0.225132f
C1066 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARN 0.175967f
C1067 a_23922_27148# VPWR 0.483246f
C1068 VPWR a_13842_35948# 0.417826f
C1069 a_5130_31196# VPWR 0.44007f
C1070 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.393049f
C1071 a_5130_30316# VPWR 0.404384f
C1072 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.327152f
C1073 uio_out[0] TIE_L 0.44106f
C1074 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_3334# 0.114704f
C1075 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3334# 0.163985f
C1076 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S 0.669708f
C1077 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.723713f
C1078 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y a_17750_42408# 0.111909f
C1079 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR 1.56028f
C1080 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.449584f
C1081 uo_out[7] uio_oe[0] 0.43252f
C1082 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1083 VPWR uio_out[0] 0.408488f
C1084 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_5808# 0.105547f
C1085 a_20250_28204# VPWR 0.361706f
C1086 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.179089f
C1087 a_3762_31196# VPWR 0.44007f
C1088 a_3762_30316# VPWR 0.404384f
C1089 VPWR a_20250_37532# 0.454392f
C1090 VPWR a_15230_42408# 0.391292f
C1091 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.15651f
C1092 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C1093 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.744161f
C1094 VPWR a_10170_35068# 0.394528f
C1095 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<6> 0.298165f
C1096 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.377598f
C1097 VPWR a_15230_41880# 0.395781f
C1098 uio_oe[0] TIE_L 1.21913f
C1099 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON a_3762_30316# 0.129098f
C1100 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.702226f
C1101 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.255261f
C1102 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.189429f
C1103 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C1104 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA2.ENO 0.363295f
C1105 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_3334# 0.118471f
C1106 VPWR SUNSAR_SAR8B_CV_0.XA6.CEO 2.28789f
C1107 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.2165f
C1108 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.126354f
C1109 SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S VPWR 0.183853f
C1110 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.D<3> 0.228326f
C1111 VPWR uio_oe[0] 1.67769f
C1112 uo_out[3] uo_out[2] 0.109993f
C1113 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.386137f
C1114 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.301485f
C1115 a_18882_28204# VPWR 0.36179f
C1116 VPWR a_18882_37532# 0.458267f
C1117 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C1118 VPWR a_13862_42408# 0.391292f
C1119 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.649845f
C1120 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C1121 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C1122 VPWR a_8802_35068# 0.394528f
C1123 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO 0.154232f
C1124 VPWR a_13862_41880# 0.395781f
C1125 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.267238f
C1126 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.191868f
C1127 VPWR a_15230_43288# 0.394205f
C1128 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.720096f
C1129 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.787331f
C1130 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.ENO 0.118161f
C1131 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y a_16382_42408# 0.113479f
C1132 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR 1.5612f
C1133 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.449584f
C1134 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.2165f
C1135 VPWR ui_in[0] 1.85366f
C1136 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.29297f
C1137 a_20250_27148# VPWR 0.470364f
C1138 VPWR a_10170_35948# 0.417826f
C1139 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR 6.88568f
C1140 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR 6.94539f
C1141 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.449584f
C1142 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.122781f
C1143 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.380687f
C1144 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO 0.3401f
C1145 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.293159f
C1146 clk TIE_L 0.146712f
C1147 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.702226f
C1148 a_13950_5094# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.160184f
C1149 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_4038# 0.135393f
C1150 a_21402_28556# SUNSAR_SAR8B_CV_0.XA7.ENO 0.134248f
C1151 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.147435f
C1152 VPWR a_13862_43288# 0.394205f
C1153 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.164325f
C1154 VPWR SUNSAR_SAR8B_CV_0.XA5.CEO 1.0603f
C1155 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO 0.13041f
C1156 SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S VPWR 0.183853f
C1157 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.175642f
C1158 uo_out[4] uo_out[3] 0.854997f
C1159 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1160 VPWR clk 0.644902f
C1161 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.318734f
C1162 a_18882_27148# VPWR 0.471462f
C1163 VPWR a_8802_35948# 0.417826f
C1164 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D 0.112098f
C1165 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.178114f
C1166 a_23922_30844# VPWR 0.425847f
C1167 a_23922_31724# VPWR 0.412398f
C1168 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C1169 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35420# 0.160931f
C1170 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.327909f
C1171 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.CEO 0.432008f
C1172 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<7> 0.294651f
C1173 uo_out[0] TIE_L 0.280844f
C1174 a_12582_5094# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.160184f
C1175 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3334# 0.163985f
C1176 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3686# 0.16579f
C1177 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA1.ENO 0.316693f
C1178 SUNSAR_CAPT8B_CV_0.XA4.MP1.G SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.138433f
C1179 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.63636f
C1180 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.723728f
C1181 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO 0.118161f
C1182 a_16542_4038# VPWR 0.379979f
C1183 SUNSAR_SAR8B_CV_0.XB2.M3.G ua[0] 0.765539f
C1184 VPWR uo_out[0] 1.02382f
C1185 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_6768# 0.105547f
C1186 SUNSAR_CAPT8B_CV_0.XE10.XA4.A a_10190_42760# 0.111734f
C1187 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y a_5150_41880# 0.100592f
C1188 a_15210_28204# VPWR 0.361706f
C1189 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.88588f
C1190 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.231927f
C1191 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D 0.112858f
C1192 a_20270_41880# SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.100592f
C1193 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.449584f
C1194 VPWR a_15210_37532# 0.459479f
C1195 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_5130_35420# 0.133834f
C1196 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.143023f
C1197 VPWR a_10190_42408# 0.391292f
C1198 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C1199 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.26609f
C1200 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C1201 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.158152f
C1202 VPWR a_5130_35068# 0.394528f
C1203 uo_out[1] TIE_L 0.50141f
C1204 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.702226f
C1205 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.ENO 0.126806f
C1206 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.EN 0.207932f
C1207 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.86675f
C1208 VPWR SUNSAR_SAR8B_CV_0.XA4.CEO 2.30385f
C1209 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO 0.129613f
C1210 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.D<4> 0.228332f
C1211 VPWR uo_out[1] 1.02322f
C1212 uo_out[5] uo_out[4] 1.16093f
C1213 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.107427f
C1214 a_13842_28204# VPWR 0.36179f
C1215 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.30589f
C1216 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 4.24834f
C1217 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR 2.45124f
C1218 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.393055f
C1219 SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR 2.62711f
C1220 VPWR a_13842_37532# 0.458324f
C1221 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA8.A 0.527529f
C1222 VPWR a_8822_42408# 0.391292f
C1223 VPWR a_3762_35068# 0.394528f
C1224 uo_out[2] TIE_L 0.156661f
C1225 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.26479f
C1226 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.126085f
C1227 VPWR a_10190_43288# 0.394205f
C1228 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.720133f
C1229 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO 0.118226f
C1230 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y a_12710_42408# 0.111909f
C1231 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.86675f
C1232 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1233 VPWR uo_out[2] 1.02322f
C1234 uo_out[6] uo_out[4] 0.843602f
C1235 a_15210_27148# VPWR 0.470364f
C1236 VPWR a_5130_35948# 0.417826f
C1237 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.231927f
C1238 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.179089f
C1239 SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR 2.62329f
C1240 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR 2.44986f
C1241 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 0.241356f
C1242 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142977f
C1243 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C1244 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN 0.473354f
C1245 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.220689f
C1246 uo_out[3] TIE_L 0.185333f
C1247 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C1248 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.702226f
C1249 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.441867f
C1250 a_17730_28556# SUNSAR_SAR8B_CV_0.XA6.ENO 0.132757f
C1251 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S 0.669708f
C1252 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.379175p
C1253 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.ENO 0.363295f
C1254 VPWR a_8822_43288# 0.394205f
C1255 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C1256 VPWR SUNSAR_SAR8B_CV_0.XA3.CEO 1.06031f
C1257 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO 0.13041f
C1258 VPWR uo_out[3] 1.25759f
C1259 uo_out[7] uo_out[4] 0.121648f
C1260 uo_out[6] uo_out[5] 0.327382f
C1261 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.318734f
C1262 a_13842_27148# VPWR 0.471462f
C1263 VPWR a_3762_35948# 0.417826f
C1264 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.11826f
C1265 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.504801f
C1266 SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR 2.62342f
C1267 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR 2.45309f
C1268 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C1269 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_3762_35420# 0.133834f
C1270 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.649845f
C1271 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.327152f
C1272 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.149144f
C1273 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN 0.145339f
C1274 uo_out[4] TIE_L 0.31941f
C1275 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3686# 0.16579f
C1276 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.233892f
C1277 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.723762f
C1278 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38576f
C1279 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C1280 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y a_11342_42408# 0.113479f
C1281 SUNSAR_SAR8B_CV_0.XB1.M3.G ua[1] 0.762388f
C1282 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO 0.118161f
C1283 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.40569f
C1284 uo_out[7] uo_out[5] 1.57818f
C1285 VPWR uo_out[4] 1.03021f
C1286 SUNSAR_CAPT8B_CV_0.XD09.XA4.A a_8822_42760# 0.113305f
C1287 a_23922_30844# SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.100515f
C1288 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 4.25569f
C1289 SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR 2.62342f
C1290 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR 2.45309f
C1291 VPWR a_10170_37532# 0.459599f
C1292 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35420# 0.160931f
C1293 VPWR a_5150_42408# 0.391292f
C1294 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142956f
C1295 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.744161f
C1296 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C1297 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 2.1352f
C1298 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.377598f
C1299 uo_out[5] TIE_L 1.3092f
C1300 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.74594f
C1301 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.441867f
C1302 a_16362_28556# SUNSAR_SAR8B_CV_0.XA5.ENO 0.135353f
C1303 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.109021f
C1304 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.143148f
C1305 VPWR SUNSAR_SAR8B_CV_0.XA2.CEO 2.30393f
C1306 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1615f
C1307 a_9990_4038# VPWR 0.379979f
C1308 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO 0.129613f
C1309 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87301f
C1310 uo_out[7] uo_out[6] 2.38922f
C1311 VPWR uo_out[5] 1.02721f
C1312 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1313 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C1314 a_5130_28204# VPWR 0.361706f
C1315 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.386137f
C1316 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y a_17750_42408# 0.100131f
C1317 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.B 1.13456f
C1318 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.178114f
C1319 SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR 2.62342f
C1320 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.386305f
C1321 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.294852f
C1322 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR 2.45309f
C1323 VPWR a_8802_37532# 0.458443f
C1324 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C1325 VPWR a_3782_42408# 0.391292f
C1326 VPWR SUNSAR_SAR8B_CV_0.XA6.DONE 0.246222f
C1327 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2165f
C1328 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO 0.152052f
C1329 uo_out[6] TIE_L 0.204625f
C1330 a_13950_5446# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.102604f
C1331 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C1332 VPWR a_5150_43288# 0.394205f
C1333 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.720114f
C1334 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR 2.50821f
C1335 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO 0.118226f
C1336 a_20250_29612# SUNSAR_SAR8B_CV_0.EN 0.142592f
C1337 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C1338 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.ENO 0.116058f
C1339 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 27.1615f
C1340 VPWR uo_out[6] 1.34623f
C1341 a_3762_28204# VPWR 0.36179f
C1342 a_10170_27148# VPWR 0.470364f
C1343 VPWR SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.774301f
C1344 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR 2.62393f
C1345 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR 2.45309f
C1346 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C1347 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA8.A 0.527529f
C1348 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142977f
C1349 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO 0.339883f
C1350 VPWR SUNSAR_SAR8B_CV_0.XA5.DONE 0.245452f
C1351 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.293159f
C1352 uo_out[7] TIE_L 0.471918f
C1353 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.748719f
C1354 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C1355 a_12582_5446# SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.101033f
C1356 VPWR a_3782_43288# 0.394205f
C1357 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.245678f
C1358 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2173f
C1359 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.CEO 0.301665f
C1360 VPWR SUNSAR_SAR8B_CV_0.XA1.CEO 1.0603f
C1361 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.57155f
C1362 SUNSAR_SAR8B_CV_0.XB2.CKN VPWR 2.34497f
C1363 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.ENO 0.13041f
C1364 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.849501f
C1365 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.ENO 0.111173f
C1366 TIE_L1 uio_oe[0] 0.902557f
C1367 VPWR uo_out[7] 1.27659f
C1368 a_8802_27148# VPWR 0.471462f
C1369 VPWR SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.780003f
C1370 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR 2.62403f
C1371 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR 2.45309f
C1372 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.686731f
C1373 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C1374 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.327909f
C1375 VPWR SUNSAR_SAR8B_CV_0.XA4.DONE 0.246222f
C1376 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.CEO 0.432008f
C1377 VPWR TIE_L 0.387688f
C1378 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.305166f
C1379 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.EN 0.37807f
C1380 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.63636f
C1381 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.728492f
C1382 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y a_7670_42408# 0.111909f
C1383 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.433299f
C1384 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.ENO 0.111217f
C1385 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.ENO 0.893904f
C1386 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1387 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO 0.144331f
C1388 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR 0.429492f
C1389 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.474658f
C1390 VPWR SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.779986f
C1391 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.535136f
C1392 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.133602f
C1393 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.179089f
C1394 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.241356f
C1395 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR 2.45309f
C1396 VPWR a_5130_37532# 0.459538f
C1397 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C1398 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.257526f
C1399 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.898003f
C1400 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142956f
C1401 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.09966f
C1402 VPWR SUNSAR_SAR8B_CV_0.XA3.DONE 0.245452f
C1403 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.158152f
C1404 a_12690_28556# SUNSAR_SAR8B_CV_0.XA4.ENO 0.132757f
C1405 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_4038# 0.135393f
C1406 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.426291f
C1407 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6519f
C1408 VPWR SUNSAR_SAR8B_CV_0.XA0.CEO 2.30575f
C1409 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.ENO 0.409858f
C1410 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.ENO 0.111173f
C1411 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.ENO 0.952619f
C1412 VPWR a_15230_40648# 0.492579f
C1413 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.318734f
C1414 a_13842_29612# VPWR 0.397362f
C1415 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D VPWR 0.137646f
C1416 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.134182f
C1417 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.107427f
C1418 VPWR SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.780003f
C1419 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D 0.112858f
C1420 a_20250_32076# VPWR 0.433941f
C1421 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.393076f
C1422 VPWR a_3762_37532# 0.458382f
C1423 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C1424 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.898003f
C1425 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.165965f
C1426 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.136678f
C1427 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.17528f
C1428 VPWR SUNSAR_SAR8B_CV_0.XA2.DONE 0.246222f
C1429 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO 0.154232f
C1430 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.303428f
C1431 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C1432 VPWR SUNSAR_CAPT8B_CV_0.XA3.Y 0.86364f
C1433 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.41635f
C1434 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y a_6302_42408# 0.113479f
C1435 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 2.31184f
C1436 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.ENO 0.111217f
C1437 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.ENO 1.02916f
C1438 VPWR a_13862_40648# 0.491225f
C1439 ui_in[0] tt_um_TT06_SAR_done_0.DONE 0.198829f
C1440 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6519f
C1441 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.142061f
C1442 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VPWR 1.06002f
C1443 a_5130_27148# VPWR 0.470364f
C1444 SUNSAR_CAPT8B_CV_0.XC08.XA4.A a_5150_42760# 0.111734f
C1445 VPWR SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.779986f
C1446 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.559553f
C1447 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.133602f
C1448 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D 0.112858f
C1449 a_18882_32076# VPWR 0.436368f
C1450 a_20250_31196# VPWR 0.437f
C1451 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142977f
C1452 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.898003f
C1453 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.744161f
C1454 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.297363f
C1455 VPWR SUNSAR_SAR8B_CV_0.XA1.DONE 0.245452f
C1456 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO 0.3401f
C1457 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.244517f
C1458 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.419738f
C1459 a_11322_28556# SUNSAR_SAR8B_CV_0.XA3.ENO 0.135353f
C1460 VPWR a_23942_43640# 0.412992f
C1461 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C1462 VPWR a_20250_37180# 0.469114f
C1463 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.98135f
C1464 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 2.31184f
C1465 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.ENO 0.111173f
C1466 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.ENO 0.952619f
C1467 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1468 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D VPWR 0.138148f
C1469 a_3762_27148# VPWR 0.471462f
C1470 VPWR SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.780003f
C1471 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 4.2492f
C1472 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.375196f
C1473 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.276413f
C1474 a_18882_31196# VPWR 0.44007f
C1475 VPWR a_28727_39955# 0.355584f
C1476 uio_out[0] tt_um_TT06_SAR_done_0.x3.MN0.S 0.165429f
C1477 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.898003f
C1478 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.649845f
C1479 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.19724f
C1480 VPWR SUNSAR_SAR8B_CV_0.XA0.DONE 0.247527f
C1481 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.250503f
C1482 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.305131f
C1483 VPWR a_18882_37180# 0.473682f
C1484 SUNSAR_SAR8B_CV_0.XB1.CKN VPWR 2.34497f
C1485 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 2.31184f
C1486 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C1487 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.ENO 0.111217f
C1488 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.ENO 1.02916f
C1489 a_10170_29612# VPWR 0.397362f
C1490 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VPWR 1.06875f
C1491 VPWR SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.779986f
C1492 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.133602f
C1493 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C1494 a_15230_41880# SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.100592f
C1495 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.898003f
C1496 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142956f
C1497 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80606f
C1498 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.18614f
C1499 VPWR a_23922_35420# 0.416528f
C1500 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.178114f
C1501 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.419738f
C1502 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.SARN 0.108405f
C1503 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.CKN 0.41624f
C1504 a_18882_29612# VPWR 0.397362f
C1505 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.245678f
C1506 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.55251f
C1507 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.TIE_L 4.28648f
C1508 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.ENO 0.438277f
C1509 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR 2.50821f
C1510 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO 4.6743f
C1511 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.ENO 0.952619f
C1512 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.ENO 0.111173f
C1513 VPWR a_10190_40648# 0.492624f
C1514 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.318734f
C1515 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO 0.144331f
C1516 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35068# 0.129098f
C1517 a_8802_29612# VPWR 0.397362f
C1518 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D VPWR 0.137646f
C1519 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C1520 VPWR SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.784656f
C1521 a_15210_32076# VPWR 0.436368f
C1522 VPWR a_28727_40307# 0.410063f
C1523 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA8.A 0.527529f
C1524 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.898003f
C1525 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.665724f
C1526 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.145048f
C1527 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1615f
C1528 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S 0.101001f
C1529 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S 0.106927f
C1530 VPWR a_10190_44168# 0.340085f
C1531 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y a_2630_42408# 0.111909f
C1532 SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR 0.665006f
C1533 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C1534 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233744f
C1535 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C1536 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.ENO 1.04628f
C1537 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.55549f
C1538 VPWR a_8822_40648# 0.491225f
C1539 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR 0.108436f
C1540 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.174845f
C1541 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43816# 0.129239f
C1542 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VPWR 1.05322f
C1543 a_20250_27500# VPWR 0.382397f
C1544 SUNSAR_CAPT8B_CV_0.XB07.XA4.A a_3782_42760# 0.113305f
C1545 VPWR a_23922_36300# 0.472384f
C1546 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 4.27988f
C1547 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C1548 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.383512f
C1549 a_13842_32076# VPWR 0.436368f
C1550 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.284482f
C1551 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.142977f
C1552 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.898003f
C1553 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.109613f
C1554 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.131536f
C1555 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.159359f
C1556 a_7650_28556# SUNSAR_SAR8B_CV_0.XA2.ENO 0.132757f
C1557 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 2.95296f
C1558 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1625f
C1559 VPWR a_8822_44168# 0.3405f
C1560 VPWR a_15210_37180# 0.474036f
C1561 a_23922_29964# SUNSAR_SAR8B_CV_0.XA20.XA2a.A 0.151031f
C1562 a_16542_4566# VPWR 0.413433f
C1563 VPWR a_20250_32956# 0.433941f
C1564 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VPWR 0.279205f
C1565 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.EN 0.343905f
C1566 TIE_L1 uo_out[5] 0.275794f
C1567 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D VPWR 0.138148f
C1568 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.12241f
C1569 a_18882_27500# VPWR 0.382189f
C1570 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.671839f
C1571 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C1572 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.293873f
C1573 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.39306f
C1574 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.898003f
C1575 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.34383f
C1576 VPWR a_20250_35420# 0.39661f
C1577 ua[2] VGND 0.117454f
C1578 ua[3] VGND 0.117454f
C1579 ua[4] VGND 0.118698f
C1580 ua[5] VGND 0.120088f
C1581 ua[6] VGND 0.120088f
C1582 ua[7] VGND 0.111009f
C1583 ua[0] VGND 7.62793f
C1584 ua[1] VGND 6.98581f
C1585 uio_out[0] VGND 8.52142f
C1586 uio_oe[0] VGND 7.87718f
C1587 ui_in[0] VGND 5.40407f
C1588 clk VGND 6.22723f
C1589 uo_out[0] VGND 2.40292f
C1590 uo_out[1] VGND 1.50319f
C1591 uo_out[2] VGND 1.42895f
C1592 uo_out[3] VGND 1.68048f
C1593 uo_out[4] VGND 1.55276f
C1594 uo_out[5] VGND 1.75883f
C1595 uo_out[6] VGND 2.73387f
C1596 uo_out[7] VGND 3.23518f
C1597 VPWR VGND 0.949773p
C1598 TIE_L1 VGND 1.33691f
C1599 TIE_L2 VGND 1.67804f
C1600 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93609f
C1601 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93609f
C1602 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.5533f
C1603 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.5533f
C1604 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.334839f
C1605 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.334839f
C1606 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.469f
C1607 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.469f
C1608 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43533f
C1609 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43533f
C1610 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67745f
C1611 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67745f
C1612 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.6684f
C1613 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.6684f
C1614 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.574499f
C1615 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.574499f
C1616 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33412f
C1617 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33412f
C1618 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.469f
C1619 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.469f
C1620 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43533f
C1621 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43533f
C1622 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67745f
C1623 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67745f
C1624 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.6684f
C1625 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.6684f
C1626 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.575099f
C1627 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.575099f
C1628 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33412f
C1629 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33412f
C1630 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.469f
C1631 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.469f
C1632 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43533f
C1633 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43533f
C1634 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67745f
C1635 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67745f
C1636 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.6684f
C1637 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.6684f
C1638 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.571799f
C1639 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.571799f
C1640 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33412f
C1641 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33412f
C1642 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.471901f
C1643 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.471901f
C1644 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.439809f
C1645 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44253f
C1646 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.3859f
C1647 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.38266f
C1648 a_15390_2630# VGND 0.542161f $ **FLOATING
C1649 a_13950_2630# VGND 0.427094f $ **FLOATING
C1650 a_12582_2630# VGND 0.426679f $ **FLOATING
C1651 a_11142_2630# VGND 0.543317f $ **FLOATING
C1652 a_15390_2982# VGND 0.491607f $ **FLOATING
C1653 a_13950_2982# VGND 0.352472f $ **FLOATING
C1654 a_12582_2982# VGND 0.352472f $ **FLOATING
C1655 a_11142_2982# VGND 0.490037f $ **FLOATING
C1656 a_15390_3334# VGND 0.374919f $ **FLOATING
C1657 a_13950_3334# VGND 0.352438f $ **FLOATING
C1658 a_12582_3334# VGND 0.352438f $ **FLOATING
C1659 a_11142_3334# VGND 0.374919f $ **FLOATING
C1660 a_13950_3686# VGND 0.352418f $ **FLOATING
C1661 a_12582_3686# VGND 0.352418f $ **FLOATING
C1662 SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND 41.5268f
C1663 SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.S VGND 0.70146f
C1664 SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND 41.5268f
C1665 SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.S VGND 0.70146f
C1666 a_15390_4038# VGND 0.397033f $ **FLOATING
C1667 a_13950_4038# VGND 0.354407f $ **FLOATING
C1668 a_12582_4038# VGND 0.354407f $ **FLOATING
C1669 a_11142_4038# VGND 0.397033f $ **FLOATING
C1670 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VGND 37.7832f
C1671 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.38998f
C1672 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND 0.103625f
C1673 a_13950_4390# VGND 0.352432f $ **FLOATING
C1674 a_12582_4390# VGND 0.352432f $ **FLOATING
C1675 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND 0.103625f
C1676 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.38998f
C1677 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VGND 37.7832f
C1678 SUNSAR_SAR8B_CV_0.XB2.M3.G VGND 3.1165f
C1679 a_15390_4566# VGND 0.389036f $ **FLOATING
C1680 SUNSAR_SAR8B_CV_0.XB1.M3.G VGND 3.07938f
C1681 a_11142_4566# VGND 0.389036f $ **FLOATING
C1682 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VGND 0.970036f
C1683 a_13950_4742# VGND 0.352456f $ **FLOATING
C1684 a_12582_4742# VGND 0.352456f $ **FLOATING
C1685 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND 0.7964f
C1686 a_15390_4918# VGND 0.470144f $ **FLOATING
C1687 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND 0.7964f
C1688 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VGND 0.970036f
C1689 a_11142_4918# VGND 0.471715f $ **FLOATING
C1690 a_13950_5094# VGND 0.353103f $ **FLOATING
C1691 a_12582_5094# VGND 0.353103f $ **FLOATING
C1692 a_15390_5270# VGND 0.492927f $ **FLOATING
C1693 a_11142_5270# VGND 0.491356f $ **FLOATING
C1694 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND 0.596866f
C1695 a_13950_5446# VGND 0.433341f $ **FLOATING
C1696 a_12582_5446# VGND 0.433756f $ **FLOATING
C1697 a_15390_5622# VGND 0.47219f $ **FLOATING
C1698 a_15390_5974# VGND 0.541341f $ **FLOATING
C1699 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND 0.596866f
C1700 a_11142_5622# VGND 0.47376f $ **FLOATING
C1701 a_11142_5974# VGND 0.540186f $ **FLOATING
C1702 a_22770_26796# VGND 0.529341f $ **FLOATING
C1703 a_21402_26796# VGND 0.531659f $ **FLOATING
C1704 a_17730_26796# VGND 0.530834f $ **FLOATING
C1705 a_16362_26796# VGND 0.531989f $ **FLOATING
C1706 a_12690_26796# VGND 0.530834f $ **FLOATING
C1707 a_11322_26796# VGND 0.531989f $ **FLOATING
C1708 a_7650_26796# VGND 0.530213f $ **FLOATING
C1709 a_6282_26796# VGND 0.530979f $ **FLOATING
C1710 a_2610_26796# VGND 0.531178f $ **FLOATING
C1711 a_22770_27148# VGND 0.499848f $ **FLOATING
C1712 a_21402_27148# VGND 0.467094f $ **FLOATING
C1713 a_17730_27148# VGND 0.471508f $ **FLOATING
C1714 a_16362_27148# VGND 0.467722f $ **FLOATING
C1715 a_12690_27148# VGND 0.471508f $ **FLOATING
C1716 a_11322_27148# VGND 0.467722f $ **FLOATING
C1717 a_7650_27148# VGND 0.470266f $ **FLOATING
C1718 a_6282_27148# VGND 0.465734f $ **FLOATING
C1719 a_2610_27148# VGND 0.47123f $ **FLOATING
C1720 a_21402_27500# VGND 0.385968f $ **FLOATING
C1721 a_17730_27500# VGND 0.387712f $ **FLOATING
C1722 a_16362_27500# VGND 0.386249f $ **FLOATING
C1723 a_12690_27500# VGND 0.387712f $ **FLOATING
C1724 a_11322_27500# VGND 0.386249f $ **FLOATING
C1725 a_7650_27500# VGND 0.38671f $ **FLOATING
C1726 a_6282_27500# VGND 0.384229f $ **FLOATING
C1727 a_2610_27500# VGND 0.387675f $ **FLOATING
C1728 a_21402_27852# VGND 0.370125f $ **FLOATING
C1729 a_17730_27852# VGND 0.370785f $ **FLOATING
C1730 a_16362_27852# VGND 0.368771f $ **FLOATING
C1731 a_12690_27852# VGND 0.370785f $ **FLOATING
C1732 a_11322_27852# VGND 0.368771f $ **FLOATING
C1733 a_7650_27852# VGND 0.369543f $ **FLOATING
C1734 a_6282_27852# VGND 0.366751f $ **FLOATING
C1735 a_2610_27852# VGND 0.370508f $ **FLOATING
C1736 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D VGND 0.506947f
C1737 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D VGND 0.502211f
C1738 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D VGND 0.477244f
C1739 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D VGND 0.502211f
C1740 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D VGND 0.477244f
C1741 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D VGND 0.502211f
C1742 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D VGND 0.477244f
C1743 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D VGND 0.502211f
C1744 a_21402_28204# VGND 0.405715f $ **FLOATING
C1745 a_17730_28204# VGND 0.406284f $ **FLOATING
C1746 a_16362_28204# VGND 0.406284f $ **FLOATING
C1747 a_12690_28204# VGND 0.406284f $ **FLOATING
C1748 a_11322_28204# VGND 0.406284f $ **FLOATING
C1749 a_7650_28204# VGND 0.405133f $ **FLOATING
C1750 a_6282_28204# VGND 0.404355f $ **FLOATING
C1751 a_2610_28204# VGND 0.406098f $ **FLOATING
C1752 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND 0.608956f
C1753 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND 0.741242f
C1754 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND 0.749251f
C1755 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND 0.735502f
C1756 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND 0.749251f
C1757 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND 0.735502f
C1758 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND 0.746591f
C1759 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND 0.73057f
C1760 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND 0.74895f
C1761 a_22770_28556# VGND 0.401649f $ **FLOATING
C1762 a_21402_28556# VGND 0.387558f $ **FLOATING
C1763 a_17730_28556# VGND 0.388127f $ **FLOATING
C1764 a_16362_28556# VGND 0.388127f $ **FLOATING
C1765 a_12690_28556# VGND 0.388127f $ **FLOATING
C1766 a_11322_28556# VGND 0.388127f $ **FLOATING
C1767 a_7650_28556# VGND 0.386976f $ **FLOATING
C1768 a_6282_28556# VGND 0.386198f $ **FLOATING
C1769 a_2610_28556# VGND 0.38794f $ **FLOATING
C1770 a_21402_28908# VGND 0.394283f $ **FLOATING
C1771 a_17730_28908# VGND 0.394852f $ **FLOATING
C1772 a_16362_28908# VGND 0.394852f $ **FLOATING
C1773 a_12690_28908# VGND 0.394852f $ **FLOATING
C1774 a_11322_28908# VGND 0.394852f $ **FLOATING
C1775 a_7650_28908# VGND 0.393701f $ **FLOATING
C1776 a_6282_28908# VGND 0.392923f $ **FLOATING
C1777 a_2610_28908# VGND 0.394666f $ **FLOATING
C1778 SUNSAR_SAR8B_CV_0.SARP VGND 70.097496f
C1779 a_21402_29612# VGND 0.395457f $ **FLOATING
C1780 a_17730_29612# VGND 0.396116f $ **FLOATING
C1781 a_16362_29612# VGND 0.395588f $ **FLOATING
C1782 a_12690_29612# VGND 0.396116f $ **FLOATING
C1783 a_11322_29612# VGND 0.395588f $ **FLOATING
C1784 a_7650_29612# VGND 0.394965f $ **FLOATING
C1785 a_6282_29612# VGND 0.393746f $ **FLOATING
C1786 a_2610_29612# VGND 0.395923f $ **FLOATING
C1787 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318647f
C1788 a_22770_29964# VGND 0.400512f $ **FLOATING
C1789 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND 0.103281f
C1790 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VGND 1.27143f
C1791 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND 0.100021f
C1792 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VGND 1.26503f
C1793 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND 0.100021f
C1794 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VGND 1.26391f
C1795 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND 0.100021f
C1796 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VGND 1.26503f
C1797 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND 0.100021f
C1798 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VGND 1.26391f
C1799 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND 0.100021f
C1800 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VGND 1.25938f
C1801 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND 0.100021f
C1802 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VGND 1.25329f
C1803 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND 0.100021f
C1804 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VGND 1.26407f
C1805 a_21402_30316# VGND 0.401758f $ **FLOATING
C1806 a_17730_30316# VGND 0.401074f $ **FLOATING
C1807 a_16362_30316# VGND 0.401074f $ **FLOATING
C1808 a_12690_30316# VGND 0.401074f $ **FLOATING
C1809 a_11322_30316# VGND 0.401074f $ **FLOATING
C1810 a_7650_30316# VGND 0.399923f $ **FLOATING
C1811 a_6282_30316# VGND 0.399145f $ **FLOATING
C1812 a_2610_30316# VGND 0.400881f $ **FLOATING
C1813 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND 15.315499f
C1814 a_22770_30844# VGND 0.421853f $ **FLOATING
C1815 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND 2.24318f
C1816 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND 2.22194f
C1817 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND 2.22198f
C1818 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND 2.22194f
C1819 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND 2.22198f
C1820 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND 2.20909f
C1821 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND 2.19751f
C1822 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND 2.21827f
C1823 a_21402_31196# VGND 0.4255f $ **FLOATING
C1824 a_17730_31196# VGND 0.426069f $ **FLOATING
C1825 a_16362_31196# VGND 0.426069f $ **FLOATING
C1826 a_12690_31196# VGND 0.426069f $ **FLOATING
C1827 a_11322_31196# VGND 0.426069f $ **FLOATING
C1828 a_7650_31196# VGND 0.424917f $ **FLOATING
C1829 a_6282_31196# VGND 0.42414f $ **FLOATING
C1830 a_2610_31196# VGND 0.425876f $ **FLOATING
C1831 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND 19.4783f
C1832 a_22770_31724# VGND 0.423601f $ **FLOATING
C1833 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.99939f
C1834 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.97987f
C1835 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.97901f
C1836 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.97987f
C1837 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.97901f
C1838 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.85828f
C1839 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.37577f
C1840 a_21402_32076# VGND 0.426091f $ **FLOATING
C1841 a_17730_32076# VGND 0.42666f $ **FLOATING
C1842 a_16362_32076# VGND 0.42666f $ **FLOATING
C1843 a_12690_32076# VGND 0.42666f $ **FLOATING
C1844 a_11322_32076# VGND 0.42666f $ **FLOATING
C1845 a_7650_32076# VGND 0.42666f $ **FLOATING
C1846 a_6282_32076# VGND 0.42666f $ **FLOATING
C1847 a_2610_32076# VGND 0.426468f $ **FLOATING
C1848 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND 1.55564f
C1849 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C1850 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND 3.19736f
C1851 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND 3.22974f
C1852 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND 3.22835f
C1853 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND 3.22974f
C1854 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND 3.22835f
C1855 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND 3.22678f
C1856 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND 3.22545f
C1857 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND 3.31413f
C1858 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND 2.68549f
C1859 a_21402_32956# VGND 0.426069f $ **FLOATING
C1860 a_17730_32956# VGND 0.426069f $ **FLOATING
C1861 a_16362_32956# VGND 0.426069f $ **FLOATING
C1862 a_12690_32956# VGND 0.426069f $ **FLOATING
C1863 a_11322_32956# VGND 0.426069f $ **FLOATING
C1864 a_7650_32956# VGND 0.426069f $ **FLOATING
C1865 a_6282_32956# VGND 0.426069f $ **FLOATING
C1866 a_2610_32956# VGND 0.425876f $ **FLOATING
C1867 SUNSAR_SAR8B_CV_0.XA20.XA2a.A VGND 2.85099f
C1868 a_22770_33132# VGND 0.403395f $ **FLOATING
C1869 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 3.01164f
C1870 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.01628f
C1871 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.01641f
C1872 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.01628f
C1873 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.01641f
C1874 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.54669f
C1875 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.78758f
C1876 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 12.1041f
C1877 a_21402_33836# VGND 0.426756f $ **FLOATING
C1878 a_17730_33836# VGND 0.426756f $ **FLOATING
C1879 a_16362_33836# VGND 0.426756f $ **FLOATING
C1880 a_12690_33836# VGND 0.426756f $ **FLOATING
C1881 a_11322_33836# VGND 0.426756f $ **FLOATING
C1882 a_7650_33836# VGND 0.426756f $ **FLOATING
C1883 a_6282_33836# VGND 0.426756f $ **FLOATING
C1884 a_2610_33836# VGND 0.426472f $ **FLOATING
C1885 SUNSAR_SAR8B_CV_0.SARN VGND 71.1589f
C1886 SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D VGND 0.149691f
C1887 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND 0.515385f
C1888 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C1889 SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D VGND 0.149691f
C1890 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.72791f
C1891 a_22770_34540# VGND 0.39377f $ **FLOATING
C1892 SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.D VGND 0.102f
C1893 SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D VGND 0.149691f
C1894 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 4.1719f
C1895 SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D VGND 0.149691f
C1896 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.27991f
C1897 SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.D VGND 0.102f
C1898 SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.D VGND 0.102f
C1899 SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D VGND 0.149691f
C1900 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.31299f
C1901 SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D VGND 0.149691f
C1902 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.68294f
C1903 SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.D VGND 0.102f
C1904 SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.D VGND 0.102f
C1905 SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D VGND 0.149691f
C1906 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 4.25175f
C1907 SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D VGND 0.149691f
C1908 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 10.150401f
C1909 SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.D VGND 0.102f
C1910 SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.D VGND 0.102f
C1911 SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.D VGND 0.102f
C1912 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 8.127279f
C1913 a_21402_34716# VGND 0.39476f $ **FLOATING
C1914 a_17730_34716# VGND 0.39476f $ **FLOATING
C1915 a_16362_34716# VGND 0.39476f $ **FLOATING
C1916 a_12690_34716# VGND 0.39476f $ **FLOATING
C1917 a_11322_34716# VGND 0.39476f $ **FLOATING
C1918 a_7650_34716# VGND 0.39476f $ **FLOATING
C1919 a_6282_34716# VGND 0.39476f $ **FLOATING
C1920 a_2610_34716# VGND 0.394567f $ **FLOATING
C1921 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND 4.75219f
C1922 a_22770_34892# VGND 0.394644f $ **FLOATING
C1923 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.67603f
C1924 SUNSAR_SAR8B_CV_0.XA6.ENO VGND 4.51439f
C1925 SUNSAR_SAR8B_CV_0.XA5.ENO VGND 4.46191f
C1926 SUNSAR_SAR8B_CV_0.XA4.ENO VGND 4.27708f
C1927 SUNSAR_SAR8B_CV_0.XA3.ENO VGND 4.50282f
C1928 SUNSAR_SAR8B_CV_0.XA2.ENO VGND 4.42572f
C1929 SUNSAR_SAR8B_CV_0.XA1.ENO VGND 4.44437f
C1930 SUNSAR_SAR8B_CV_0.XA0.ENO VGND 4.39222f
C1931 a_21402_35068# VGND 0.389563f $ **FLOATING
C1932 a_17730_35068# VGND 0.389563f $ **FLOATING
C1933 a_16362_35068# VGND 0.389563f $ **FLOATING
C1934 a_12690_35068# VGND 0.389563f $ **FLOATING
C1935 a_11322_35068# VGND 0.389563f $ **FLOATING
C1936 a_7650_35068# VGND 0.389563f $ **FLOATING
C1937 a_6282_35068# VGND 0.389563f $ **FLOATING
C1938 a_2610_35068# VGND 0.38937f $ **FLOATING
C1939 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND 4.54316f
C1940 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C1941 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C1942 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C1943 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C1944 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C1945 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C1946 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557214f
C1947 a_22770_35420# VGND 0.395535f $ **FLOATING
C1948 a_21402_35420# VGND 0.389041f $ **FLOATING
C1949 a_17730_35420# VGND 0.388925f $ **FLOATING
C1950 a_16362_35420# VGND 0.389297f $ **FLOATING
C1951 a_12690_35420# VGND 0.388925f $ **FLOATING
C1952 a_11322_35420# VGND 0.389297f $ **FLOATING
C1953 a_7650_35420# VGND 0.388925f $ **FLOATING
C1954 a_6282_35420# VGND 0.389297f $ **FLOATING
C1955 a_2610_35420# VGND 0.389015f $ **FLOATING
C1956 SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND 1.07685f
C1957 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND 0.112889f
C1958 SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND 1.50901f
C1959 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VGND 1.53168f
C1960 SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND 1.50964f
C1961 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND 0.112889f
C1962 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VGND 1.54335f
C1963 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND 0.112889f
C1964 SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND 1.51005f
C1965 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VGND 1.53305f
C1966 SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND 1.50964f
C1967 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND 0.112889f
C1968 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VGND 1.54335f
C1969 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND 0.112889f
C1970 SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND 1.51005f
C1971 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VGND 1.53305f
C1972 SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND 1.50964f
C1973 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND 0.112889f
C1974 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VGND 1.54335f
C1975 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND 0.112889f
C1976 SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND 1.51005f
C1977 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VGND 1.53305f
C1978 SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND 1.51935f
C1979 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND 0.112889f
C1980 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VGND 1.61753f
C1981 a_22770_35948# VGND 0.414038f $ **FLOATING
C1982 a_21402_35948# VGND 0.390722f $ **FLOATING
C1983 a_17730_35948# VGND 0.391291f $ **FLOATING
C1984 a_16362_35948# VGND 0.391291f $ **FLOATING
C1985 a_12690_35948# VGND 0.391291f $ **FLOATING
C1986 a_11322_35948# VGND 0.391291f $ **FLOATING
C1987 a_7650_35948# VGND 0.391291f $ **FLOATING
C1988 a_6282_35948# VGND 0.391291f $ **FLOATING
C1989 a_2610_35948# VGND 0.391099f $ **FLOATING
C1990 SUNSAR_SAR8B_CV_0.XA20.XA10.B VGND 0.789814f
C1991 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C1992 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C1993 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C1994 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C1995 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C1996 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C1997 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C1998 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.895311f
C1999 a_22770_36300# VGND 0.472701f $ **FLOATING
C2000 a_21402_36300# VGND 0.393831f $ **FLOATING
C2001 a_17730_36300# VGND 0.394738f $ **FLOATING
C2002 a_16362_36300# VGND 0.3944f $ **FLOATING
C2003 a_12690_36300# VGND 0.394718f $ **FLOATING
C2004 a_11322_36300# VGND 0.3944f $ **FLOATING
C2005 a_7650_36300# VGND 0.394715f $ **FLOATING
C2006 a_6282_36300# VGND 0.3944f $ **FLOATING
C2007 a_2610_36300# VGND 0.394523f $ **FLOATING
C2008 a_22770_36652# VGND 0.542245f $ **FLOATING
C2009 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND 0.881626f
C2010 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND 0.884627f
C2011 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND 0.877071f
C2012 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND 0.884604f
C2013 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND 0.877059f
C2014 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND 0.884603f
C2015 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND 0.877071f
C2016 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND 0.892649f
C2017 SUNSAR_SAR8B_CV_0.XB1.TIE_L VGND 32.9183f
C2018 a_21402_36828# VGND 0.414041f $ **FLOATING
C2019 a_17730_36828# VGND 0.413952f $ **FLOATING
C2020 a_16362_36828# VGND 0.413659f $ **FLOATING
C2021 a_12690_36828# VGND 0.413942f $ **FLOATING
C2022 a_11322_36828# VGND 0.413658f $ **FLOATING
C2023 a_7650_36828# VGND 0.413944f $ **FLOATING
C2024 a_6282_36828# VGND 0.413659f $ **FLOATING
C2025 a_2610_36828# VGND 0.413594f $ **FLOATING
C2026 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND 1.08552f
C2027 SUNSAR_SAR8B_CV_0.XA7.CEO VGND 2.06017f
C2028 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND 1.10839f
C2029 SUNSAR_SAR8B_CV_0.XA6.CEO VGND 1.45333f
C2030 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND 1.06778f
C2031 SUNSAR_SAR8B_CV_0.XA5.CEO VGND 1.71757f
C2032 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND 1.10834f
C2033 SUNSAR_SAR8B_CV_0.XA4.CEO VGND 1.52588f
C2034 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND 1.06777f
C2035 SUNSAR_SAR8B_CV_0.XA3.CEO VGND 1.71756f
C2036 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND 1.10835f
C2037 SUNSAR_SAR8B_CV_0.XA2.CEO VGND 1.52589f
C2038 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND 1.06778f
C2039 SUNSAR_SAR8B_CV_0.XA1.CEO VGND 1.71756f
C2040 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND 1.11927f
C2041 SUNSAR_SAR8B_CV_0.XA0.CEO VGND 1.53308f
C2042 a_21402_37180# VGND 0.47501f $ **FLOATING
C2043 a_17730_37180# VGND 0.474809f $ **FLOATING
C2044 a_16362_37180# VGND 0.476355f $ **FLOATING
C2045 a_12690_37180# VGND 0.47479f $ **FLOATING
C2046 a_11322_37180# VGND 0.476354f $ **FLOATING
C2047 a_7650_37180# VGND 0.474794f $ **FLOATING
C2048 a_6282_37180# VGND 0.476355f $ **FLOATING
C2049 a_2610_37180# VGND 0.474277f $ **FLOATING
C2050 a_21402_37532# VGND 0.546649f $ **FLOATING
C2051 a_17730_37532# VGND 0.548986f $ **FLOATING
C2052 a_16362_37532# VGND 0.547631f $ **FLOATING
C2053 a_12690_37532# VGND 0.548815f $ **FLOATING
C2054 a_11322_37532# VGND 0.547631f $ **FLOATING
C2055 a_7650_37532# VGND 0.548857f $ **FLOATING
C2056 a_6282_37532# VGND 0.547634f $ **FLOATING
C2057 a_2610_37532# VGND 0.546853f $ **FLOATING
C2058 a_27575_39955# VGND 0.440387f $ **FLOATING
C2059 a_27575_40307# VGND 0.408627f $ **FLOATING
C2060 tt_um_TT06_SAR_done_0.x3.MN0.S VGND 1.07773f
C2061 a_27575_40659# VGND 0.389133f $ **FLOATING
C2062 tt_um_TT06_SAR_done_0.x4.MN0.G VGND 0.822801f
C2063 a_27575_41011# VGND 0.472703f $ **FLOATING
C2064 a_27575_41363# VGND 0.532318f $ **FLOATING
C2065 a_22790_40296# VGND 0.546732f $ **FLOATING
C2066 a_21422_40296# VGND 0.54563f $ **FLOATING
C2067 a_17750_40296# VGND 0.546813f $ **FLOATING
C2068 a_16382_40296# VGND 0.547966f $ **FLOATING
C2069 a_12710_40296# VGND 0.546813f $ **FLOATING
C2070 a_11342_40296# VGND 0.547969f $ **FLOATING
C2071 a_7670_40296# VGND 0.54681f $ **FLOATING
C2072 a_6302_40296# VGND 0.547966f $ **FLOATING
C2073 a_2630_40296# VGND 0.54539f $ **FLOATING
C2074 a_22790_40648# VGND 0.492438f $ **FLOATING
C2075 a_21422_40648# VGND 0.49034f $ **FLOATING
C2076 a_17750_40648# VGND 0.492453f $ **FLOATING
C2077 a_16382_40648# VGND 0.490883f $ **FLOATING
C2078 a_12710_40648# VGND 0.492453f $ **FLOATING
C2079 a_11342_40648# VGND 0.490883f $ **FLOATING
C2080 a_7670_40648# VGND 0.492453f $ **FLOATING
C2081 a_6302_40648# VGND 0.490883f $ **FLOATING
C2082 a_2630_40648# VGND 0.492826f $ **FLOATING
C2083 tt_um_TT06_SAR_done_0.DONE VGND 22.5195f
C2084 a_22790_41000# VGND 0.388777f $ **FLOATING
C2085 a_21422_41000# VGND 0.388174f $ **FLOATING
C2086 a_17750_41000# VGND 0.388174f $ **FLOATING
C2087 a_16382_41000# VGND 0.388174f $ **FLOATING
C2088 a_12710_41000# VGND 0.388174f $ **FLOATING
C2089 a_11342_41000# VGND 0.388174f $ **FLOATING
C2090 a_7670_41000# VGND 0.388174f $ **FLOATING
C2091 a_6302_41000# VGND 0.388174f $ **FLOATING
C2092 a_2630_41000# VGND 0.388638f $ **FLOATING
C2093 a_22790_41352# VGND 0.374594f $ **FLOATING
C2094 a_21422_41352# VGND 0.393558f $ **FLOATING
C2095 a_17750_41352# VGND 0.393558f $ **FLOATING
C2096 a_16382_41352# VGND 0.393558f $ **FLOATING
C2097 a_12710_41352# VGND 0.393558f $ **FLOATING
C2098 a_11342_41352# VGND 0.393558f $ **FLOATING
C2099 a_7670_41352# VGND 0.393558f $ **FLOATING
C2100 a_6302_41352# VGND 0.393558f $ **FLOATING
C2101 a_2630_41352# VGND 0.394022f $ **FLOATING
C2102 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND 0.803097f
C2103 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND 0.107737f
C2104 SUNSAR_SAR8B_CV_0.D<0> VGND 5.87227f
C2105 SUNSAR_SAR8B_CV_0.D<1> VGND 13.789701f
C2106 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND 0.107643f
C2107 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND 0.107643f
C2108 SUNSAR_SAR8B_CV_0.D<2> VGND 12.5832f
C2109 SUNSAR_SAR8B_CV_0.D<3> VGND 11.4395f
C2110 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND 0.107643f
C2111 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND 0.107643f
C2112 SUNSAR_SAR8B_CV_0.D<4> VGND 11.8306f
C2113 SUNSAR_SAR8B_CV_0.D<5> VGND 12.7012f
C2114 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND 0.107643f
C2115 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND 0.107643f
C2116 SUNSAR_SAR8B_CV_0.D<6> VGND 12.0145f
C2117 SUNSAR_SAR8B_CV_0.D<7> VGND 17.833302f
C2118 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND 0.107643f
C2119 a_22790_41880# VGND 0.394408f $ **FLOATING
C2120 a_21422_41880# VGND 0.395138f $ **FLOATING
C2121 a_17750_41880# VGND 0.395707f $ **FLOATING
C2122 a_16382_41880# VGND 0.395707f $ **FLOATING
C2123 a_12710_41880# VGND 0.395707f $ **FLOATING
C2124 a_11342_41880# VGND 0.395707f $ **FLOATING
C2125 a_7670_41880# VGND 0.395707f $ **FLOATING
C2126 a_6302_41880# VGND 0.395707f $ **FLOATING
C2127 a_2630_41880# VGND 0.396052f $ **FLOATING
C2128 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND 1.96193f
C2129 a_22790_42408# VGND 0.410698f $ **FLOATING
C2130 a_21422_42408# VGND 0.389697f $ **FLOATING
C2131 a_17750_42408# VGND 0.390266f $ **FLOATING
C2132 a_16382_42408# VGND 0.390266f $ **FLOATING
C2133 a_12710_42408# VGND 0.390266f $ **FLOATING
C2134 a_11342_42408# VGND 0.390266f $ **FLOATING
C2135 a_7670_42408# VGND 0.390266f $ **FLOATING
C2136 a_6302_42408# VGND 0.390266f $ **FLOATING
C2137 a_2630_42408# VGND 0.390612f $ **FLOATING
C2138 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C2139 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND 1.28758f
C2140 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND 1.27933f
C2141 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND 1.27933f
C2142 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND 1.27933f
C2143 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND 1.27933f
C2144 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND 1.27933f
C2145 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND 1.27933f
C2146 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND 1.29578f
C2147 a_22790_42760# VGND 0.378208f $ **FLOATING
C2148 a_21422_42760# VGND 0.393027f $ **FLOATING
C2149 a_17750_42760# VGND 0.393596f $ **FLOATING
C2150 a_16382_42760# VGND 0.393596f $ **FLOATING
C2151 a_12710_42760# VGND 0.393596f $ **FLOATING
C2152 a_11342_42760# VGND 0.393596f $ **FLOATING
C2153 a_7670_42760# VGND 0.393596f $ **FLOATING
C2154 a_6302_42760# VGND 0.393596f $ **FLOATING
C2155 a_2630_42760# VGND 0.393942f $ **FLOATING
C2156 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 24.6885f
C2157 SUNSAR_SAR8B_CV_0.EN VGND 10.9728f
C2158 a_22790_43112# VGND 0.388427f $ **FLOATING
C2159 SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND 1.29446f
C2160 SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND 1.29655f
C2161 SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND 1.29655f
C2162 SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND 1.29655f
C2163 SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND 1.29655f
C2164 SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND 1.29655f
C2165 SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND 1.29655f
C2166 SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND 1.29893f
C2167 SUNSAR_CAPT8B_CV_0.XA4.Y VGND 2.38038f
C2168 a_21422_43288# VGND 0.394124f $ **FLOATING
C2169 a_17750_43288# VGND 0.394693f $ **FLOATING
C2170 a_16382_43288# VGND 0.394693f $ **FLOATING
C2171 a_12710_43288# VGND 0.394693f $ **FLOATING
C2172 a_11342_43288# VGND 0.394693f $ **FLOATING
C2173 a_7670_43288# VGND 0.394693f $ **FLOATING
C2174 a_6302_43288# VGND 0.394693f $ **FLOATING
C2175 a_2630_43288# VGND 0.395039f $ **FLOATING
C2176 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND 0.103608f
C2177 SUNSAR_CAPT8B_CV_0.XA3.Y VGND 1.65375f
C2178 a_22790_43640# VGND 0.387806f $ **FLOATING
C2179 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND 0.112889f
C2180 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND 2.60322f
C2181 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VGND 1.69058f
C2182 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND 0.112889f
C2183 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VGND 1.69315f
C2184 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND 2.58593f
C2185 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND 0.112889f
C2186 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND 2.63669f
C2187 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VGND 1.69315f
C2188 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND 0.112889f
C2189 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VGND 1.69315f
C2190 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND 2.63655f
C2191 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND 0.112889f
C2192 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND 2.59274f
C2193 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VGND 1.69797f
C2194 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND 0.112889f
C2195 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VGND 1.69797f
C2196 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND 2.5926f
C2197 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND 0.112889f
C2198 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND 2.6374f
C2199 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VGND 1.69797f
C2200 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND 0.112889f
C2201 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VGND 1.69726f
C2202 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND 2.70316f
C2203 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.88269f
C2204 a_21422_43816# VGND 0.390629f $ **FLOATING
C2205 a_17750_43816# VGND 0.391198f $ **FLOATING
C2206 a_16382_43816# VGND 0.391198f $ **FLOATING
C2207 a_12710_43816# VGND 0.391198f $ **FLOATING
C2208 a_11342_43816# VGND 0.391198f $ **FLOATING
C2209 a_7670_43816# VGND 0.391198f $ **FLOATING
C2210 a_6302_43816# VGND 0.391198f $ **FLOATING
C2211 a_2630_43816# VGND 0.391544f $ **FLOATING
C2212 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 26.5938f
C2213 a_22790_43992# VGND 0.384235f $ **FLOATING
C2214 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.23582f
C2215 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.23517f
C2216 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.23517f
C2217 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.23517f
C2218 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26123f
C2219 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C2220 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C2221 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C2222 SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND 0.5774f
C2223 a_21422_44168# VGND 0.425534f $ **FLOATING
C2224 a_17750_44168# VGND 0.425449f $ **FLOATING
C2225 a_16382_44168# VGND 0.425864f $ **FLOATING
C2226 a_12710_44168# VGND 0.425449f $ **FLOATING
C2227 a_11342_44168# VGND 0.425864f $ **FLOATING
C2228 a_7670_44168# VGND 0.425449f $ **FLOATING
C2229 a_6302_44168# VGND 0.425864f $ **FLOATING
C2230 a_2630_44168# VGND 0.426034f $ **FLOATING
C2231 TIE_L VGND 6.36945f
C2232 a_22790_44344# VGND 0.423601f $ **FLOATING
.ends

