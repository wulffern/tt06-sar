magic
tech sky130B
magscale 1 2
timestamp 1708687947
<< locali >>
rect 6142 44434 6202 44440
rect 6142 44386 6148 44434
rect 6196 44386 6202 44434
rect 3398 44082 3458 44230
rect 6142 44166 6202 44386
rect 16220 44390 16280 44396
rect 16220 44342 16226 44390
rect 16274 44342 16280 44390
rect 3398 44034 3404 44082
rect 3452 44034 3458 44082
rect 8474 44090 8534 44230
rect 8474 44042 8480 44090
rect 8528 44042 8534 44090
rect 10896 44118 10956 44226
rect 10896 44070 10902 44118
rect 10950 44070 10956 44118
rect 10896 44064 10956 44070
rect 13498 44110 13558 44240
rect 16220 44172 16280 44342
rect 13498 44062 13504 44110
rect 13552 44062 13558 44110
rect 13498 44056 13558 44062
rect 18692 44076 18752 44228
rect 8474 44036 8534 44042
rect 3398 44028 3458 44034
rect 18692 44028 18698 44076
rect 18746 44028 18752 44076
rect 18692 44022 18752 44028
rect 21298 44068 21361 44243
rect 21298 44017 21304 44068
rect 21355 44017 21361 44068
rect 21298 44011 21361 44017
rect 23318 44006 26726 44074
rect 23318 43650 23386 44006
rect 22646 43022 22886 43090
rect 22646 41848 22714 43022
rect 23840 42760 24252 42828
rect 22916 42530 22984 42736
rect 22916 42462 23270 42530
rect 23202 42408 23270 42462
rect 23754 42408 24252 42476
rect 22646 41780 22966 41848
rect 22898 41650 22966 41780
rect 22898 41582 23270 41650
rect 23202 41528 23270 41582
rect 2641 41349 2711 41501
rect 2641 41291 2647 41349
rect 2705 41291 2711 41349
rect 6860 41374 6928 41502
rect 6860 41318 6866 41374
rect 6922 41318 6928 41374
rect 7772 41380 7840 41498
rect 7772 41324 7778 41380
rect 7834 41324 7840 41380
rect 7772 41318 7840 41324
rect 6860 41312 6928 41318
rect 2641 41285 2711 41291
rect 11918 41300 11986 41506
rect 11918 41244 11924 41300
rect 11980 41244 11986 41300
rect 12766 41316 12834 41496
rect 12766 41260 12772 41316
rect 12828 41260 12834 41316
rect 16952 41360 17020 41500
rect 16952 41304 16958 41360
rect 17014 41304 17020 41360
rect 16952 41298 17020 41304
rect 17816 41326 17884 41506
rect 17816 41270 17822 41326
rect 17878 41270 17884 41326
rect 21968 41340 22036 41494
rect 21968 41284 21974 41340
rect 22030 41284 22036 41340
rect 21968 41278 22036 41284
rect 17816 41264 17884 41270
rect 12766 41254 12834 41260
rect 22764 41246 22824 41344
rect 11918 41238 11986 41244
rect 22644 41240 22824 41246
rect 22644 41192 22650 41240
rect 22698 41192 22824 41240
rect 22644 41186 22824 41192
rect 22732 40734 22736 40794
rect 22796 40734 22880 40794
rect 2686 40492 2754 40628
rect 6862 40470 6930 40628
rect 7718 40516 7786 40628
rect 11910 40458 11978 40628
rect 12764 40516 12832 40628
rect 16948 40470 17016 40628
rect 17808 40502 17876 40628
rect 21986 40408 22054 40628
rect 22820 40576 22880 40734
rect 12390 38800 12574 39710
rect 26658 39502 26726 44006
rect 22570 38738 22638 38750
rect 22570 38682 22578 38738
rect 22634 38682 22638 38738
rect 22570 38634 22638 38682
rect 2686 38632 24980 38634
rect 2686 38628 12770 38632
rect 2686 38572 2692 38628
rect 2748 38626 12770 38628
rect 2748 38572 6868 38626
rect 2686 38570 6868 38572
rect 6924 38570 7724 38626
rect 7780 38570 11916 38626
rect 11972 38576 12770 38626
rect 12826 38630 24980 38632
rect 12826 38626 17814 38630
rect 12826 38576 16954 38626
rect 11972 38570 16954 38576
rect 17010 38574 17814 38626
rect 17870 38624 24980 38630
rect 17870 38574 21992 38624
rect 17010 38570 21992 38574
rect 2686 38568 21992 38570
rect 22048 38568 24980 38624
rect 2686 38566 24980 38568
<< viali >>
rect 6148 44386 6196 44434
rect 16226 44342 16274 44390
rect 3404 44034 3452 44082
rect 8480 44042 8528 44090
rect 10902 44070 10950 44118
rect 13504 44062 13552 44110
rect 18698 44028 18746 44076
rect 21304 44017 21355 44068
rect 24252 42760 24320 42828
rect 24252 42408 24320 42476
rect 2647 41291 2705 41349
rect 6866 41318 6922 41374
rect 7778 41324 7834 41380
rect 11924 41244 11980 41300
rect 12772 41260 12828 41316
rect 16958 41304 17014 41360
rect 17822 41270 17878 41326
rect 21974 41284 22030 41340
rect 22650 41192 22698 41240
rect 22736 40734 22796 40794
rect 2686 40424 2754 40492
rect 6862 40402 6930 40470
rect 7718 40448 7786 40516
rect 11910 40390 11978 40458
rect 12764 40448 12832 40516
rect 16948 40402 17016 40470
rect 17808 40434 17876 40502
rect 21986 40340 22054 40408
rect 22578 38682 22634 38738
rect 2692 38572 2748 38628
rect 6868 38570 6924 38626
rect 7724 38570 7780 38626
rect 11916 38570 11972 38626
rect 12770 38576 12826 38632
rect 16954 38570 17010 38626
rect 17814 38574 17870 38630
rect 21992 38568 22048 38624
<< metal1 >>
rect 13034 44440 13094 44446
rect 6136 44434 13034 44440
rect 6136 44386 6148 44434
rect 6196 44386 13034 44434
rect 6136 44380 13034 44386
rect 13034 44374 13094 44380
rect 16060 44336 16066 44396
rect 16126 44390 16286 44396
rect 16126 44342 16226 44390
rect 16274 44342 16286 44390
rect 16126 44336 16286 44342
rect 11218 44124 11278 44130
rect 10890 44118 11218 44124
rect 8468 44090 8710 44096
rect 3392 44082 3654 44088
rect 3392 44034 3404 44082
rect 3452 44034 3654 44082
rect 3392 44028 3654 44034
rect 3714 44028 3720 44088
rect 8468 44042 8480 44090
rect 8528 44042 8710 44090
rect 8468 44036 8710 44042
rect 8770 44036 8776 44096
rect 10890 44070 10902 44118
rect 10950 44070 11218 44118
rect 10890 44064 11218 44070
rect 11218 44058 11278 44064
rect 13492 44110 13718 44116
rect 13492 44062 13504 44110
rect 13552 44062 13718 44110
rect 13492 44056 13718 44062
rect 13778 44056 13784 44116
rect 18450 44022 18456 44082
rect 18516 44076 18758 44082
rect 18516 44028 18698 44076
rect 18746 44028 18758 44076
rect 18516 44022 18758 44028
rect 21141 44074 21204 44080
rect 21298 44074 21361 44080
rect 21204 44068 21361 44074
rect 21204 44017 21304 44068
rect 21355 44017 21361 44068
rect 21204 44011 21361 44017
rect 21141 44005 21204 44011
rect 21298 44005 21361 44011
rect 24246 42828 24326 42840
rect 24474 42828 24542 42834
rect 24246 42760 24252 42828
rect 24320 42760 24474 42828
rect 24246 42748 24326 42760
rect 24474 42754 24542 42760
rect 25596 42828 25664 42834
rect 24246 42476 24326 42488
rect 25344 42476 25412 42482
rect 24246 42408 24252 42476
rect 24320 42408 24336 42476
rect 24404 42408 24410 42476
rect 25342 42408 25344 42460
rect 24246 42396 24326 42408
rect 25342 42402 25412 42408
rect 6860 41374 6928 41386
rect 2641 41349 2711 41361
rect 2641 41291 2647 41349
rect 2705 41291 2711 41349
rect 2641 41145 2711 41291
rect 6860 41318 6866 41374
rect 6922 41318 6928 41374
rect 6860 41238 6928 41318
rect 7772 41380 7840 41392
rect 7772 41324 7778 41380
rect 7834 41324 7840 41380
rect 16952 41360 17020 41372
rect 7772 41260 7840 41324
rect 12766 41316 12834 41328
rect 11918 41300 11986 41312
rect 6854 41170 6860 41238
rect 6928 41170 6934 41238
rect 7086 41156 7590 41224
rect 7766 41192 7772 41260
rect 7840 41192 7846 41260
rect 9582 41174 9650 41290
rect 11918 41244 11924 41300
rect 11980 41244 11986 41300
rect 11918 41174 11986 41244
rect 12766 41260 12772 41316
rect 12828 41260 12834 41316
rect 12132 41180 12630 41222
rect 2635 41075 2641 41145
rect 2711 41075 2717 41145
rect 9582 41106 10084 41174
rect 11912 41106 11918 41174
rect 11986 41106 11992 41174
rect 12102 41154 12630 41180
rect 12766 41164 12834 41260
rect 16952 41304 16958 41360
rect 17014 41304 17020 41360
rect 21968 41340 22036 41352
rect 16952 41216 17020 41304
rect 17816 41326 17884 41338
rect 17816 41270 17822 41326
rect 17878 41270 17884 41326
rect 2488 40736 2494 40804
rect 2562 40736 2568 40804
rect 7062 40762 7130 41036
rect 7062 40688 7130 40694
rect 9582 40756 9650 41106
rect 12102 40762 12170 41154
rect 12760 41096 12766 41164
rect 12834 41096 12840 41164
rect 16946 41148 16952 41216
rect 17020 41148 17026 41216
rect 12102 40688 12170 40694
rect 14622 41082 14690 41148
rect 17142 41100 17210 41212
rect 17816 41194 17884 41270
rect 21968 41284 21974 41340
rect 22030 41284 22036 41340
rect 17810 41126 17816 41194
rect 17884 41126 17890 41194
rect 21968 41186 22036 41284
rect 14622 41014 15150 41082
rect 17142 41032 17662 41100
rect 19662 41078 19730 41128
rect 21962 41118 21968 41186
rect 22036 41118 22042 41186
rect 22182 41090 22250 41712
rect 22638 41268 22644 41328
rect 22704 41268 22710 41328
rect 22644 41240 22704 41268
rect 22644 41192 22650 41240
rect 22698 41192 22704 41240
rect 22644 41180 22704 41192
rect 14622 40754 14690 41014
rect 9582 40682 9650 40688
rect 14622 40680 14690 40686
rect 17142 40756 17210 41032
rect 19662 41010 20144 41078
rect 19662 40762 19730 41010
rect 19662 40688 19730 40694
rect 22182 40758 22250 41022
rect 22730 40794 22802 40806
rect 22588 40734 22594 40794
rect 22654 40734 22736 40794
rect 22796 40734 22802 40794
rect 22730 40722 22802 40734
rect 17142 40682 17210 40688
rect 22182 40684 22250 40690
rect 7706 40516 7798 40522
rect 2674 40492 2766 40498
rect 2674 40424 2686 40492
rect 2754 40424 2766 40492
rect 2674 40418 2766 40424
rect 6850 40470 6942 40476
rect 2686 38628 2754 40418
rect 6850 40402 6862 40470
rect 6930 40402 6942 40470
rect 7706 40448 7718 40516
rect 7786 40448 7798 40516
rect 12752 40516 12844 40522
rect 7706 40442 7798 40448
rect 11898 40458 11990 40464
rect 6850 40396 6942 40402
rect 2686 38572 2692 38628
rect 2748 38572 2754 38628
rect 2686 38560 2754 38572
rect 6862 38626 6930 40396
rect 6862 38570 6868 38626
rect 6924 38570 6930 38626
rect 6862 38558 6930 38570
rect 7718 38626 7786 40442
rect 11898 40390 11910 40458
rect 11978 40390 11990 40458
rect 12752 40448 12764 40516
rect 12832 40448 12844 40516
rect 17796 40502 17888 40508
rect 12752 40442 12844 40448
rect 16936 40470 17028 40476
rect 11898 40384 11990 40390
rect 7718 38570 7724 38626
rect 7780 38570 7786 38626
rect 7718 38558 7786 38570
rect 11910 38626 11978 40384
rect 11910 38570 11916 38626
rect 11972 38570 11978 38626
rect 11910 38558 11978 38570
rect 12764 38632 12832 40442
rect 16936 40402 16948 40470
rect 17016 40402 17028 40470
rect 17796 40434 17808 40502
rect 17876 40434 17888 40502
rect 17796 40428 17888 40434
rect 16936 40396 17028 40402
rect 12764 38576 12770 38632
rect 12826 38576 12832 38632
rect 12764 38564 12832 38576
rect 16948 38626 17016 40396
rect 16948 38570 16954 38626
rect 17010 38570 17016 38626
rect 16948 38558 17016 38570
rect 17808 38630 17876 40428
rect 21974 40408 22066 40414
rect 21974 40340 21986 40408
rect 22054 40340 22066 40408
rect 21974 40334 22066 40340
rect 17808 38574 17814 38630
rect 17870 38574 17876 38630
rect 17808 38562 17876 38574
rect 21986 38624 22054 40334
rect 21986 38568 21992 38624
rect 22048 38568 22054 38624
rect 21986 38556 22054 38568
rect 22572 38738 22640 38750
rect 22572 38682 22578 38738
rect 22634 38682 22640 38738
rect 22572 38546 22640 38682
rect 22566 38478 22572 38546
rect 22640 38478 22646 38546
rect 25342 34112 25410 42402
rect 25596 39612 25664 42760
rect 25596 39388 25684 39612
rect 25590 39272 25702 39388
rect 25616 37946 25684 39272
rect 25616 37872 25684 37878
rect 25342 34038 25410 34044
<< via1 >>
rect 13034 44380 13094 44440
rect 16066 44336 16126 44396
rect 3654 44028 3714 44088
rect 8710 44036 8770 44096
rect 11218 44064 11278 44124
rect 13718 44056 13778 44116
rect 18456 44022 18516 44082
rect 21141 44011 21204 44074
rect 24474 42760 24542 42828
rect 25596 42760 25664 42828
rect 24336 42408 24404 42476
rect 25344 42408 25412 42476
rect 6860 41170 6928 41238
rect 7772 41192 7840 41260
rect 2641 41075 2711 41145
rect 11918 41106 11986 41174
rect 2494 40736 2562 40804
rect 7062 40694 7130 40762
rect 9582 40688 9650 40756
rect 12766 41096 12834 41164
rect 16952 41148 17020 41216
rect 12102 40694 12170 40762
rect 17816 41126 17884 41194
rect 21968 41118 22036 41186
rect 22644 41268 22704 41328
rect 14622 40686 14690 40754
rect 17142 40688 17210 40756
rect 22182 41022 22250 41090
rect 19662 40694 19730 40762
rect 22182 40690 22250 40758
rect 22594 40734 22654 40794
rect 22572 38478 22640 38546
rect 25616 37878 25684 37946
rect 25342 34044 25410 34112
<< metal2 >>
rect 21144 44847 21200 44852
rect 21141 44843 21204 44847
rect 21141 44787 21144 44843
rect 21200 44787 21204 44843
rect 8712 44776 8768 44783
rect 8710 44774 8770 44776
rect 8710 44718 8712 44774
rect 8768 44718 8770 44774
rect 3656 44440 3712 44447
rect 3654 44438 3714 44440
rect 3654 44382 3656 44438
rect 3712 44382 3714 44438
rect 3654 44088 3714 44382
rect 8710 44096 8770 44718
rect 18458 44676 18514 44683
rect 18456 44674 18516 44676
rect 18456 44618 18458 44674
rect 18514 44618 18516 44674
rect 11220 44608 11276 44615
rect 11218 44606 11278 44608
rect 11218 44550 11220 44606
rect 11276 44550 11278 44606
rect 11218 44124 11278 44550
rect 13178 44440 13234 44447
rect 13028 44380 13034 44440
rect 13094 44438 13236 44440
rect 13094 44382 13178 44438
rect 13234 44382 13236 44438
rect 13718 44404 13778 44406
rect 13094 44380 13236 44382
rect 13178 44373 13234 44380
rect 13711 44348 13720 44404
rect 13776 44348 13785 44404
rect 16066 44396 16126 44402
rect 11212 44064 11218 44124
rect 11278 44064 11284 44124
rect 13718 44116 13778 44348
rect 16066 44126 16126 44336
rect 16066 44070 16068 44126
rect 16124 44070 16126 44126
rect 16066 44068 16126 44070
rect 18456 44082 18516 44618
rect 16068 44061 16124 44068
rect 13718 44050 13778 44056
rect 8710 44030 8770 44036
rect 3654 44022 3714 44028
rect 21141 44074 21204 44787
rect 18456 44016 18516 44022
rect 21135 44011 21141 44074
rect 21204 44011 21210 44074
rect 24468 42760 24474 42828
rect 24542 42760 25596 42828
rect 25664 42760 25670 42828
rect 24336 42476 24404 42482
rect 24404 42408 25344 42476
rect 25412 42408 25418 42476
rect 24336 42402 24404 42408
rect 22644 41446 22704 41448
rect 22637 41390 22646 41446
rect 22702 41390 22711 41446
rect 22644 41328 22704 41390
rect 7772 41260 7840 41266
rect 22644 41262 22704 41268
rect 6860 41238 6928 41244
rect 2641 41145 2711 41151
rect 2641 41004 2711 41075
rect 6860 41061 6928 41170
rect 7772 41137 7840 41192
rect 16952 41216 17020 41222
rect 11918 41174 11986 41180
rect 7768 41079 7777 41137
rect 7835 41079 7844 41137
rect 7772 41074 7840 41079
rect 2637 40944 2646 41004
rect 2706 40944 2715 41004
rect 6856 41003 6865 41061
rect 6923 41003 6932 41061
rect 11918 41033 11986 41106
rect 12766 41164 12834 41170
rect 6860 40998 6928 41003
rect 11914 40975 11923 41033
rect 11981 40975 11990 41033
rect 12766 41015 12834 41096
rect 16952 41017 17020 41148
rect 17816 41194 17884 41200
rect 17816 41049 17884 41126
rect 21968 41186 22036 41192
rect 11918 40970 11986 40975
rect 12762 40957 12771 41015
rect 12829 40957 12838 41015
rect 16948 40959 16957 41017
rect 17015 40959 17024 41017
rect 17812 40991 17821 41049
rect 17879 40991 17888 41049
rect 21968 41007 22036 41118
rect 22176 41022 22182 41090
rect 22250 41022 23544 41090
rect 17816 40986 17884 40991
rect 12766 40952 12834 40957
rect 16952 40954 17020 40959
rect 21964 40949 21973 41007
rect 22031 40949 22040 41007
rect 21968 40944 22036 40949
rect 2641 40939 2711 40944
rect 22594 40892 22654 40901
rect 2494 40804 2562 40810
rect 22594 40794 22654 40832
rect 7056 40756 7062 40762
rect 2562 40736 7062 40756
rect 2494 40694 7062 40736
rect 7130 40756 7136 40762
rect 12096 40756 12102 40762
rect 7130 40694 9582 40756
rect 2494 40688 9582 40694
rect 9650 40694 12102 40756
rect 12170 40756 12176 40762
rect 19656 40756 19662 40762
rect 12170 40754 17142 40756
rect 12170 40694 14622 40754
rect 9650 40688 14622 40694
rect 14616 40686 14622 40688
rect 14690 40688 17142 40754
rect 17210 40694 19662 40756
rect 19730 40756 19736 40762
rect 22176 40756 22182 40758
rect 19730 40694 22182 40756
rect 17210 40690 22182 40694
rect 22250 40756 22256 40758
rect 22250 40690 22376 40756
rect 22594 40728 22654 40734
rect 17210 40688 22376 40690
rect 14690 40686 14696 40688
rect 6211 39881 6860 39886
rect 6207 39823 6216 39881
rect 6274 39823 6860 39881
rect 6211 39818 6860 39823
rect 6928 39818 6937 39886
rect 11251 39869 11918 39874
rect 7763 39782 7772 39850
rect 7840 39845 8440 39850
rect 7840 39787 8377 39845
rect 8435 39787 8444 39845
rect 11247 39811 11256 39869
rect 11314 39811 11918 39869
rect 11251 39806 11918 39811
rect 11986 39806 11995 39874
rect 16291 39851 16952 39856
rect 7840 39782 8440 39787
rect 12757 39782 12766 39850
rect 12834 39845 13480 39850
rect 12834 39787 13417 39845
rect 13475 39787 13484 39845
rect 16287 39793 16296 39851
rect 16354 39793 16952 39851
rect 16291 39788 16952 39793
rect 17020 39788 17029 39856
rect 17807 39802 17816 39870
rect 17884 39865 18520 39870
rect 17884 39807 18457 39865
rect 18515 39807 18524 39865
rect 21331 39859 21968 39864
rect 17884 39802 18520 39807
rect 21327 39801 21336 39859
rect 21394 39801 21968 39859
rect 21331 39796 21968 39801
rect 22036 39796 22045 39864
rect 12834 39782 13480 39787
rect 22572 38546 22640 38552
rect 22572 38445 22640 38478
rect 22568 38387 22577 38445
rect 22635 38387 22644 38445
rect 22572 38382 22640 38387
rect 20510 37941 25616 37946
rect 20506 37883 20515 37941
rect 20573 37883 25616 37941
rect 20510 37878 25616 37883
rect 25684 37878 25690 37946
rect 22572 35824 22640 35833
rect 22572 35747 22640 35756
rect 22044 34044 25342 34112
rect 25410 34044 25416 34112
rect 20114 30124 20510 30192
rect 20578 30124 20587 30192
rect 12694 413 12814 2926
rect 14498 695 14618 2932
rect 14498 585 14503 695
rect 14613 585 14618 695
rect 14498 580 14618 585
rect 14503 576 14613 580
rect 12690 303 12699 413
rect 12809 303 12818 413
rect 12694 298 12814 303
<< via2 >>
rect 21144 44787 21200 44843
rect 8712 44718 8768 44774
rect 3656 44382 3712 44438
rect 18458 44618 18514 44674
rect 11220 44550 11276 44606
rect 13178 44382 13234 44438
rect 13720 44348 13776 44404
rect 16068 44070 16124 44126
rect 22646 41390 22702 41446
rect 7777 41079 7835 41137
rect 2646 40944 2706 41004
rect 6865 41003 6923 41061
rect 11923 40975 11981 41033
rect 12771 40957 12829 41015
rect 16957 40959 17015 41017
rect 17821 40991 17879 41049
rect 21973 40949 22031 41007
rect 22594 40832 22654 40892
rect 6216 39823 6274 39881
rect 6860 39818 6928 39886
rect 7772 39782 7840 39850
rect 8377 39787 8435 39845
rect 11256 39811 11314 39869
rect 11918 39806 11986 39874
rect 12766 39782 12834 39850
rect 13417 39787 13475 39845
rect 16296 39793 16354 39851
rect 16952 39788 17020 39856
rect 17816 39802 17884 39870
rect 18457 39807 18515 39865
rect 21336 39801 21394 39859
rect 21968 39796 22036 39864
rect 22577 38387 22635 38445
rect 20515 37883 20573 37941
rect 22572 35756 22640 35824
rect 20510 30124 20578 30192
rect 14503 585 14613 695
rect 12699 303 12809 413
<< metal3 >>
rect 21139 44846 21205 44848
rect 17718 44782 17724 44846
rect 17788 44844 17794 44846
rect 18501 44844 21205 44846
rect 17788 44843 21205 44844
rect 17788 44787 21144 44843
rect 21200 44787 21205 44843
rect 17788 44784 21205 44787
rect 17788 44782 17794 44784
rect 18501 44783 21205 44784
rect 21139 44782 21205 44783
rect 8707 44776 8773 44779
rect 14038 44776 14044 44778
rect 8707 44774 14044 44776
rect 8707 44718 8712 44774
rect 8768 44718 14044 44774
rect 8707 44716 14044 44718
rect 8707 44713 8773 44716
rect 14038 44714 14044 44716
rect 14108 44714 14114 44778
rect 11215 44608 11281 44611
rect 14780 44610 14844 44616
rect 16982 44614 16988 44678
rect 17052 44676 17058 44678
rect 18453 44676 18519 44679
rect 17052 44674 18519 44676
rect 17052 44618 18458 44674
rect 18514 44618 18519 44674
rect 22636 44668 22642 44732
rect 22706 44730 22712 44732
rect 30966 44730 30972 44732
rect 22706 44670 30972 44730
rect 22706 44668 22712 44670
rect 30966 44668 30972 44670
rect 31036 44668 31042 44732
rect 17052 44616 18519 44618
rect 17052 44614 17058 44616
rect 18453 44613 18519 44616
rect 11215 44606 14780 44608
rect 11215 44550 11220 44606
rect 11276 44550 14780 44606
rect 11215 44548 14780 44550
rect 11215 44545 11281 44548
rect 14780 44540 14844 44546
rect 15510 44498 15516 44500
rect 13708 44463 13802 44476
rect 14956 44463 15516 44498
rect 3651 44440 3717 44443
rect 12566 44440 12572 44442
rect 3651 44438 12572 44440
rect 3651 44382 3656 44438
rect 3712 44382 12572 44438
rect 3651 44380 12572 44382
rect 3651 44377 3717 44380
rect 12566 44378 12572 44380
rect 12636 44378 12642 44442
rect 13173 44440 13239 44443
rect 13302 44440 13308 44442
rect 13173 44438 13308 44440
rect 13173 44382 13178 44438
rect 13234 44382 13308 44438
rect 13173 44380 13308 44382
rect 13173 44377 13239 44380
rect 13302 44378 13308 44380
rect 13372 44378 13378 44442
rect 13708 44438 15516 44463
rect 13708 44404 15017 44438
rect 15510 44436 15516 44438
rect 15580 44436 15586 44500
rect 22448 44462 22454 44526
rect 22518 44524 22524 44526
rect 29494 44524 29500 44526
rect 22518 44464 29500 44524
rect 22518 44462 22524 44464
rect 29494 44462 29500 44464
rect 29564 44462 29570 44526
rect 13708 44348 13720 44404
rect 13776 44402 15017 44404
rect 13776 44348 13802 44402
rect 13708 44340 13802 44348
rect 16063 44128 16129 44131
rect 16246 44128 16252 44130
rect 16063 44126 16252 44128
rect 16063 44070 16068 44126
rect 16124 44070 16252 44126
rect 16063 44068 16252 44070
rect 16063 44065 16129 44068
rect 16246 44066 16252 44068
rect 16316 44066 16322 44130
rect 22636 41558 22720 41568
rect 2641 41004 2711 41009
rect 2641 40944 2646 41004
rect 2706 40944 2711 41004
rect 2641 29275 2711 40944
rect 3042 37740 3226 41532
rect 22636 41494 22642 41558
rect 22706 41494 22720 41558
rect 22636 41446 22720 41494
rect 22636 41390 22646 41446
rect 22702 41390 22720 41446
rect 22636 41384 22720 41390
rect 7772 41137 7840 41142
rect 3834 39424 4018 41084
rect 7772 41079 7777 41137
rect 7835 41079 7840 41137
rect 6860 41061 6928 41066
rect 6860 41003 6865 41061
rect 6923 41003 6928 41061
rect 4552 39424 5074 39452
rect 5594 39424 5778 40752
rect 3834 39423 5778 39424
rect 3834 39125 4711 39423
rect 5009 39125 5778 39423
rect 3834 39124 5778 39125
rect 3834 37818 4018 39124
rect 4552 39102 5074 39124
rect 5594 38304 5778 39124
rect 6211 39881 6279 39886
rect 6211 39823 6216 39881
rect 6274 39823 6279 39881
rect 6211 30970 6279 39823
rect 6386 37728 6570 40610
rect 6860 39891 6928 41003
rect 6855 39886 6933 39891
rect 6855 39818 6860 39886
rect 6928 39818 6933 39886
rect 7772 39855 7840 41079
rect 17816 41049 17884 41054
rect 11918 41033 11986 41038
rect 11918 40975 11923 41033
rect 11981 40975 11986 41033
rect 6855 39813 6933 39818
rect 7767 39850 7845 39855
rect 7767 39782 7772 39850
rect 7840 39782 7845 39850
rect 7767 39777 7845 39782
rect 8082 37804 8266 40650
rect 8372 39845 8440 39850
rect 8372 39787 8377 39845
rect 8435 39787 8440 39845
rect 8372 27636 8440 39787
rect 8874 39424 9058 40598
rect 10634 39429 10818 40904
rect 11251 39869 11319 39874
rect 11251 39811 11256 39869
rect 11314 39811 11319 39869
rect 10579 39424 10877 39429
rect 8856 39423 10878 39424
rect 8856 39125 10579 39423
rect 10877 39125 10878 39423
rect 8856 39124 10878 39125
rect 8874 37676 9058 39124
rect 10579 39119 10877 39124
rect 10634 38418 10818 39119
rect 11251 28232 11319 39811
rect 11426 38382 11610 40662
rect 11918 39879 11986 40975
rect 12766 41015 12834 41020
rect 12766 40957 12771 41015
rect 12829 40957 12834 41015
rect 11913 39874 11991 39879
rect 11913 39806 11918 39874
rect 11986 39806 11991 39874
rect 12766 39855 12834 40957
rect 16952 41017 17020 41022
rect 16952 40959 16957 41017
rect 17015 40959 17020 41017
rect 11913 39801 11991 39806
rect 12761 39850 12839 39855
rect 12761 39782 12766 39850
rect 12834 39782 12839 39850
rect 12761 39777 12839 39782
rect 12301 38382 12599 38387
rect 13122 38382 13306 40444
rect 11426 38381 13306 38382
rect 11426 38083 12301 38381
rect 12599 38083 13306 38381
rect 11426 38082 13306 38083
rect 11426 37740 11610 38082
rect 12301 38077 12599 38082
rect 13122 37766 13306 38082
rect 13412 39845 13480 39850
rect 13412 39787 13417 39845
rect 13475 39787 13480 39845
rect 13412 26386 13480 39787
rect 13914 39429 14098 40598
rect 13851 39424 14149 39429
rect 15674 39424 15858 40458
rect 13850 39423 15858 39424
rect 13850 39125 13851 39423
rect 14149 39125 15858 39423
rect 13850 39124 15858 39125
rect 13851 39119 14149 39124
rect 13914 37818 14098 39119
rect 15674 38368 15858 39124
rect 16291 39851 16359 39856
rect 16291 39793 16296 39851
rect 16354 39793 16359 39851
rect 16291 29204 16359 39793
rect 16466 37780 16650 40700
rect 16952 39861 17020 40959
rect 17816 40991 17821 41049
rect 17879 40991 17884 41049
rect 17816 39875 17884 40991
rect 21968 41007 22036 41012
rect 21968 40949 21973 41007
rect 22031 40949 22036 41007
rect 17811 39870 17889 39875
rect 16947 39856 17025 39861
rect 16947 39788 16952 39856
rect 17020 39788 17025 39856
rect 17811 39802 17816 39870
rect 17884 39802 17889 39870
rect 17811 39797 17889 39802
rect 16947 39783 17025 39788
rect 18162 37766 18346 40636
rect 18452 39865 18520 39870
rect 18452 39807 18457 39865
rect 18515 39807 18520 39865
rect 18452 26436 18520 39807
rect 18954 39424 19138 40662
rect 19875 39424 20173 39429
rect 20714 39424 20898 40586
rect 18954 39423 20898 39424
rect 18954 39125 19875 39423
rect 20173 39125 20898 39423
rect 18954 39124 20898 39125
rect 18954 37754 19138 39124
rect 19875 39119 20173 39124
rect 20714 38482 20898 39124
rect 21331 39859 21399 39864
rect 21331 39801 21336 39859
rect 21394 39801 21399 39859
rect 20510 37941 20578 38358
rect 20510 37883 20515 37941
rect 20573 37883 20578 37941
rect 20510 30197 20578 37883
rect 21331 31422 21399 39801
rect 21506 37716 21690 40546
rect 21968 39869 22036 40949
rect 22456 40894 22520 40900
rect 22589 40892 22659 40897
rect 22520 40832 22594 40892
rect 22654 40832 22659 40892
rect 23202 40880 23386 40892
rect 22456 40824 22520 40830
rect 22589 40827 22659 40832
rect 21963 39864 22041 39869
rect 21963 39796 21968 39864
rect 22036 39796 22041 39864
rect 21963 39791 22041 39796
rect 22572 38445 22640 38450
rect 22572 38387 22577 38445
rect 22635 38387 22640 38445
rect 22572 35829 22640 38387
rect 23202 37600 23386 40696
rect 23994 39429 24178 40696
rect 23913 39423 24211 39429
rect 23913 39119 24211 39125
rect 23994 38342 24178 39119
rect 22567 35824 22645 35829
rect 22567 35756 22572 35824
rect 22640 35756 22645 35824
rect 22567 35751 22645 35756
rect 20505 30192 20583 30197
rect 20505 30124 20510 30192
rect 20578 30124 20583 30192
rect 20505 30119 20583 30124
rect 31313 700 31431 705
rect 14498 699 31432 700
rect 14498 695 31313 699
rect 14498 585 14503 695
rect 14613 585 31313 695
rect 14498 581 31313 585
rect 31431 581 31432 699
rect 14498 580 31432 581
rect 31313 575 31431 580
rect 12694 417 27016 418
rect 12694 413 26897 417
rect 12694 303 12699 413
rect 12809 303 26897 413
rect 12694 299 26897 303
rect 27015 299 27021 417
rect 12694 298 27016 299
<< via3 >>
rect 17724 44782 17788 44846
rect 14044 44714 14108 44778
rect 16988 44614 17052 44678
rect 22642 44668 22706 44732
rect 30972 44668 31036 44732
rect 14780 44546 14844 44610
rect 12572 44378 12636 44442
rect 13308 44378 13372 44442
rect 15516 44436 15580 44500
rect 22454 44462 22518 44526
rect 29500 44462 29564 44526
rect 16252 44066 16316 44130
rect 22642 41494 22706 41558
rect 4711 39125 5009 39423
rect 10579 39125 10877 39423
rect 12301 38083 12599 38381
rect 13851 39125 14149 39423
rect 19875 39125 20173 39423
rect 22456 40830 22520 40894
rect 23913 39125 24211 39423
rect 31313 581 31431 699
rect 26897 299 27015 417
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44443 12634 45152
rect 13310 44443 13370 45152
rect 14046 44779 14106 45152
rect 14043 44778 14109 44779
rect 14043 44714 14044 44778
rect 14108 44714 14109 44778
rect 14043 44713 14109 44714
rect 14782 44611 14842 45152
rect 14779 44610 14845 44611
rect 14779 44546 14780 44610
rect 14844 44546 14845 44610
rect 14779 44545 14845 44546
rect 15518 44501 15578 45152
rect 15515 44500 15581 44501
rect 12571 44442 12637 44443
rect 12571 44378 12572 44442
rect 12636 44378 12637 44442
rect 12571 44377 12637 44378
rect 13307 44442 13373 44443
rect 13307 44378 13308 44442
rect 13372 44378 13373 44442
rect 15515 44436 15516 44500
rect 15580 44436 15581 44500
rect 15515 44435 15581 44436
rect 15518 44409 15578 44435
rect 13307 44377 13373 44378
rect 200 39424 500 44152
rect 16254 44131 16314 45152
rect 16990 44679 17050 45152
rect 17726 44847 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 17723 44846 17789 44847
rect 17723 44782 17724 44846
rect 17788 44782 17789 44846
rect 17723 44781 17789 44782
rect 22641 44732 22707 44733
rect 16987 44678 17053 44679
rect 16987 44614 16988 44678
rect 17052 44614 17053 44678
rect 22641 44668 22642 44732
rect 22706 44668 22707 44732
rect 22641 44667 22707 44668
rect 16987 44613 17053 44614
rect 22458 44527 22518 44538
rect 22453 44526 22519 44527
rect 22453 44462 22454 44526
rect 22518 44462 22519 44526
rect 22453 44461 22519 44462
rect 16251 44130 16317 44131
rect 16251 44066 16252 44130
rect 16316 44066 16317 44130
rect 16251 44065 16317 44066
rect 22458 40895 22518 44461
rect 22644 41559 22704 44667
rect 29502 44527 29562 45152
rect 30238 44952 30298 45152
rect 30974 44733 31034 45152
rect 31710 44952 31770 45152
rect 30971 44732 31037 44733
rect 30971 44668 30972 44732
rect 31036 44668 31037 44732
rect 30971 44667 31037 44668
rect 29499 44526 29565 44527
rect 29499 44462 29500 44526
rect 29564 44462 29565 44526
rect 29499 44461 29565 44462
rect 22641 41558 22707 41559
rect 22641 41494 22642 41558
rect 22706 41494 22707 41558
rect 22641 41493 22707 41494
rect 22455 40894 22521 40895
rect 22455 40830 22456 40894
rect 22520 40830 22521 40894
rect 22455 40829 22521 40830
rect 200 39423 24224 39424
rect 200 39125 4711 39423
rect 5009 39125 10579 39423
rect 10877 39125 13851 39423
rect 14149 39125 19875 39423
rect 20173 39125 23913 39423
rect 24211 39125 24224 39423
rect 200 39124 24224 39125
rect 200 1000 500 39124
rect 31200 38382 31500 44152
rect 1958 38381 31500 38382
rect 1958 38083 12301 38381
rect 12599 38083 31500 38381
rect 1958 38082 31500 38083
rect 31200 1000 31500 38082
rect 31312 699 31432 700
rect 31312 581 31313 699
rect 31431 581 31432 699
rect 26896 417 27016 418
rect 26896 299 26897 417
rect 27015 299 27016 417
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 299
rect 31312 0 31432 581
use SUNSAR_SAR8B_CV  SUNSAR_SAR8B_CV_0 SUN_SAR9B_SKY130NM
timestamp 1708687947
transform 1 0 2448 0 1 2648
box -1922 -1864 24278 37062
use SUNSAR_SARCAPTURE_CV  SUNSAR_SARCAPTURE_CV_0 SUN_SAR9B_SKY130NM
timestamp 1708687947
transform 1 0 2286 0 1 40066
box -180 -132 22860 4356
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 200 1000 500 44152 0 FreeSans 2000 90 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 s 31200 1000 31500 44152 0 FreeSans 2000 90 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
