VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_TT06_SAR_wulffern
  CLASS BLOCK ;
  FOREIGN tt_um_TT06_SAR_wulffern ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 156.000 5.000 157.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 13.060 138.570 20.260 212.050 ;
      LAYER nwell ;
        RECT 20.260 138.570 32.860 212.050 ;
      LAYER pwell ;
        RECT 32.860 138.570 45.460 212.050 ;
      LAYER nwell ;
        RECT 45.460 138.570 58.060 212.050 ;
      LAYER pwell ;
        RECT 58.060 138.570 70.660 212.050 ;
      LAYER nwell ;
        RECT 70.660 138.570 83.260 212.050 ;
      LAYER pwell ;
        RECT 83.260 138.570 95.860 212.050 ;
      LAYER nwell ;
        RECT 95.860 138.570 108.460 212.050 ;
      LAYER pwell ;
        RECT 108.460 210.290 115.660 212.050 ;
        RECT 108.460 138.570 121.060 210.290 ;
      LAYER nwell ;
        RECT 121.060 138.570 128.260 210.290 ;
        RECT 49.960 12.580 57.160 33.260 ;
      LAYER pwell ;
        RECT 57.160 27.980 64.360 33.260 ;
        RECT 76.960 27.980 84.160 33.260 ;
        RECT 57.160 12.580 84.160 27.980 ;
      LAYER nwell ;
        RECT 84.160 12.580 91.360 33.260 ;
      LAYER pwell ;
        RECT 139.000 2.000 146.200 223.320 ;
      LAYER nwell ;
        RECT 146.200 2.000 153.400 223.320 ;
      LAYER li1 ;
        RECT 4.020 207.450 4.320 222.190 ;
        RECT 5.040 221.190 135.520 222.190 ;
        RECT 5.040 217.590 135.520 218.590 ;
        RECT 4.000 206.530 4.340 207.450 ;
        RECT 4.020 4.300 4.320 206.530 ;
        RECT 5.040 7.040 6.040 217.590 ;
        RECT 8.640 213.990 131.920 214.990 ;
        RECT 8.640 10.640 9.640 213.990 ;
        RECT 13.420 210.660 14.500 211.610 ;
        RECT 17.740 211.100 18.660 211.140 ;
        RECT 21.700 211.100 22.620 211.140 ;
        RECT 16.960 210.800 18.820 211.100 ;
        RECT 21.700 210.800 23.380 211.100 ;
        RECT 16.960 210.660 17.260 210.800 ;
        RECT 13.420 210.360 17.260 210.660 ;
        RECT 13.420 140.260 14.500 210.360 ;
        RECT 16.960 210.220 17.260 210.360 ;
        RECT 23.080 210.660 23.380 210.800 ;
        RECT 26.020 210.660 27.100 211.610 ;
        RECT 30.500 211.100 31.420 211.140 ;
        RECT 34.460 211.100 35.380 211.140 ;
        RECT 29.740 210.800 31.420 211.100 ;
        RECT 34.300 210.800 36.160 211.100 ;
        RECT 29.740 210.660 30.040 210.800 ;
        RECT 23.080 210.360 30.040 210.660 ;
        RECT 17.740 210.220 18.660 210.260 ;
        RECT 21.700 210.220 22.620 210.260 ;
        RECT 23.080 210.220 23.380 210.360 ;
        RECT 16.960 209.920 18.820 210.220 ;
        RECT 21.700 209.920 23.380 210.220 ;
        RECT 21.700 209.340 22.620 209.570 ;
        RECT 17.740 209.040 22.780 209.340 ;
        RECT 15.580 208.600 17.260 208.900 ;
        RECT 23.860 208.600 24.940 208.900 ;
        RECT 15.580 207.140 16.500 207.180 ;
        RECT 15.580 206.840 16.660 207.140 ;
        RECT 16.960 206.700 17.260 208.600 ;
        RECT 17.740 208.460 18.660 208.500 ;
        RECT 21.700 208.460 22.620 208.500 ;
        RECT 17.740 208.160 18.820 208.460 ;
        RECT 21.700 208.160 22.780 208.460 ;
        RECT 17.740 207.580 18.660 207.620 ;
        RECT 17.740 207.280 18.820 207.580 ;
        RECT 19.120 207.280 22.780 207.580 ;
        RECT 19.120 206.700 19.420 207.280 ;
        RECT 23.860 206.840 24.940 207.140 ;
        RECT 16.960 206.400 19.420 206.700 ;
        RECT 21.700 206.400 22.780 206.700 ;
        RECT 19.120 205.820 19.420 206.400 ;
        RECT 22.090 205.820 22.390 206.400 ;
        RECT 17.740 205.520 19.420 205.820 ;
        RECT 21.700 205.520 22.780 205.820 ;
        RECT 15.580 205.080 16.660 205.380 ;
        RECT 23.860 205.080 24.940 205.380 ;
        RECT 16.360 204.780 17.260 205.080 ;
        RECT 16.960 204.060 17.260 204.780 ;
        RECT 17.740 204.940 18.660 204.980 ;
        RECT 21.700 204.940 22.620 204.980 ;
        RECT 17.740 204.640 18.820 204.940 ;
        RECT 21.700 204.640 22.780 204.940 ;
        RECT 16.960 203.760 22.780 204.060 ;
        RECT 15.580 203.320 16.660 203.620 ;
        RECT 23.860 203.320 24.940 203.620 ;
        RECT 16.360 203.020 17.260 203.320 ;
        RECT 16.960 202.300 17.260 203.020 ;
        RECT 17.740 203.180 18.660 203.220 ;
        RECT 21.700 203.180 22.620 203.220 ;
        RECT 17.740 202.880 18.820 203.180 ;
        RECT 21.700 202.880 22.780 203.180 ;
        RECT 21.700 202.300 22.620 202.340 ;
        RECT 16.960 202.000 19.420 202.300 ;
        RECT 21.700 202.000 22.780 202.300 ;
        RECT 15.580 201.860 16.500 201.900 ;
        RECT 15.580 201.560 16.660 201.860 ;
        RECT 19.120 201.420 19.420 202.000 ;
        RECT 23.860 201.560 24.940 201.860 ;
        RECT 17.740 201.120 18.820 201.420 ;
        RECT 19.120 201.120 22.780 201.420 ;
        RECT 18.130 200.540 18.430 201.120 ;
        RECT 19.120 200.540 19.420 201.120 ;
        RECT 17.740 200.240 18.820 200.540 ;
        RECT 19.120 200.240 22.780 200.540 ;
        RECT 15.580 199.800 16.660 200.100 ;
        RECT 23.860 199.800 24.940 200.100 ;
        RECT 15.970 198.340 16.270 199.800 ;
        RECT 17.740 199.660 18.660 199.700 ;
        RECT 21.700 199.660 22.620 199.700 ;
        RECT 17.740 199.360 18.820 199.660 ;
        RECT 21.700 199.360 22.780 199.660 ;
        RECT 17.740 198.480 22.780 198.780 ;
        RECT 15.580 198.040 17.260 198.340 ;
        RECT 23.860 198.040 24.940 198.340 ;
        RECT 16.960 197.020 17.260 198.040 ;
        RECT 17.740 197.900 18.660 197.940 ;
        RECT 21.700 197.900 22.620 197.940 ;
        RECT 17.740 197.600 18.820 197.900 ;
        RECT 21.700 197.600 22.780 197.900 ;
        RECT 16.960 196.720 22.780 197.020 ;
        RECT 23.860 196.580 24.780 196.620 ;
        RECT 15.580 196.280 16.660 196.580 ;
        RECT 23.860 196.280 24.940 196.580 ;
        RECT 17.740 196.140 18.660 196.180 ;
        RECT 21.700 196.140 22.620 196.180 ;
        RECT 17.740 195.840 18.820 196.140 ;
        RECT 21.700 195.840 22.780 196.140 ;
        RECT 17.740 195.260 18.660 195.300 ;
        RECT 17.740 194.960 22.780 195.260 ;
        RECT 15.580 194.520 16.660 194.820 ;
        RECT 15.970 193.060 16.270 194.520 ;
        RECT 17.740 194.080 18.820 194.380 ;
        RECT 18.130 193.500 18.430 194.080 ;
        RECT 17.740 193.200 18.820 193.500 ;
        RECT 15.580 192.760 16.660 193.060 ;
        RECT 15.970 191.340 16.270 192.760 ;
        RECT 17.740 192.620 18.660 192.660 ;
        RECT 17.740 192.320 18.820 192.620 ;
        RECT 18.130 191.780 18.430 192.320 ;
        RECT 17.740 191.740 18.660 191.780 ;
        RECT 17.740 191.440 18.820 191.740 ;
        RECT 15.580 191.300 16.500 191.340 ;
        RECT 15.580 191.000 16.660 191.300 ;
        RECT 15.970 189.540 16.270 191.000 ;
        RECT 17.740 190.560 18.820 190.860 ;
        RECT 18.130 189.980 18.430 190.560 ;
        RECT 17.740 189.680 18.820 189.980 ;
        RECT 15.580 189.240 16.660 189.540 ;
        RECT 17.740 189.100 18.660 189.140 ;
        RECT 19.120 189.100 19.420 194.960 ;
        RECT 23.860 194.520 24.940 194.820 ;
        RECT 21.700 194.080 22.780 194.380 ;
        RECT 22.090 193.500 22.390 194.080 ;
        RECT 21.700 193.200 22.780 193.500 ;
        RECT 24.250 193.100 24.550 194.520 ;
        RECT 23.860 193.060 24.780 193.100 ;
        RECT 23.860 192.760 24.940 193.060 ;
        RECT 21.700 192.620 22.620 192.660 ;
        RECT 21.700 192.320 22.780 192.620 ;
        RECT 22.090 191.780 22.390 192.320 ;
        RECT 21.700 191.740 22.620 191.780 ;
        RECT 21.700 191.440 22.780 191.740 ;
        RECT 23.860 191.000 24.940 191.300 ;
        RECT 21.700 190.560 22.780 190.860 ;
        RECT 22.090 189.980 22.390 190.560 ;
        RECT 21.700 189.680 22.780 189.980 ;
        RECT 24.250 189.540 24.550 191.000 ;
        RECT 23.080 189.240 24.940 189.540 ;
        RECT 17.740 188.800 18.820 189.100 ;
        RECT 19.120 188.800 22.780 189.100 ;
        RECT 17.740 188.220 18.660 188.260 ;
        RECT 21.700 188.220 22.620 188.260 ;
        RECT 17.740 187.920 18.820 188.220 ;
        RECT 21.700 187.920 22.780 188.220 ;
        RECT 15.580 187.480 16.660 187.780 ;
        RECT 15.970 186.020 16.270 187.480 ;
        RECT 17.740 187.040 18.820 187.340 ;
        RECT 21.700 187.040 22.780 187.340 ;
        RECT 18.130 186.460 18.430 187.040 ;
        RECT 22.090 186.460 22.390 187.040 ;
        RECT 17.740 186.160 22.780 186.460 ;
        RECT 15.580 185.720 16.660 186.020 ;
        RECT 15.970 184.260 16.270 185.720 ;
        RECT 17.740 185.580 18.660 185.620 ;
        RECT 17.740 185.280 18.820 185.580 ;
        RECT 18.130 184.740 18.430 185.280 ;
        RECT 17.740 184.700 18.660 184.740 ;
        RECT 17.740 184.400 18.820 184.700 ;
        RECT 15.580 183.960 16.660 184.260 ;
        RECT 15.970 182.500 16.270 183.960 ;
        RECT 17.740 183.520 18.820 183.820 ;
        RECT 18.130 182.940 18.430 183.520 ;
        RECT 19.120 182.940 19.420 186.160 ;
        RECT 21.700 185.280 22.780 185.580 ;
        RECT 22.090 184.740 22.390 185.280 ;
        RECT 21.700 184.700 22.620 184.740 ;
        RECT 21.700 184.400 22.780 184.700 ;
        RECT 21.700 183.520 22.780 183.820 ;
        RECT 20.910 182.940 21.250 183.210 ;
        RECT 22.090 182.940 22.390 183.520 ;
        RECT 23.080 182.940 23.380 189.240 ;
        RECT 23.860 187.480 24.940 187.780 ;
        RECT 24.250 186.020 24.550 187.480 ;
        RECT 23.860 185.720 24.940 186.020 ;
        RECT 24.250 184.260 24.550 185.720 ;
        RECT 23.860 183.960 24.940 184.260 ;
        RECT 17.740 182.640 23.380 182.940 ;
        RECT 15.580 182.200 17.260 182.500 ;
        RECT 20.910 182.290 21.250 182.640 ;
        RECT 24.250 182.500 24.550 183.960 ;
        RECT 23.860 182.200 24.940 182.500 ;
        RECT 15.580 180.440 16.660 180.740 ;
        RECT 15.970 178.980 16.270 180.440 ;
        RECT 15.580 178.680 16.660 178.980 ;
        RECT 15.970 177.220 16.270 178.680 ;
        RECT 15.580 176.920 16.660 177.220 ;
        RECT 15.970 175.500 16.270 176.920 ;
        RECT 16.960 175.900 17.260 182.200 ;
        RECT 17.740 182.060 18.660 182.100 ;
        RECT 21.700 182.060 22.620 182.100 ;
        RECT 17.740 181.760 18.820 182.060 ;
        RECT 21.700 181.760 22.780 182.060 ;
        RECT 17.740 181.180 18.660 181.220 ;
        RECT 21.700 181.180 22.620 181.220 ;
        RECT 17.740 180.880 18.820 181.180 ;
        RECT 21.700 180.880 22.780 181.180 ;
        RECT 23.860 180.440 24.940 180.740 ;
        RECT 17.740 180.000 18.820 180.300 ;
        RECT 21.700 180.000 22.780 180.300 ;
        RECT 18.130 179.420 18.430 180.000 ;
        RECT 22.090 179.420 22.390 180.000 ;
        RECT 17.740 179.120 22.780 179.420 ;
        RECT 17.740 178.540 18.660 178.580 ;
        RECT 17.740 178.240 18.820 178.540 ;
        RECT 18.130 177.700 18.430 178.240 ;
        RECT 17.740 177.660 18.660 177.700 ;
        RECT 17.740 177.360 18.820 177.660 ;
        RECT 17.740 176.480 18.820 176.780 ;
        RECT 18.130 175.900 18.430 176.480 ;
        RECT 19.120 175.900 19.420 179.120 ;
        RECT 24.250 178.980 24.550 180.440 ;
        RECT 23.860 178.680 24.940 178.980 ;
        RECT 21.700 178.240 22.780 178.540 ;
        RECT 22.090 177.700 22.390 178.240 ;
        RECT 21.700 177.660 22.620 177.700 ;
        RECT 21.700 177.360 22.780 177.660 ;
        RECT 24.250 177.220 24.550 178.680 ;
        RECT 23.860 176.920 24.940 177.220 ;
        RECT 21.700 176.480 22.780 176.780 ;
        RECT 20.035 175.900 20.375 176.170 ;
        RECT 22.090 175.900 22.390 176.480 ;
        RECT 16.960 175.600 22.780 175.900 ;
        RECT 15.580 175.460 16.500 175.500 ;
        RECT 15.580 175.160 16.660 175.460 ;
        RECT 20.035 175.250 20.375 175.600 ;
        RECT 24.250 175.460 24.550 176.920 ;
        RECT 23.860 175.160 24.940 175.460 ;
        RECT 17.740 175.020 18.660 175.060 ;
        RECT 21.700 175.020 22.620 175.060 ;
        RECT 17.740 174.720 18.820 175.020 ;
        RECT 21.700 174.720 22.780 175.020 ;
        RECT 17.740 174.140 18.660 174.180 ;
        RECT 21.700 174.140 22.620 174.180 ;
        RECT 17.740 173.840 18.820 174.140 ;
        RECT 21.700 173.840 22.780 174.140 ;
        RECT 15.580 173.400 16.660 173.700 ;
        RECT 23.860 173.400 24.940 173.700 ;
        RECT 15.970 171.940 16.270 173.400 ;
        RECT 17.740 172.960 18.820 173.260 ;
        RECT 21.700 172.960 22.780 173.260 ;
        RECT 18.130 172.380 18.430 172.960 ;
        RECT 22.090 172.380 22.390 172.960 ;
        RECT 17.740 172.080 22.780 172.380 ;
        RECT 15.580 171.640 16.660 171.940 ;
        RECT 15.970 170.180 16.270 171.640 ;
        RECT 17.740 171.500 18.660 171.540 ;
        RECT 17.740 171.200 18.820 171.500 ;
        RECT 18.130 170.660 18.430 171.200 ;
        RECT 17.740 170.620 18.660 170.660 ;
        RECT 17.740 170.320 18.820 170.620 ;
        RECT 15.580 169.880 16.660 170.180 ;
        RECT 15.970 168.420 16.270 169.880 ;
        RECT 17.740 169.440 18.820 169.740 ;
        RECT 18.130 168.860 18.430 169.440 ;
        RECT 19.120 169.130 19.420 172.080 ;
        RECT 24.250 171.940 24.550 173.400 ;
        RECT 23.860 171.640 24.940 171.940 ;
        RECT 21.700 171.200 22.780 171.500 ;
        RECT 22.090 170.660 22.390 171.200 ;
        RECT 21.700 170.620 22.620 170.660 ;
        RECT 21.700 170.320 22.780 170.620 ;
        RECT 24.250 170.180 24.550 171.640 ;
        RECT 23.860 169.880 24.940 170.180 ;
        RECT 21.700 169.440 22.780 169.740 ;
        RECT 19.120 168.860 19.575 169.130 ;
        RECT 22.090 168.900 22.390 169.440 ;
        RECT 21.700 168.860 22.620 168.900 ;
        RECT 17.740 168.560 22.780 168.860 ;
        RECT 15.580 168.120 17.260 168.420 ;
        RECT 19.235 168.210 19.575 168.560 ;
        RECT 24.250 168.420 24.550 169.880 ;
        RECT 23.860 168.120 24.940 168.420 ;
        RECT 15.660 168.080 16.580 168.120 ;
        RECT 15.580 166.360 16.660 166.660 ;
        RECT 15.970 164.900 16.270 166.360 ;
        RECT 15.580 164.600 16.660 164.900 ;
        RECT 15.970 163.140 16.270 164.600 ;
        RECT 15.580 162.840 16.660 163.140 ;
        RECT 15.970 161.380 16.270 162.840 ;
        RECT 16.960 161.820 17.260 168.120 ;
        RECT 17.740 167.980 18.660 168.020 ;
        RECT 21.700 167.980 22.620 168.020 ;
        RECT 17.740 167.680 18.820 167.980 ;
        RECT 21.700 167.680 22.780 167.980 ;
        RECT 17.740 167.100 18.660 167.140 ;
        RECT 21.700 167.100 22.620 167.140 ;
        RECT 17.740 166.800 18.820 167.100 ;
        RECT 21.700 166.800 22.780 167.100 ;
        RECT 23.860 166.360 24.940 166.660 ;
        RECT 17.740 165.920 18.820 166.220 ;
        RECT 21.700 165.920 22.780 166.220 ;
        RECT 18.130 165.340 18.430 165.920 ;
        RECT 22.090 165.340 22.390 165.920 ;
        RECT 17.740 165.040 22.780 165.340 ;
        RECT 17.740 164.460 18.660 164.500 ;
        RECT 17.740 164.160 18.820 164.460 ;
        RECT 18.130 163.620 18.430 164.160 ;
        RECT 17.740 163.580 18.660 163.620 ;
        RECT 17.740 163.280 18.820 163.580 ;
        RECT 17.740 162.400 18.820 162.700 ;
        RECT 18.130 161.820 18.430 162.400 ;
        RECT 19.120 161.820 19.420 165.040 ;
        RECT 24.250 164.900 24.550 166.360 ;
        RECT 23.860 164.600 24.940 164.900 ;
        RECT 21.700 164.160 22.780 164.460 ;
        RECT 22.090 163.620 22.390 164.160 ;
        RECT 21.700 163.580 22.620 163.620 ;
        RECT 21.700 163.280 22.780 163.580 ;
        RECT 24.250 163.140 24.550 164.600 ;
        RECT 23.860 162.840 24.940 163.140 ;
        RECT 21.700 162.400 22.780 162.700 ;
        RECT 22.090 161.820 22.390 162.400 ;
        RECT 16.960 161.520 22.780 161.820 ;
        RECT 24.250 161.380 24.550 162.840 ;
        RECT 15.580 161.080 16.660 161.380 ;
        RECT 23.260 161.080 24.940 161.380 ;
        RECT 17.740 160.940 18.660 160.980 ;
        RECT 21.700 160.940 22.620 160.980 ;
        RECT 17.740 160.640 18.820 160.940 ;
        RECT 21.700 160.640 22.780 160.940 ;
        RECT 23.260 160.060 23.560 161.080 ;
        RECT 17.740 159.760 23.560 160.060 ;
        RECT 15.580 159.620 16.500 159.660 ;
        RECT 23.860 159.620 24.780 159.660 ;
        RECT 15.580 159.320 16.660 159.620 ;
        RECT 23.860 159.320 25.540 159.620 ;
        RECT 17.740 158.880 18.820 159.180 ;
        RECT 21.700 158.880 22.780 159.180 ;
        RECT 18.130 158.300 18.430 158.880 ;
        RECT 22.090 158.300 22.390 158.880 ;
        RECT 17.740 158.000 18.820 158.300 ;
        RECT 21.700 158.000 22.780 158.300 ;
        RECT 24.250 157.860 24.550 159.320 ;
        RECT 15.580 157.560 17.260 157.860 ;
        RECT 23.860 157.560 24.940 157.860 ;
        RECT 15.580 156.100 16.500 156.140 ;
        RECT 14.980 155.800 16.660 156.100 ;
        RECT 14.980 143.780 15.280 155.800 ;
        RECT 15.580 154.340 16.500 154.380 ;
        RECT 15.580 154.040 16.660 154.340 ;
        RECT 16.960 152.580 17.260 157.560 ;
        RECT 17.740 157.120 18.820 157.420 ;
        RECT 21.700 157.120 22.780 157.420 ;
        RECT 18.130 156.540 18.430 157.120 ;
        RECT 22.090 156.540 22.390 157.120 ;
        RECT 17.740 156.240 18.820 156.540 ;
        RECT 21.700 156.240 22.780 156.540 ;
        RECT 24.250 156.100 24.550 157.560 ;
        RECT 23.860 155.800 24.940 156.100 ;
        RECT 17.740 155.660 18.660 155.700 ;
        RECT 21.700 155.660 22.620 155.700 ;
        RECT 17.740 155.360 18.820 155.660 ;
        RECT 21.700 155.360 22.780 155.660 ;
        RECT 17.740 154.780 18.660 154.820 ;
        RECT 17.740 154.480 22.780 154.780 ;
        RECT 25.240 154.340 25.540 159.320 ;
        RECT 23.860 154.040 25.540 154.340 ;
        RECT 17.740 153.600 18.820 153.900 ;
        RECT 21.700 153.600 22.780 153.900 ;
        RECT 18.130 153.020 18.430 153.600 ;
        RECT 22.090 153.020 22.390 153.600 ;
        RECT 17.740 152.720 18.820 153.020 ;
        RECT 21.700 152.720 22.780 153.020 ;
        RECT 24.250 152.580 24.550 154.040 ;
        RECT 15.580 152.280 17.260 152.580 ;
        RECT 23.860 152.280 24.940 152.580 ;
        RECT 15.740 150.820 16.660 150.860 ;
        RECT 15.580 150.520 16.660 150.820 ;
        RECT 16.960 149.500 17.260 152.280 ;
        RECT 17.740 151.840 18.820 152.140 ;
        RECT 21.700 151.840 22.780 152.140 ;
        RECT 18.130 151.260 18.430 151.840 ;
        RECT 22.090 151.260 22.390 151.840 ;
        RECT 17.740 150.960 18.820 151.260 ;
        RECT 21.700 150.960 22.780 151.260 ;
        RECT 24.250 150.820 24.550 152.280 ;
        RECT 23.860 150.520 24.940 150.820 ;
        RECT 17.740 150.380 18.660 150.420 ;
        RECT 21.700 150.380 22.620 150.420 ;
        RECT 17.740 150.080 18.820 150.380 ;
        RECT 21.700 150.080 22.780 150.380 ;
        RECT 16.960 149.200 22.780 149.500 ;
        RECT 15.580 148.760 16.660 149.060 ;
        RECT 23.860 148.760 24.940 149.060 ;
        RECT 16.360 148.460 17.260 148.760 ;
        RECT 16.960 147.740 17.260 148.460 ;
        RECT 17.740 148.620 18.660 148.660 ;
        RECT 21.700 148.620 22.620 148.660 ;
        RECT 17.740 148.320 18.820 148.620 ;
        RECT 21.700 148.320 22.780 148.620 ;
        RECT 21.700 147.740 22.620 147.780 ;
        RECT 16.960 147.440 21.400 147.740 ;
        RECT 21.700 147.440 22.780 147.740 ;
        RECT 15.580 147.000 16.660 147.300 ;
        RECT 17.740 146.860 18.660 146.900 ;
        RECT 17.740 146.560 18.820 146.860 ;
        RECT 17.740 145.980 18.660 146.020 ;
        RECT 17.740 145.680 18.820 145.980 ;
        RECT 15.740 145.540 16.660 145.580 ;
        RECT 15.580 145.240 16.660 145.540 ;
        RECT 17.740 144.800 19.420 145.100 ;
        RECT 19.120 144.220 19.420 144.800 ;
        RECT 17.740 143.920 19.420 144.220 ;
        RECT 14.980 143.480 16.660 143.780 ;
        RECT 17.740 143.340 18.660 143.380 ;
        RECT 17.740 143.040 18.820 143.340 ;
        RECT 19.120 142.460 19.420 143.920 ;
        RECT 21.100 143.340 21.400 147.440 ;
        RECT 23.080 147.000 24.940 147.300 ;
        RECT 21.700 146.560 22.780 146.860 ;
        RECT 22.090 145.980 22.390 146.560 ;
        RECT 21.700 145.680 22.780 145.980 ;
        RECT 21.700 144.800 22.780 145.100 ;
        RECT 22.090 144.220 22.390 144.800 ;
        RECT 21.700 143.920 22.780 144.220 ;
        RECT 21.700 143.340 22.620 143.380 ;
        RECT 21.100 143.040 22.780 143.340 ;
        RECT 17.740 142.160 19.420 142.460 ;
        RECT 21.700 142.460 22.620 142.500 ;
        RECT 21.700 142.160 22.780 142.460 ;
        RECT 15.580 142.020 16.500 142.060 ;
        RECT 15.580 141.720 16.660 142.020 ;
        RECT 23.080 141.580 23.380 147.000 ;
        RECT 23.860 145.240 24.940 145.540 ;
        RECT 23.860 143.480 24.940 143.780 ;
        RECT 25.240 142.020 25.540 154.040 ;
        RECT 23.860 141.720 25.540 142.020 ;
        RECT 17.740 141.280 23.380 141.580 ;
        RECT 17.740 140.700 18.660 140.740 ;
        RECT 21.700 140.700 22.620 140.740 ;
        RECT 16.960 140.400 18.820 140.700 ;
        RECT 21.700 140.400 23.380 140.700 ;
        RECT 16.960 140.260 17.260 140.400 ;
        RECT 13.420 139.960 17.260 140.260 ;
        RECT 13.420 139.010 14.500 139.960 ;
        RECT 16.960 139.820 17.260 139.960 ;
        RECT 23.080 140.260 23.380 140.400 ;
        RECT 26.020 140.260 27.100 210.360 ;
        RECT 29.740 210.220 30.040 210.360 ;
        RECT 35.860 210.660 36.160 210.800 ;
        RECT 38.620 210.660 39.700 211.610 ;
        RECT 42.940 211.100 43.860 211.140 ;
        RECT 46.900 211.100 47.820 211.140 ;
        RECT 42.160 210.800 44.020 211.100 ;
        RECT 46.900 210.800 48.580 211.100 ;
        RECT 42.160 210.660 42.460 210.800 ;
        RECT 35.860 210.360 42.460 210.660 ;
        RECT 30.500 210.220 31.420 210.260 ;
        RECT 34.460 210.220 35.380 210.260 ;
        RECT 35.860 210.220 36.160 210.360 ;
        RECT 29.740 209.920 31.420 210.220 ;
        RECT 34.300 209.920 36.160 210.220 ;
        RECT 30.340 209.340 31.260 209.380 ;
        RECT 30.340 209.040 35.380 209.340 ;
        RECT 28.180 208.600 29.260 208.900 ;
        RECT 35.860 208.600 37.540 208.900 ;
        RECT 30.500 208.460 31.420 208.500 ;
        RECT 34.460 208.460 35.380 208.500 ;
        RECT 30.340 208.160 31.420 208.460 ;
        RECT 34.300 208.160 35.380 208.460 ;
        RECT 34.460 207.580 35.380 207.620 ;
        RECT 30.340 207.280 34.000 207.580 ;
        RECT 34.300 207.280 35.380 207.580 ;
        RECT 28.180 206.840 29.260 207.140 ;
        RECT 33.700 206.700 34.000 207.280 ;
        RECT 35.860 206.700 36.160 208.600 ;
        RECT 36.460 207.140 37.380 207.180 ;
        RECT 36.460 206.840 37.540 207.140 ;
        RECT 30.340 206.400 31.420 206.700 ;
        RECT 33.700 206.400 36.160 206.700 ;
        RECT 30.730 205.820 31.030 206.400 ;
        RECT 33.700 205.820 34.000 206.400 ;
        RECT 30.340 205.520 31.420 205.820 ;
        RECT 33.700 205.520 35.380 205.820 ;
        RECT 28.180 205.080 29.260 205.380 ;
        RECT 36.460 205.080 37.540 205.380 ;
        RECT 30.500 204.940 31.420 204.980 ;
        RECT 34.460 204.940 35.380 204.980 ;
        RECT 30.340 204.640 31.420 204.940 ;
        RECT 34.300 204.640 35.380 204.940 ;
        RECT 35.860 204.780 36.760 205.080 ;
        RECT 35.860 204.060 36.160 204.780 ;
        RECT 30.340 203.760 36.160 204.060 ;
        RECT 28.180 203.320 29.260 203.620 ;
        RECT 36.460 203.320 37.540 203.620 ;
        RECT 30.500 203.180 31.420 203.220 ;
        RECT 34.460 203.180 35.380 203.220 ;
        RECT 30.340 202.880 31.420 203.180 ;
        RECT 34.300 202.880 35.380 203.180 ;
        RECT 35.860 203.020 36.760 203.320 ;
        RECT 30.500 202.300 31.420 202.340 ;
        RECT 35.860 202.300 36.160 203.020 ;
        RECT 30.340 202.000 31.420 202.300 ;
        RECT 33.700 202.000 36.160 202.300 ;
        RECT 28.180 201.560 29.260 201.860 ;
        RECT 33.700 201.420 34.000 202.000 ;
        RECT 36.620 201.860 37.540 201.900 ;
        RECT 36.460 201.560 37.540 201.860 ;
        RECT 30.340 201.120 34.000 201.420 ;
        RECT 34.300 201.120 35.380 201.420 ;
        RECT 33.700 200.540 34.000 201.120 ;
        RECT 34.690 200.540 34.990 201.120 ;
        RECT 30.340 200.240 34.000 200.540 ;
        RECT 34.300 200.240 35.380 200.540 ;
        RECT 28.180 199.800 29.260 200.100 ;
        RECT 36.460 199.800 37.540 200.100 ;
        RECT 30.500 199.660 31.420 199.700 ;
        RECT 34.460 199.660 35.380 199.700 ;
        RECT 30.340 199.360 31.420 199.660 ;
        RECT 34.300 199.360 35.380 199.660 ;
        RECT 30.340 198.480 35.380 198.780 ;
        RECT 36.850 198.340 37.150 199.800 ;
        RECT 28.180 198.040 29.260 198.340 ;
        RECT 35.860 198.040 37.540 198.340 ;
        RECT 30.500 197.900 31.420 197.940 ;
        RECT 34.460 197.900 35.380 197.940 ;
        RECT 30.340 197.600 31.420 197.900 ;
        RECT 34.300 197.600 35.380 197.900 ;
        RECT 35.860 197.020 36.160 198.040 ;
        RECT 30.340 196.720 36.160 197.020 ;
        RECT 28.340 196.580 29.260 196.620 ;
        RECT 28.180 196.280 29.260 196.580 ;
        RECT 36.460 196.280 37.540 196.580 ;
        RECT 30.500 196.140 31.420 196.180 ;
        RECT 34.460 196.140 35.380 196.180 ;
        RECT 30.340 195.840 31.420 196.140 ;
        RECT 34.300 195.840 35.380 196.140 ;
        RECT 34.460 195.260 35.380 195.300 ;
        RECT 30.340 194.960 35.380 195.260 ;
        RECT 28.180 194.520 29.260 194.820 ;
        RECT 28.570 193.100 28.870 194.520 ;
        RECT 30.340 194.080 31.420 194.380 ;
        RECT 30.730 193.500 31.030 194.080 ;
        RECT 30.340 193.200 31.420 193.500 ;
        RECT 28.340 193.060 29.260 193.100 ;
        RECT 28.180 192.760 29.260 193.060 ;
        RECT 30.500 192.620 31.420 192.660 ;
        RECT 30.340 192.320 31.420 192.620 ;
        RECT 30.730 191.780 31.030 192.320 ;
        RECT 30.500 191.740 31.420 191.780 ;
        RECT 30.340 191.440 31.420 191.740 ;
        RECT 28.180 191.000 29.260 191.300 ;
        RECT 28.570 189.540 28.870 191.000 ;
        RECT 30.340 190.560 31.420 190.860 ;
        RECT 30.730 189.980 31.030 190.560 ;
        RECT 30.340 189.680 31.420 189.980 ;
        RECT 28.180 189.240 30.040 189.540 ;
        RECT 28.180 187.480 29.260 187.780 ;
        RECT 28.570 186.020 28.870 187.480 ;
        RECT 28.180 185.720 29.260 186.020 ;
        RECT 28.570 184.260 28.870 185.720 ;
        RECT 28.180 183.960 29.260 184.260 ;
        RECT 28.570 182.500 28.870 183.960 ;
        RECT 29.740 182.940 30.040 189.240 ;
        RECT 33.700 189.100 34.000 194.960 ;
        RECT 36.460 194.520 37.540 194.820 ;
        RECT 34.300 194.080 35.380 194.380 ;
        RECT 34.690 193.500 34.990 194.080 ;
        RECT 34.300 193.200 35.380 193.500 ;
        RECT 36.850 193.060 37.150 194.520 ;
        RECT 36.460 192.760 37.540 193.060 ;
        RECT 34.460 192.620 35.380 192.660 ;
        RECT 34.300 192.320 35.380 192.620 ;
        RECT 34.690 191.780 34.990 192.320 ;
        RECT 34.460 191.740 35.380 191.780 ;
        RECT 34.300 191.440 35.380 191.740 ;
        RECT 36.850 191.340 37.150 192.760 ;
        RECT 36.460 191.300 37.380 191.340 ;
        RECT 36.460 191.000 37.540 191.300 ;
        RECT 34.300 190.560 35.380 190.860 ;
        RECT 34.690 189.980 34.990 190.560 ;
        RECT 34.300 189.680 35.380 189.980 ;
        RECT 36.850 189.540 37.150 191.000 ;
        RECT 36.460 189.240 37.540 189.540 ;
        RECT 34.460 189.100 35.380 189.140 ;
        RECT 30.340 188.800 34.000 189.100 ;
        RECT 34.300 188.800 35.380 189.100 ;
        RECT 30.500 188.220 31.420 188.260 ;
        RECT 34.460 188.220 35.380 188.260 ;
        RECT 30.340 187.920 31.420 188.220 ;
        RECT 34.300 187.920 35.380 188.220 ;
        RECT 36.460 187.480 37.540 187.780 ;
        RECT 30.340 187.040 31.420 187.340 ;
        RECT 34.300 187.040 35.380 187.340 ;
        RECT 30.730 186.460 31.030 187.040 ;
        RECT 34.690 186.460 34.990 187.040 ;
        RECT 30.340 186.160 35.380 186.460 ;
        RECT 30.340 185.280 31.420 185.580 ;
        RECT 30.730 184.740 31.030 185.280 ;
        RECT 30.500 184.700 31.420 184.740 ;
        RECT 30.340 184.400 31.420 184.700 ;
        RECT 30.340 183.520 31.420 183.820 ;
        RECT 30.730 182.940 31.030 183.520 ;
        RECT 31.870 182.940 32.210 183.210 ;
        RECT 33.700 182.940 34.000 186.160 ;
        RECT 36.850 186.020 37.150 187.480 ;
        RECT 36.460 185.720 37.540 186.020 ;
        RECT 34.460 185.580 35.380 185.620 ;
        RECT 34.300 185.280 35.380 185.580 ;
        RECT 34.690 184.740 34.990 185.280 ;
        RECT 34.460 184.700 35.380 184.740 ;
        RECT 34.300 184.400 35.380 184.700 ;
        RECT 36.850 184.260 37.150 185.720 ;
        RECT 36.460 183.960 37.540 184.260 ;
        RECT 34.300 183.520 35.380 183.820 ;
        RECT 34.690 182.940 34.990 183.520 ;
        RECT 29.740 182.640 35.380 182.940 ;
        RECT 28.180 182.200 29.260 182.500 ;
        RECT 31.870 182.290 32.210 182.640 ;
        RECT 36.850 182.500 37.150 183.960 ;
        RECT 35.860 182.200 37.540 182.500 ;
        RECT 30.500 182.060 31.420 182.100 ;
        RECT 34.460 182.060 35.380 182.100 ;
        RECT 30.340 181.760 31.420 182.060 ;
        RECT 34.300 181.760 35.380 182.060 ;
        RECT 30.500 181.180 31.420 181.220 ;
        RECT 34.460 181.180 35.380 181.220 ;
        RECT 30.340 180.880 31.420 181.180 ;
        RECT 34.300 180.880 35.380 181.180 ;
        RECT 28.180 180.440 29.260 180.740 ;
        RECT 28.570 178.980 28.870 180.440 ;
        RECT 30.340 180.000 31.420 180.300 ;
        RECT 34.300 180.000 35.380 180.300 ;
        RECT 30.730 179.420 31.030 180.000 ;
        RECT 34.690 179.420 34.990 180.000 ;
        RECT 30.340 179.120 35.380 179.420 ;
        RECT 28.180 178.680 29.260 178.980 ;
        RECT 28.570 177.220 28.870 178.680 ;
        RECT 30.340 178.240 31.420 178.540 ;
        RECT 30.730 177.700 31.030 178.240 ;
        RECT 30.500 177.660 31.420 177.700 ;
        RECT 30.340 177.360 31.420 177.660 ;
        RECT 28.180 176.920 29.260 177.220 ;
        RECT 28.570 175.460 28.870 176.920 ;
        RECT 30.340 176.480 31.420 176.780 ;
        RECT 30.730 175.900 31.030 176.480 ;
        RECT 32.745 175.900 33.085 176.170 ;
        RECT 33.700 175.900 34.000 179.120 ;
        RECT 34.460 178.540 35.380 178.580 ;
        RECT 34.300 178.240 35.380 178.540 ;
        RECT 34.690 177.700 34.990 178.240 ;
        RECT 34.460 177.660 35.380 177.700 ;
        RECT 34.300 177.360 35.380 177.660 ;
        RECT 34.300 176.480 35.380 176.780 ;
        RECT 34.690 175.900 34.990 176.480 ;
        RECT 35.860 175.900 36.160 182.200 ;
        RECT 36.460 180.440 37.540 180.740 ;
        RECT 36.850 178.980 37.150 180.440 ;
        RECT 36.460 178.680 37.540 178.980 ;
        RECT 36.850 177.220 37.150 178.680 ;
        RECT 36.460 176.920 37.540 177.220 ;
        RECT 30.340 175.600 36.160 175.900 ;
        RECT 28.180 175.160 29.260 175.460 ;
        RECT 32.745 175.250 33.085 175.600 ;
        RECT 36.850 175.500 37.150 176.920 ;
        RECT 36.620 175.460 37.540 175.500 ;
        RECT 36.460 175.160 37.540 175.460 ;
        RECT 30.500 175.020 31.420 175.060 ;
        RECT 34.460 175.020 35.380 175.060 ;
        RECT 30.340 174.720 31.420 175.020 ;
        RECT 34.300 174.720 35.380 175.020 ;
        RECT 30.500 174.140 31.420 174.180 ;
        RECT 34.460 174.140 35.380 174.180 ;
        RECT 30.340 173.840 31.420 174.140 ;
        RECT 34.300 173.840 35.380 174.140 ;
        RECT 28.180 173.400 29.260 173.700 ;
        RECT 36.460 173.400 37.540 173.700 ;
        RECT 28.570 171.940 28.870 173.400 ;
        RECT 30.340 172.960 31.420 173.260 ;
        RECT 34.300 172.960 35.380 173.260 ;
        RECT 30.730 172.380 31.030 172.960 ;
        RECT 34.690 172.380 34.990 172.960 ;
        RECT 30.340 172.080 35.380 172.380 ;
        RECT 28.180 171.640 29.260 171.940 ;
        RECT 28.570 170.180 28.870 171.640 ;
        RECT 30.340 171.200 31.420 171.500 ;
        RECT 30.730 170.660 31.030 171.200 ;
        RECT 30.500 170.620 31.420 170.660 ;
        RECT 30.340 170.320 31.420 170.620 ;
        RECT 28.180 169.880 29.260 170.180 ;
        RECT 28.570 168.420 28.870 169.880 ;
        RECT 30.340 169.440 31.420 169.740 ;
        RECT 30.730 168.900 31.030 169.440 ;
        RECT 33.700 169.130 34.000 172.080 ;
        RECT 36.850 171.940 37.150 173.400 ;
        RECT 36.460 171.640 37.540 171.940 ;
        RECT 34.460 171.500 35.380 171.540 ;
        RECT 34.300 171.200 35.380 171.500 ;
        RECT 34.690 170.660 34.990 171.200 ;
        RECT 34.460 170.620 35.380 170.660 ;
        RECT 34.300 170.320 35.380 170.620 ;
        RECT 36.850 170.180 37.150 171.640 ;
        RECT 36.460 169.880 37.540 170.180 ;
        RECT 34.300 169.440 35.380 169.740 ;
        RECT 30.500 168.860 31.420 168.900 ;
        RECT 33.545 168.860 34.000 169.130 ;
        RECT 34.690 168.860 34.990 169.440 ;
        RECT 30.340 168.560 35.380 168.860 ;
        RECT 28.180 168.120 29.260 168.420 ;
        RECT 33.545 168.210 33.885 168.560 ;
        RECT 36.850 168.420 37.150 169.880 ;
        RECT 35.860 168.120 37.540 168.420 ;
        RECT 30.500 167.980 31.420 168.020 ;
        RECT 34.460 167.980 35.380 168.020 ;
        RECT 30.340 167.680 31.420 167.980 ;
        RECT 34.300 167.680 35.380 167.980 ;
        RECT 30.500 167.100 31.420 167.140 ;
        RECT 34.460 167.100 35.380 167.140 ;
        RECT 30.340 166.800 31.420 167.100 ;
        RECT 34.300 166.800 35.380 167.100 ;
        RECT 28.180 166.360 29.260 166.660 ;
        RECT 28.570 164.900 28.870 166.360 ;
        RECT 30.340 165.920 31.420 166.220 ;
        RECT 34.300 165.920 35.380 166.220 ;
        RECT 30.730 165.340 31.030 165.920 ;
        RECT 34.690 165.340 34.990 165.920 ;
        RECT 30.340 165.040 35.380 165.340 ;
        RECT 28.180 164.600 29.260 164.900 ;
        RECT 28.570 163.140 28.870 164.600 ;
        RECT 30.340 164.160 31.420 164.460 ;
        RECT 30.730 163.620 31.030 164.160 ;
        RECT 30.500 163.580 31.420 163.620 ;
        RECT 30.340 163.280 31.420 163.580 ;
        RECT 28.180 162.840 29.260 163.140 ;
        RECT 28.570 161.380 28.870 162.840 ;
        RECT 30.340 162.400 31.420 162.700 ;
        RECT 30.730 161.820 31.030 162.400 ;
        RECT 33.700 161.820 34.000 165.040 ;
        RECT 34.460 164.460 35.380 164.500 ;
        RECT 34.300 164.160 35.380 164.460 ;
        RECT 34.690 163.620 34.990 164.160 ;
        RECT 34.460 163.580 35.380 163.620 ;
        RECT 34.300 163.280 35.380 163.580 ;
        RECT 34.300 162.400 35.380 162.700 ;
        RECT 34.690 161.820 34.990 162.400 ;
        RECT 35.860 161.820 36.160 168.120 ;
        RECT 36.540 168.080 37.460 168.120 ;
        RECT 36.460 166.360 37.540 166.660 ;
        RECT 36.850 164.900 37.150 166.360 ;
        RECT 36.460 164.600 37.540 164.900 ;
        RECT 36.850 163.140 37.150 164.600 ;
        RECT 36.460 162.840 37.540 163.140 ;
        RECT 30.340 161.520 36.160 161.820 ;
        RECT 36.850 161.380 37.150 162.840 ;
        RECT 28.180 161.080 29.860 161.380 ;
        RECT 36.460 161.080 37.540 161.380 ;
        RECT 29.560 160.060 29.860 161.080 ;
        RECT 30.500 160.940 31.420 160.980 ;
        RECT 34.460 160.940 35.380 160.980 ;
        RECT 30.340 160.640 31.420 160.940 ;
        RECT 34.300 160.640 35.380 160.940 ;
        RECT 29.560 159.760 35.380 160.060 ;
        RECT 28.180 159.620 29.100 159.660 ;
        RECT 36.620 159.620 37.540 159.660 ;
        RECT 27.580 159.320 29.260 159.620 ;
        RECT 36.460 159.320 37.540 159.620 ;
        RECT 27.580 154.340 27.880 159.320 ;
        RECT 28.570 157.860 28.870 159.320 ;
        RECT 30.340 158.880 31.420 159.180 ;
        RECT 34.300 158.880 35.380 159.180 ;
        RECT 30.730 158.300 31.030 158.880 ;
        RECT 34.690 158.300 34.990 158.880 ;
        RECT 30.340 158.000 31.420 158.300 ;
        RECT 34.300 158.000 35.380 158.300 ;
        RECT 28.180 157.560 29.260 157.860 ;
        RECT 35.860 157.560 37.540 157.860 ;
        RECT 28.570 156.100 28.870 157.560 ;
        RECT 30.340 157.120 31.420 157.420 ;
        RECT 34.300 157.120 35.380 157.420 ;
        RECT 30.730 156.540 31.030 157.120 ;
        RECT 34.690 156.540 34.990 157.120 ;
        RECT 30.340 156.240 31.420 156.540 ;
        RECT 34.300 156.240 35.380 156.540 ;
        RECT 28.180 155.800 29.260 156.100 ;
        RECT 30.500 155.660 31.420 155.700 ;
        RECT 34.460 155.660 35.380 155.700 ;
        RECT 30.340 155.360 31.420 155.660 ;
        RECT 34.300 155.360 35.380 155.660 ;
        RECT 34.460 154.780 35.380 154.820 ;
        RECT 30.340 154.480 35.380 154.780 ;
        RECT 27.580 154.040 29.260 154.340 ;
        RECT 27.580 142.020 27.880 154.040 ;
        RECT 28.570 152.580 28.870 154.040 ;
        RECT 30.340 153.600 31.420 153.900 ;
        RECT 34.300 153.600 35.380 153.900 ;
        RECT 30.730 153.020 31.030 153.600 ;
        RECT 34.690 153.020 34.990 153.600 ;
        RECT 30.340 152.720 31.420 153.020 ;
        RECT 34.300 152.720 35.380 153.020 ;
        RECT 35.860 152.580 36.160 157.560 ;
        RECT 36.460 156.100 37.380 156.140 ;
        RECT 36.460 155.800 38.140 156.100 ;
        RECT 36.620 154.340 37.540 154.380 ;
        RECT 36.460 154.040 37.540 154.340 ;
        RECT 28.180 152.280 29.260 152.580 ;
        RECT 35.860 152.280 37.540 152.580 ;
        RECT 28.570 150.820 28.870 152.280 ;
        RECT 30.340 151.840 31.420 152.140 ;
        RECT 34.300 151.840 35.380 152.140 ;
        RECT 30.730 151.260 31.030 151.840 ;
        RECT 34.690 151.260 34.990 151.840 ;
        RECT 30.340 150.960 31.420 151.260 ;
        RECT 34.300 150.960 35.380 151.260 ;
        RECT 28.180 150.520 29.260 150.820 ;
        RECT 30.500 150.380 31.420 150.420 ;
        RECT 34.460 150.380 35.380 150.420 ;
        RECT 30.340 150.080 31.420 150.380 ;
        RECT 34.300 150.080 35.380 150.380 ;
        RECT 35.860 149.500 36.160 152.280 ;
        RECT 36.460 150.820 37.380 150.860 ;
        RECT 36.460 150.520 37.540 150.820 ;
        RECT 30.340 149.200 36.160 149.500 ;
        RECT 28.180 148.760 29.260 149.060 ;
        RECT 36.460 148.760 37.540 149.060 ;
        RECT 30.500 148.620 31.420 148.660 ;
        RECT 34.460 148.620 35.380 148.660 ;
        RECT 30.340 148.320 31.420 148.620 ;
        RECT 34.300 148.320 35.380 148.620 ;
        RECT 35.860 148.460 36.760 148.760 ;
        RECT 30.500 147.740 31.420 147.780 ;
        RECT 35.860 147.740 36.160 148.460 ;
        RECT 30.340 147.440 31.420 147.740 ;
        RECT 31.720 147.440 36.160 147.740 ;
        RECT 28.180 147.000 30.040 147.300 ;
        RECT 28.180 145.240 29.260 145.540 ;
        RECT 28.180 143.480 29.260 143.780 ;
        RECT 27.580 141.720 29.260 142.020 ;
        RECT 29.740 141.580 30.040 147.000 ;
        RECT 30.340 146.560 31.420 146.860 ;
        RECT 30.730 145.980 31.030 146.560 ;
        RECT 30.340 145.680 31.420 145.980 ;
        RECT 30.340 144.800 31.420 145.100 ;
        RECT 30.730 144.220 31.030 144.800 ;
        RECT 30.340 143.920 31.420 144.220 ;
        RECT 30.500 143.340 31.420 143.380 ;
        RECT 31.720 143.340 32.020 147.440 ;
        RECT 36.460 147.000 37.540 147.300 ;
        RECT 34.460 146.860 35.380 146.900 ;
        RECT 34.300 146.560 35.380 146.860 ;
        RECT 34.460 145.980 35.380 146.020 ;
        RECT 34.300 145.680 35.380 145.980 ;
        RECT 36.460 145.540 37.380 145.580 ;
        RECT 36.460 145.240 37.540 145.540 ;
        RECT 30.340 143.040 32.020 143.340 ;
        RECT 33.700 144.800 35.380 145.100 ;
        RECT 33.700 144.220 34.000 144.800 ;
        RECT 33.700 143.920 35.380 144.220 ;
        RECT 30.500 142.460 31.420 142.500 ;
        RECT 30.340 142.160 31.420 142.460 ;
        RECT 33.700 142.460 34.000 143.920 ;
        RECT 37.840 143.780 38.140 155.800 ;
        RECT 36.460 143.480 38.140 143.780 ;
        RECT 34.460 143.340 35.380 143.380 ;
        RECT 34.300 143.040 35.380 143.340 ;
        RECT 33.700 142.160 35.380 142.460 ;
        RECT 36.620 142.020 37.540 142.060 ;
        RECT 36.460 141.720 37.540 142.020 ;
        RECT 29.740 141.280 35.380 141.580 ;
        RECT 30.500 140.700 31.420 140.740 ;
        RECT 34.460 140.700 35.380 140.740 ;
        RECT 29.740 140.400 31.420 140.700 ;
        RECT 34.300 140.400 36.160 140.700 ;
        RECT 29.740 140.260 30.040 140.400 ;
        RECT 23.080 139.960 30.040 140.260 ;
        RECT 17.740 139.820 18.660 139.860 ;
        RECT 21.700 139.820 22.620 139.860 ;
        RECT 23.080 139.820 23.380 139.960 ;
        RECT 16.960 139.520 18.820 139.820 ;
        RECT 21.700 139.520 23.380 139.820 ;
        RECT 26.020 139.010 27.100 139.960 ;
        RECT 29.740 139.820 30.040 139.960 ;
        RECT 35.860 140.260 36.160 140.400 ;
        RECT 38.620 140.260 39.700 210.360 ;
        RECT 42.160 210.220 42.460 210.360 ;
        RECT 48.280 210.660 48.580 210.800 ;
        RECT 51.220 210.660 52.300 211.610 ;
        RECT 55.700 211.100 56.620 211.140 ;
        RECT 59.660 211.100 60.580 211.140 ;
        RECT 54.940 210.800 56.620 211.100 ;
        RECT 59.500 210.800 61.360 211.100 ;
        RECT 54.940 210.660 55.240 210.800 ;
        RECT 48.280 210.360 55.240 210.660 ;
        RECT 42.940 210.220 43.860 210.260 ;
        RECT 46.900 210.220 47.820 210.260 ;
        RECT 48.280 210.220 48.580 210.360 ;
        RECT 42.160 209.920 44.020 210.220 ;
        RECT 46.900 209.920 48.580 210.220 ;
        RECT 46.900 209.340 47.820 209.570 ;
        RECT 42.940 209.040 47.980 209.340 ;
        RECT 40.780 208.600 42.460 208.900 ;
        RECT 49.060 208.600 50.140 208.900 ;
        RECT 40.780 207.140 41.700 207.180 ;
        RECT 40.780 206.840 41.860 207.140 ;
        RECT 42.160 206.700 42.460 208.600 ;
        RECT 42.940 208.460 43.860 208.500 ;
        RECT 46.900 208.460 47.820 208.500 ;
        RECT 42.940 208.160 44.020 208.460 ;
        RECT 46.900 208.160 47.980 208.460 ;
        RECT 42.940 207.580 43.860 207.620 ;
        RECT 42.940 207.280 44.020 207.580 ;
        RECT 44.320 207.280 47.980 207.580 ;
        RECT 44.320 206.700 44.620 207.280 ;
        RECT 49.060 206.840 50.140 207.140 ;
        RECT 42.160 206.400 44.620 206.700 ;
        RECT 46.900 206.400 47.980 206.700 ;
        RECT 44.320 205.820 44.620 206.400 ;
        RECT 47.290 205.820 47.590 206.400 ;
        RECT 42.940 205.520 44.620 205.820 ;
        RECT 46.900 205.520 47.980 205.820 ;
        RECT 40.780 205.080 41.860 205.380 ;
        RECT 49.060 205.080 50.140 205.380 ;
        RECT 41.560 204.780 42.460 205.080 ;
        RECT 42.160 204.060 42.460 204.780 ;
        RECT 42.940 204.940 43.860 204.980 ;
        RECT 46.900 204.940 47.820 204.980 ;
        RECT 42.940 204.640 44.020 204.940 ;
        RECT 46.900 204.640 47.980 204.940 ;
        RECT 42.160 203.760 47.980 204.060 ;
        RECT 40.780 203.320 41.860 203.620 ;
        RECT 49.060 203.320 50.140 203.620 ;
        RECT 41.560 203.020 42.460 203.320 ;
        RECT 42.160 202.300 42.460 203.020 ;
        RECT 42.940 203.180 43.860 203.220 ;
        RECT 46.900 203.180 47.820 203.220 ;
        RECT 42.940 202.880 44.020 203.180 ;
        RECT 46.900 202.880 47.980 203.180 ;
        RECT 46.900 202.300 47.820 202.340 ;
        RECT 42.160 202.000 44.620 202.300 ;
        RECT 46.900 202.000 47.980 202.300 ;
        RECT 40.780 201.860 41.700 201.900 ;
        RECT 40.780 201.560 41.860 201.860 ;
        RECT 44.320 201.420 44.620 202.000 ;
        RECT 49.060 201.560 50.140 201.860 ;
        RECT 42.940 201.120 44.020 201.420 ;
        RECT 44.320 201.120 47.980 201.420 ;
        RECT 43.330 200.540 43.630 201.120 ;
        RECT 44.320 200.540 44.620 201.120 ;
        RECT 42.940 200.240 44.020 200.540 ;
        RECT 44.320 200.240 47.980 200.540 ;
        RECT 40.780 199.800 41.860 200.100 ;
        RECT 49.060 199.800 50.140 200.100 ;
        RECT 41.170 198.340 41.470 199.800 ;
        RECT 42.940 199.660 43.860 199.700 ;
        RECT 46.900 199.660 47.820 199.700 ;
        RECT 42.940 199.360 44.020 199.660 ;
        RECT 46.900 199.360 47.980 199.660 ;
        RECT 42.940 198.480 47.980 198.780 ;
        RECT 40.780 198.040 42.460 198.340 ;
        RECT 49.060 198.040 50.140 198.340 ;
        RECT 42.160 197.020 42.460 198.040 ;
        RECT 42.940 197.900 43.860 197.940 ;
        RECT 46.900 197.900 47.820 197.940 ;
        RECT 42.940 197.600 44.020 197.900 ;
        RECT 46.900 197.600 47.980 197.900 ;
        RECT 42.160 196.720 47.980 197.020 ;
        RECT 49.060 196.580 49.980 196.620 ;
        RECT 40.780 196.280 41.860 196.580 ;
        RECT 49.060 196.280 50.140 196.580 ;
        RECT 42.940 196.140 43.860 196.180 ;
        RECT 46.900 196.140 47.820 196.180 ;
        RECT 42.940 195.840 44.020 196.140 ;
        RECT 46.900 195.840 47.980 196.140 ;
        RECT 42.940 195.260 43.860 195.300 ;
        RECT 42.940 194.960 47.980 195.260 ;
        RECT 40.780 194.520 41.860 194.820 ;
        RECT 41.170 193.060 41.470 194.520 ;
        RECT 42.940 194.080 44.020 194.380 ;
        RECT 43.330 193.500 43.630 194.080 ;
        RECT 42.940 193.200 44.020 193.500 ;
        RECT 40.780 192.760 41.860 193.060 ;
        RECT 41.170 191.340 41.470 192.760 ;
        RECT 42.940 192.620 43.860 192.660 ;
        RECT 42.940 192.320 44.020 192.620 ;
        RECT 43.330 191.780 43.630 192.320 ;
        RECT 42.940 191.740 43.860 191.780 ;
        RECT 42.940 191.440 44.020 191.740 ;
        RECT 40.780 191.300 41.700 191.340 ;
        RECT 40.780 191.000 41.860 191.300 ;
        RECT 41.170 189.540 41.470 191.000 ;
        RECT 42.940 190.560 44.020 190.860 ;
        RECT 43.330 189.980 43.630 190.560 ;
        RECT 42.940 189.680 44.020 189.980 ;
        RECT 40.780 189.240 41.860 189.540 ;
        RECT 42.940 189.100 43.860 189.140 ;
        RECT 44.320 189.100 44.620 194.960 ;
        RECT 49.060 194.520 50.140 194.820 ;
        RECT 46.900 194.080 47.980 194.380 ;
        RECT 47.290 193.500 47.590 194.080 ;
        RECT 46.900 193.200 47.980 193.500 ;
        RECT 49.450 193.100 49.750 194.520 ;
        RECT 49.060 193.060 49.980 193.100 ;
        RECT 49.060 192.760 50.140 193.060 ;
        RECT 46.900 192.620 47.820 192.660 ;
        RECT 46.900 192.320 47.980 192.620 ;
        RECT 47.290 191.780 47.590 192.320 ;
        RECT 46.900 191.740 47.820 191.780 ;
        RECT 46.900 191.440 47.980 191.740 ;
        RECT 49.060 191.000 50.140 191.300 ;
        RECT 46.900 190.560 47.980 190.860 ;
        RECT 47.290 189.980 47.590 190.560 ;
        RECT 46.900 189.680 47.980 189.980 ;
        RECT 49.450 189.540 49.750 191.000 ;
        RECT 48.280 189.240 50.140 189.540 ;
        RECT 42.940 188.800 44.020 189.100 ;
        RECT 44.320 188.800 47.980 189.100 ;
        RECT 42.940 188.220 43.860 188.260 ;
        RECT 46.900 188.220 47.820 188.260 ;
        RECT 42.940 187.920 44.020 188.220 ;
        RECT 46.900 187.920 47.980 188.220 ;
        RECT 40.780 187.480 41.860 187.780 ;
        RECT 41.170 186.020 41.470 187.480 ;
        RECT 42.940 187.040 44.020 187.340 ;
        RECT 46.900 187.040 47.980 187.340 ;
        RECT 43.330 186.460 43.630 187.040 ;
        RECT 47.290 186.460 47.590 187.040 ;
        RECT 42.940 186.160 47.980 186.460 ;
        RECT 40.780 185.720 41.860 186.020 ;
        RECT 41.170 184.260 41.470 185.720 ;
        RECT 42.940 185.580 43.860 185.620 ;
        RECT 42.940 185.280 44.020 185.580 ;
        RECT 43.330 184.740 43.630 185.280 ;
        RECT 42.940 184.700 43.860 184.740 ;
        RECT 42.940 184.400 44.020 184.700 ;
        RECT 40.780 183.960 41.860 184.260 ;
        RECT 41.170 182.500 41.470 183.960 ;
        RECT 42.940 183.520 44.020 183.820 ;
        RECT 43.330 182.940 43.630 183.520 ;
        RECT 44.320 182.940 44.620 186.160 ;
        RECT 46.900 185.280 47.980 185.580 ;
        RECT 47.290 184.740 47.590 185.280 ;
        RECT 46.900 184.700 47.820 184.740 ;
        RECT 46.900 184.400 47.980 184.700 ;
        RECT 46.900 183.520 47.980 183.820 ;
        RECT 46.110 182.940 46.450 183.210 ;
        RECT 47.290 182.940 47.590 183.520 ;
        RECT 48.280 182.940 48.580 189.240 ;
        RECT 49.060 187.480 50.140 187.780 ;
        RECT 49.450 186.020 49.750 187.480 ;
        RECT 49.060 185.720 50.140 186.020 ;
        RECT 49.450 184.260 49.750 185.720 ;
        RECT 49.060 183.960 50.140 184.260 ;
        RECT 42.940 182.640 48.580 182.940 ;
        RECT 40.780 182.200 42.460 182.500 ;
        RECT 46.110 182.290 46.450 182.640 ;
        RECT 49.450 182.500 49.750 183.960 ;
        RECT 49.060 182.200 50.140 182.500 ;
        RECT 40.780 180.440 41.860 180.740 ;
        RECT 41.170 178.980 41.470 180.440 ;
        RECT 40.780 178.680 41.860 178.980 ;
        RECT 41.170 177.220 41.470 178.680 ;
        RECT 40.780 176.920 41.860 177.220 ;
        RECT 41.170 175.500 41.470 176.920 ;
        RECT 42.160 175.900 42.460 182.200 ;
        RECT 42.940 182.060 43.860 182.100 ;
        RECT 46.900 182.060 47.820 182.100 ;
        RECT 42.940 181.760 44.020 182.060 ;
        RECT 46.900 181.760 47.980 182.060 ;
        RECT 42.940 181.180 43.860 181.220 ;
        RECT 46.900 181.180 47.820 181.220 ;
        RECT 42.940 180.880 44.020 181.180 ;
        RECT 46.900 180.880 47.980 181.180 ;
        RECT 49.060 180.440 50.140 180.740 ;
        RECT 42.940 180.000 44.020 180.300 ;
        RECT 46.900 180.000 47.980 180.300 ;
        RECT 43.330 179.420 43.630 180.000 ;
        RECT 47.290 179.420 47.590 180.000 ;
        RECT 42.940 179.120 47.980 179.420 ;
        RECT 42.940 178.540 43.860 178.580 ;
        RECT 42.940 178.240 44.020 178.540 ;
        RECT 43.330 177.700 43.630 178.240 ;
        RECT 42.940 177.660 43.860 177.700 ;
        RECT 42.940 177.360 44.020 177.660 ;
        RECT 42.940 176.480 44.020 176.780 ;
        RECT 43.330 175.900 43.630 176.480 ;
        RECT 44.320 175.900 44.620 179.120 ;
        RECT 49.450 178.980 49.750 180.440 ;
        RECT 49.060 178.680 50.140 178.980 ;
        RECT 46.900 178.240 47.980 178.540 ;
        RECT 47.290 177.700 47.590 178.240 ;
        RECT 46.900 177.660 47.820 177.700 ;
        RECT 46.900 177.360 47.980 177.660 ;
        RECT 49.450 177.220 49.750 178.680 ;
        RECT 49.060 176.920 50.140 177.220 ;
        RECT 46.900 176.480 47.980 176.780 ;
        RECT 45.235 175.900 45.575 176.170 ;
        RECT 47.290 175.900 47.590 176.480 ;
        RECT 42.160 175.600 47.980 175.900 ;
        RECT 40.780 175.460 41.700 175.500 ;
        RECT 40.780 175.160 41.860 175.460 ;
        RECT 45.235 175.250 45.575 175.600 ;
        RECT 49.450 175.460 49.750 176.920 ;
        RECT 49.060 175.160 50.140 175.460 ;
        RECT 42.940 175.020 43.860 175.060 ;
        RECT 46.900 175.020 47.820 175.060 ;
        RECT 42.940 174.720 44.020 175.020 ;
        RECT 46.900 174.720 47.980 175.020 ;
        RECT 42.940 174.140 43.860 174.180 ;
        RECT 46.900 174.140 47.820 174.180 ;
        RECT 42.940 173.840 44.020 174.140 ;
        RECT 46.900 173.840 47.980 174.140 ;
        RECT 40.780 173.400 41.860 173.700 ;
        RECT 49.060 173.400 50.140 173.700 ;
        RECT 41.170 171.940 41.470 173.400 ;
        RECT 42.940 172.960 44.020 173.260 ;
        RECT 46.900 172.960 47.980 173.260 ;
        RECT 43.330 172.380 43.630 172.960 ;
        RECT 47.290 172.380 47.590 172.960 ;
        RECT 42.940 172.080 47.980 172.380 ;
        RECT 40.780 171.640 41.860 171.940 ;
        RECT 41.170 170.180 41.470 171.640 ;
        RECT 42.940 171.500 43.860 171.540 ;
        RECT 42.940 171.200 44.020 171.500 ;
        RECT 43.330 170.660 43.630 171.200 ;
        RECT 42.940 170.620 43.860 170.660 ;
        RECT 42.940 170.320 44.020 170.620 ;
        RECT 40.780 169.880 41.860 170.180 ;
        RECT 41.170 168.420 41.470 169.880 ;
        RECT 42.940 169.440 44.020 169.740 ;
        RECT 43.330 168.860 43.630 169.440 ;
        RECT 44.320 169.130 44.620 172.080 ;
        RECT 49.450 171.940 49.750 173.400 ;
        RECT 49.060 171.640 50.140 171.940 ;
        RECT 46.900 171.200 47.980 171.500 ;
        RECT 47.290 170.660 47.590 171.200 ;
        RECT 46.900 170.620 47.820 170.660 ;
        RECT 46.900 170.320 47.980 170.620 ;
        RECT 49.450 170.180 49.750 171.640 ;
        RECT 49.060 169.880 50.140 170.180 ;
        RECT 46.900 169.440 47.980 169.740 ;
        RECT 44.320 168.860 44.775 169.130 ;
        RECT 47.290 168.900 47.590 169.440 ;
        RECT 46.900 168.860 47.820 168.900 ;
        RECT 42.940 168.560 47.980 168.860 ;
        RECT 40.780 168.120 42.460 168.420 ;
        RECT 44.435 168.210 44.775 168.560 ;
        RECT 49.450 168.420 49.750 169.880 ;
        RECT 49.060 168.120 50.140 168.420 ;
        RECT 40.860 168.080 41.780 168.120 ;
        RECT 40.780 166.360 41.860 166.660 ;
        RECT 41.170 164.900 41.470 166.360 ;
        RECT 40.780 164.600 41.860 164.900 ;
        RECT 41.170 163.140 41.470 164.600 ;
        RECT 40.780 162.840 41.860 163.140 ;
        RECT 41.170 161.380 41.470 162.840 ;
        RECT 42.160 161.820 42.460 168.120 ;
        RECT 42.940 167.980 43.860 168.020 ;
        RECT 46.900 167.980 47.820 168.020 ;
        RECT 42.940 167.680 44.020 167.980 ;
        RECT 46.900 167.680 47.980 167.980 ;
        RECT 42.940 167.100 43.860 167.140 ;
        RECT 46.900 167.100 47.820 167.140 ;
        RECT 42.940 166.800 44.020 167.100 ;
        RECT 46.900 166.800 47.980 167.100 ;
        RECT 49.060 166.360 50.140 166.660 ;
        RECT 42.940 165.920 44.020 166.220 ;
        RECT 46.900 165.920 47.980 166.220 ;
        RECT 43.330 165.340 43.630 165.920 ;
        RECT 47.290 165.340 47.590 165.920 ;
        RECT 42.940 165.040 47.980 165.340 ;
        RECT 42.940 164.460 43.860 164.500 ;
        RECT 42.940 164.160 44.020 164.460 ;
        RECT 43.330 163.620 43.630 164.160 ;
        RECT 42.940 163.580 43.860 163.620 ;
        RECT 42.940 163.280 44.020 163.580 ;
        RECT 42.940 162.400 44.020 162.700 ;
        RECT 43.330 161.820 43.630 162.400 ;
        RECT 44.320 161.820 44.620 165.040 ;
        RECT 49.450 164.900 49.750 166.360 ;
        RECT 49.060 164.600 50.140 164.900 ;
        RECT 46.900 164.160 47.980 164.460 ;
        RECT 47.290 163.620 47.590 164.160 ;
        RECT 46.900 163.580 47.820 163.620 ;
        RECT 46.900 163.280 47.980 163.580 ;
        RECT 49.450 163.140 49.750 164.600 ;
        RECT 49.060 162.840 50.140 163.140 ;
        RECT 46.900 162.400 47.980 162.700 ;
        RECT 47.290 161.820 47.590 162.400 ;
        RECT 42.160 161.520 47.980 161.820 ;
        RECT 49.450 161.380 49.750 162.840 ;
        RECT 40.780 161.080 41.860 161.380 ;
        RECT 48.460 161.080 50.140 161.380 ;
        RECT 42.940 160.940 43.860 160.980 ;
        RECT 46.900 160.940 47.820 160.980 ;
        RECT 42.940 160.640 44.020 160.940 ;
        RECT 46.900 160.640 47.980 160.940 ;
        RECT 48.460 160.060 48.760 161.080 ;
        RECT 42.940 159.760 48.760 160.060 ;
        RECT 40.780 159.620 41.700 159.660 ;
        RECT 49.060 159.620 49.980 159.660 ;
        RECT 40.780 159.320 41.860 159.620 ;
        RECT 49.060 159.320 50.740 159.620 ;
        RECT 42.940 158.880 44.020 159.180 ;
        RECT 46.900 158.880 47.980 159.180 ;
        RECT 43.330 158.300 43.630 158.880 ;
        RECT 47.290 158.300 47.590 158.880 ;
        RECT 42.940 158.000 44.020 158.300 ;
        RECT 46.900 158.000 47.980 158.300 ;
        RECT 49.450 157.860 49.750 159.320 ;
        RECT 40.780 157.560 42.460 157.860 ;
        RECT 49.060 157.560 50.140 157.860 ;
        RECT 40.780 156.100 41.700 156.140 ;
        RECT 40.180 155.800 41.860 156.100 ;
        RECT 40.180 143.780 40.480 155.800 ;
        RECT 40.780 154.340 41.700 154.380 ;
        RECT 40.780 154.040 41.860 154.340 ;
        RECT 42.160 152.580 42.460 157.560 ;
        RECT 42.940 157.120 44.020 157.420 ;
        RECT 46.900 157.120 47.980 157.420 ;
        RECT 43.330 156.540 43.630 157.120 ;
        RECT 47.290 156.540 47.590 157.120 ;
        RECT 42.940 156.240 44.020 156.540 ;
        RECT 46.900 156.240 47.980 156.540 ;
        RECT 49.450 156.100 49.750 157.560 ;
        RECT 49.060 155.800 50.140 156.100 ;
        RECT 42.940 155.660 43.860 155.700 ;
        RECT 46.900 155.660 47.820 155.700 ;
        RECT 42.940 155.360 44.020 155.660 ;
        RECT 46.900 155.360 47.980 155.660 ;
        RECT 42.940 154.780 43.860 154.820 ;
        RECT 42.940 154.480 47.980 154.780 ;
        RECT 50.440 154.340 50.740 159.320 ;
        RECT 49.060 154.040 50.740 154.340 ;
        RECT 42.940 153.600 44.020 153.900 ;
        RECT 46.900 153.600 47.980 153.900 ;
        RECT 43.330 153.020 43.630 153.600 ;
        RECT 47.290 153.020 47.590 153.600 ;
        RECT 42.940 152.720 44.020 153.020 ;
        RECT 46.900 152.720 47.980 153.020 ;
        RECT 49.450 152.580 49.750 154.040 ;
        RECT 40.780 152.280 42.460 152.580 ;
        RECT 49.060 152.280 50.140 152.580 ;
        RECT 40.940 150.820 41.860 150.860 ;
        RECT 40.780 150.520 41.860 150.820 ;
        RECT 42.160 149.500 42.460 152.280 ;
        RECT 42.940 151.840 44.020 152.140 ;
        RECT 46.900 151.840 47.980 152.140 ;
        RECT 43.330 151.260 43.630 151.840 ;
        RECT 47.290 151.260 47.590 151.840 ;
        RECT 42.940 150.960 44.020 151.260 ;
        RECT 46.900 150.960 47.980 151.260 ;
        RECT 49.450 150.820 49.750 152.280 ;
        RECT 49.060 150.520 50.140 150.820 ;
        RECT 42.940 150.380 43.860 150.420 ;
        RECT 46.900 150.380 47.820 150.420 ;
        RECT 42.940 150.080 44.020 150.380 ;
        RECT 46.900 150.080 47.980 150.380 ;
        RECT 42.160 149.200 47.980 149.500 ;
        RECT 40.780 148.760 41.860 149.060 ;
        RECT 49.060 148.760 50.140 149.060 ;
        RECT 41.560 148.460 42.460 148.760 ;
        RECT 42.160 147.740 42.460 148.460 ;
        RECT 42.940 148.620 43.860 148.660 ;
        RECT 46.900 148.620 47.820 148.660 ;
        RECT 42.940 148.320 44.020 148.620 ;
        RECT 46.900 148.320 47.980 148.620 ;
        RECT 46.900 147.740 47.820 147.780 ;
        RECT 42.160 147.440 46.600 147.740 ;
        RECT 46.900 147.440 47.980 147.740 ;
        RECT 40.780 147.000 41.860 147.300 ;
        RECT 42.940 146.860 43.860 146.900 ;
        RECT 42.940 146.560 44.020 146.860 ;
        RECT 42.940 145.980 43.860 146.020 ;
        RECT 42.940 145.680 44.020 145.980 ;
        RECT 40.940 145.540 41.860 145.580 ;
        RECT 40.780 145.240 41.860 145.540 ;
        RECT 42.940 144.800 44.620 145.100 ;
        RECT 44.320 144.220 44.620 144.800 ;
        RECT 42.940 143.920 44.620 144.220 ;
        RECT 40.180 143.480 41.860 143.780 ;
        RECT 42.940 143.340 43.860 143.380 ;
        RECT 42.940 143.040 44.020 143.340 ;
        RECT 44.320 142.460 44.620 143.920 ;
        RECT 46.300 143.340 46.600 147.440 ;
        RECT 48.280 147.000 50.140 147.300 ;
        RECT 46.900 146.560 47.980 146.860 ;
        RECT 47.290 145.980 47.590 146.560 ;
        RECT 46.900 145.680 47.980 145.980 ;
        RECT 46.900 144.800 47.980 145.100 ;
        RECT 47.290 144.220 47.590 144.800 ;
        RECT 46.900 143.920 47.980 144.220 ;
        RECT 46.900 143.340 47.820 143.380 ;
        RECT 46.300 143.040 47.980 143.340 ;
        RECT 42.940 142.160 44.620 142.460 ;
        RECT 46.900 142.460 47.820 142.500 ;
        RECT 46.900 142.160 47.980 142.460 ;
        RECT 40.780 142.020 41.700 142.060 ;
        RECT 40.780 141.720 41.860 142.020 ;
        RECT 48.280 141.580 48.580 147.000 ;
        RECT 49.060 145.240 50.140 145.540 ;
        RECT 49.060 143.480 50.140 143.780 ;
        RECT 50.440 142.020 50.740 154.040 ;
        RECT 49.060 141.720 50.740 142.020 ;
        RECT 42.940 141.280 48.580 141.580 ;
        RECT 42.940 140.700 43.860 140.740 ;
        RECT 46.900 140.700 47.820 140.740 ;
        RECT 42.160 140.400 44.020 140.700 ;
        RECT 46.900 140.400 48.580 140.700 ;
        RECT 42.160 140.260 42.460 140.400 ;
        RECT 35.860 139.960 42.460 140.260 ;
        RECT 30.500 139.820 31.420 139.860 ;
        RECT 34.460 139.820 35.380 139.860 ;
        RECT 35.860 139.820 36.160 139.960 ;
        RECT 29.740 139.520 31.420 139.820 ;
        RECT 34.300 139.520 36.160 139.820 ;
        RECT 38.620 139.010 39.700 139.960 ;
        RECT 42.160 139.820 42.460 139.960 ;
        RECT 48.280 140.260 48.580 140.400 ;
        RECT 51.220 140.260 52.300 210.360 ;
        RECT 54.940 210.220 55.240 210.360 ;
        RECT 61.060 210.660 61.360 210.800 ;
        RECT 63.820 210.660 64.900 211.610 ;
        RECT 68.140 211.100 69.060 211.140 ;
        RECT 72.100 211.100 73.020 211.140 ;
        RECT 67.360 210.800 69.220 211.100 ;
        RECT 72.100 210.800 73.780 211.100 ;
        RECT 67.360 210.660 67.660 210.800 ;
        RECT 61.060 210.360 67.660 210.660 ;
        RECT 55.700 210.220 56.620 210.260 ;
        RECT 59.660 210.220 60.580 210.260 ;
        RECT 61.060 210.220 61.360 210.360 ;
        RECT 54.940 209.920 56.620 210.220 ;
        RECT 59.500 209.920 61.360 210.220 ;
        RECT 55.540 209.340 56.460 209.380 ;
        RECT 55.540 209.040 60.580 209.340 ;
        RECT 53.380 208.600 54.460 208.900 ;
        RECT 61.060 208.600 62.740 208.900 ;
        RECT 55.700 208.460 56.620 208.500 ;
        RECT 59.660 208.460 60.580 208.500 ;
        RECT 55.540 208.160 56.620 208.460 ;
        RECT 59.500 208.160 60.580 208.460 ;
        RECT 59.660 207.580 60.580 207.620 ;
        RECT 55.540 207.280 59.200 207.580 ;
        RECT 59.500 207.280 60.580 207.580 ;
        RECT 53.380 206.840 54.460 207.140 ;
        RECT 58.900 206.700 59.200 207.280 ;
        RECT 61.060 206.700 61.360 208.600 ;
        RECT 61.660 207.140 62.580 207.180 ;
        RECT 61.660 206.840 62.740 207.140 ;
        RECT 55.540 206.400 56.620 206.700 ;
        RECT 58.900 206.400 61.360 206.700 ;
        RECT 55.930 205.820 56.230 206.400 ;
        RECT 58.900 205.820 59.200 206.400 ;
        RECT 55.540 205.520 56.620 205.820 ;
        RECT 58.900 205.520 60.580 205.820 ;
        RECT 53.380 205.080 54.460 205.380 ;
        RECT 61.660 205.080 62.740 205.380 ;
        RECT 55.700 204.940 56.620 204.980 ;
        RECT 59.660 204.940 60.580 204.980 ;
        RECT 55.540 204.640 56.620 204.940 ;
        RECT 59.500 204.640 60.580 204.940 ;
        RECT 61.060 204.780 61.960 205.080 ;
        RECT 61.060 204.060 61.360 204.780 ;
        RECT 55.540 203.760 61.360 204.060 ;
        RECT 53.380 203.320 54.460 203.620 ;
        RECT 61.660 203.320 62.740 203.620 ;
        RECT 55.700 203.180 56.620 203.220 ;
        RECT 59.660 203.180 60.580 203.220 ;
        RECT 55.540 202.880 56.620 203.180 ;
        RECT 59.500 202.880 60.580 203.180 ;
        RECT 61.060 203.020 61.960 203.320 ;
        RECT 55.700 202.300 56.620 202.340 ;
        RECT 61.060 202.300 61.360 203.020 ;
        RECT 55.540 202.000 56.620 202.300 ;
        RECT 58.900 202.000 61.360 202.300 ;
        RECT 53.380 201.560 54.460 201.860 ;
        RECT 58.900 201.420 59.200 202.000 ;
        RECT 61.820 201.860 62.740 201.900 ;
        RECT 61.660 201.560 62.740 201.860 ;
        RECT 55.540 201.120 59.200 201.420 ;
        RECT 59.500 201.120 60.580 201.420 ;
        RECT 58.900 200.540 59.200 201.120 ;
        RECT 59.890 200.540 60.190 201.120 ;
        RECT 55.540 200.240 59.200 200.540 ;
        RECT 59.500 200.240 60.580 200.540 ;
        RECT 53.380 199.800 54.460 200.100 ;
        RECT 61.660 199.800 62.740 200.100 ;
        RECT 55.700 199.660 56.620 199.700 ;
        RECT 59.660 199.660 60.580 199.700 ;
        RECT 55.540 199.360 56.620 199.660 ;
        RECT 59.500 199.360 60.580 199.660 ;
        RECT 55.540 198.480 60.580 198.780 ;
        RECT 62.050 198.340 62.350 199.800 ;
        RECT 53.380 198.040 54.460 198.340 ;
        RECT 61.060 198.040 62.740 198.340 ;
        RECT 55.700 197.900 56.620 197.940 ;
        RECT 59.660 197.900 60.580 197.940 ;
        RECT 55.540 197.600 56.620 197.900 ;
        RECT 59.500 197.600 60.580 197.900 ;
        RECT 61.060 197.020 61.360 198.040 ;
        RECT 55.540 196.720 61.360 197.020 ;
        RECT 53.540 196.580 54.460 196.620 ;
        RECT 53.380 196.280 54.460 196.580 ;
        RECT 61.660 196.280 62.740 196.580 ;
        RECT 55.700 196.140 56.620 196.180 ;
        RECT 59.660 196.140 60.580 196.180 ;
        RECT 55.540 195.840 56.620 196.140 ;
        RECT 59.500 195.840 60.580 196.140 ;
        RECT 59.660 195.260 60.580 195.300 ;
        RECT 55.540 194.960 60.580 195.260 ;
        RECT 53.380 194.520 54.460 194.820 ;
        RECT 53.770 193.100 54.070 194.520 ;
        RECT 55.540 194.080 56.620 194.380 ;
        RECT 55.930 193.500 56.230 194.080 ;
        RECT 55.540 193.200 56.620 193.500 ;
        RECT 53.540 193.060 54.460 193.100 ;
        RECT 53.380 192.760 54.460 193.060 ;
        RECT 55.700 192.620 56.620 192.660 ;
        RECT 55.540 192.320 56.620 192.620 ;
        RECT 55.930 191.780 56.230 192.320 ;
        RECT 55.700 191.740 56.620 191.780 ;
        RECT 55.540 191.440 56.620 191.740 ;
        RECT 53.380 191.000 54.460 191.300 ;
        RECT 53.770 189.540 54.070 191.000 ;
        RECT 55.540 190.560 56.620 190.860 ;
        RECT 55.930 189.980 56.230 190.560 ;
        RECT 55.540 189.680 56.620 189.980 ;
        RECT 53.380 189.240 55.240 189.540 ;
        RECT 53.380 187.480 54.460 187.780 ;
        RECT 53.770 186.020 54.070 187.480 ;
        RECT 53.380 185.720 54.460 186.020 ;
        RECT 53.770 184.260 54.070 185.720 ;
        RECT 53.380 183.960 54.460 184.260 ;
        RECT 53.770 182.500 54.070 183.960 ;
        RECT 54.940 182.940 55.240 189.240 ;
        RECT 58.900 189.100 59.200 194.960 ;
        RECT 61.660 194.520 62.740 194.820 ;
        RECT 59.500 194.080 60.580 194.380 ;
        RECT 59.890 193.500 60.190 194.080 ;
        RECT 59.500 193.200 60.580 193.500 ;
        RECT 62.050 193.060 62.350 194.520 ;
        RECT 61.660 192.760 62.740 193.060 ;
        RECT 59.660 192.620 60.580 192.660 ;
        RECT 59.500 192.320 60.580 192.620 ;
        RECT 59.890 191.780 60.190 192.320 ;
        RECT 59.660 191.740 60.580 191.780 ;
        RECT 59.500 191.440 60.580 191.740 ;
        RECT 62.050 191.340 62.350 192.760 ;
        RECT 61.660 191.300 62.580 191.340 ;
        RECT 61.660 191.000 62.740 191.300 ;
        RECT 59.500 190.560 60.580 190.860 ;
        RECT 59.890 189.980 60.190 190.560 ;
        RECT 59.500 189.680 60.580 189.980 ;
        RECT 62.050 189.540 62.350 191.000 ;
        RECT 61.660 189.240 62.740 189.540 ;
        RECT 59.660 189.100 60.580 189.140 ;
        RECT 55.540 188.800 59.200 189.100 ;
        RECT 59.500 188.800 60.580 189.100 ;
        RECT 55.700 188.220 56.620 188.260 ;
        RECT 59.660 188.220 60.580 188.260 ;
        RECT 55.540 187.920 56.620 188.220 ;
        RECT 59.500 187.920 60.580 188.220 ;
        RECT 61.660 187.480 62.740 187.780 ;
        RECT 55.540 187.040 56.620 187.340 ;
        RECT 59.500 187.040 60.580 187.340 ;
        RECT 55.930 186.460 56.230 187.040 ;
        RECT 59.890 186.460 60.190 187.040 ;
        RECT 55.540 186.160 60.580 186.460 ;
        RECT 55.540 185.280 56.620 185.580 ;
        RECT 55.930 184.740 56.230 185.280 ;
        RECT 55.700 184.700 56.620 184.740 ;
        RECT 55.540 184.400 56.620 184.700 ;
        RECT 55.540 183.520 56.620 183.820 ;
        RECT 55.930 182.940 56.230 183.520 ;
        RECT 57.070 182.940 57.410 183.210 ;
        RECT 58.900 182.940 59.200 186.160 ;
        RECT 62.050 186.020 62.350 187.480 ;
        RECT 61.660 185.720 62.740 186.020 ;
        RECT 59.660 185.580 60.580 185.620 ;
        RECT 59.500 185.280 60.580 185.580 ;
        RECT 59.890 184.740 60.190 185.280 ;
        RECT 59.660 184.700 60.580 184.740 ;
        RECT 59.500 184.400 60.580 184.700 ;
        RECT 62.050 184.260 62.350 185.720 ;
        RECT 61.660 183.960 62.740 184.260 ;
        RECT 59.500 183.520 60.580 183.820 ;
        RECT 59.890 182.940 60.190 183.520 ;
        RECT 54.940 182.640 60.580 182.940 ;
        RECT 53.380 182.200 54.460 182.500 ;
        RECT 57.070 182.290 57.410 182.640 ;
        RECT 62.050 182.500 62.350 183.960 ;
        RECT 61.060 182.200 62.740 182.500 ;
        RECT 55.700 182.060 56.620 182.100 ;
        RECT 59.660 182.060 60.580 182.100 ;
        RECT 55.540 181.760 56.620 182.060 ;
        RECT 59.500 181.760 60.580 182.060 ;
        RECT 55.700 181.180 56.620 181.220 ;
        RECT 59.660 181.180 60.580 181.220 ;
        RECT 55.540 180.880 56.620 181.180 ;
        RECT 59.500 180.880 60.580 181.180 ;
        RECT 53.380 180.440 54.460 180.740 ;
        RECT 53.770 178.980 54.070 180.440 ;
        RECT 55.540 180.000 56.620 180.300 ;
        RECT 59.500 180.000 60.580 180.300 ;
        RECT 55.930 179.420 56.230 180.000 ;
        RECT 59.890 179.420 60.190 180.000 ;
        RECT 55.540 179.120 60.580 179.420 ;
        RECT 53.380 178.680 54.460 178.980 ;
        RECT 53.770 177.220 54.070 178.680 ;
        RECT 55.540 178.240 56.620 178.540 ;
        RECT 55.930 177.700 56.230 178.240 ;
        RECT 55.700 177.660 56.620 177.700 ;
        RECT 55.540 177.360 56.620 177.660 ;
        RECT 53.380 176.920 54.460 177.220 ;
        RECT 53.770 175.460 54.070 176.920 ;
        RECT 55.540 176.480 56.620 176.780 ;
        RECT 55.930 175.900 56.230 176.480 ;
        RECT 57.945 175.900 58.285 176.170 ;
        RECT 58.900 175.900 59.200 179.120 ;
        RECT 59.660 178.540 60.580 178.580 ;
        RECT 59.500 178.240 60.580 178.540 ;
        RECT 59.890 177.700 60.190 178.240 ;
        RECT 59.660 177.660 60.580 177.700 ;
        RECT 59.500 177.360 60.580 177.660 ;
        RECT 59.500 176.480 60.580 176.780 ;
        RECT 59.890 175.900 60.190 176.480 ;
        RECT 61.060 175.900 61.360 182.200 ;
        RECT 61.660 180.440 62.740 180.740 ;
        RECT 62.050 178.980 62.350 180.440 ;
        RECT 61.660 178.680 62.740 178.980 ;
        RECT 62.050 177.220 62.350 178.680 ;
        RECT 61.660 176.920 62.740 177.220 ;
        RECT 55.540 175.600 61.360 175.900 ;
        RECT 53.380 175.160 54.460 175.460 ;
        RECT 57.945 175.250 58.285 175.600 ;
        RECT 62.050 175.500 62.350 176.920 ;
        RECT 61.820 175.460 62.740 175.500 ;
        RECT 61.660 175.160 62.740 175.460 ;
        RECT 55.700 175.020 56.620 175.060 ;
        RECT 59.660 175.020 60.580 175.060 ;
        RECT 55.540 174.720 56.620 175.020 ;
        RECT 59.500 174.720 60.580 175.020 ;
        RECT 55.700 174.140 56.620 174.180 ;
        RECT 59.660 174.140 60.580 174.180 ;
        RECT 55.540 173.840 56.620 174.140 ;
        RECT 59.500 173.840 60.580 174.140 ;
        RECT 53.380 173.400 54.460 173.700 ;
        RECT 61.660 173.400 62.740 173.700 ;
        RECT 53.770 171.940 54.070 173.400 ;
        RECT 55.540 172.960 56.620 173.260 ;
        RECT 59.500 172.960 60.580 173.260 ;
        RECT 55.930 172.380 56.230 172.960 ;
        RECT 59.890 172.380 60.190 172.960 ;
        RECT 55.540 172.080 60.580 172.380 ;
        RECT 53.380 171.640 54.460 171.940 ;
        RECT 53.770 170.180 54.070 171.640 ;
        RECT 55.540 171.200 56.620 171.500 ;
        RECT 55.930 170.660 56.230 171.200 ;
        RECT 55.700 170.620 56.620 170.660 ;
        RECT 55.540 170.320 56.620 170.620 ;
        RECT 53.380 169.880 54.460 170.180 ;
        RECT 53.770 168.420 54.070 169.880 ;
        RECT 55.540 169.440 56.620 169.740 ;
        RECT 55.930 168.900 56.230 169.440 ;
        RECT 58.900 169.130 59.200 172.080 ;
        RECT 62.050 171.940 62.350 173.400 ;
        RECT 61.660 171.640 62.740 171.940 ;
        RECT 59.660 171.500 60.580 171.540 ;
        RECT 59.500 171.200 60.580 171.500 ;
        RECT 59.890 170.660 60.190 171.200 ;
        RECT 59.660 170.620 60.580 170.660 ;
        RECT 59.500 170.320 60.580 170.620 ;
        RECT 62.050 170.180 62.350 171.640 ;
        RECT 61.660 169.880 62.740 170.180 ;
        RECT 59.500 169.440 60.580 169.740 ;
        RECT 55.700 168.860 56.620 168.900 ;
        RECT 58.745 168.860 59.200 169.130 ;
        RECT 59.890 168.860 60.190 169.440 ;
        RECT 55.540 168.560 60.580 168.860 ;
        RECT 53.380 168.120 54.460 168.420 ;
        RECT 58.745 168.210 59.085 168.560 ;
        RECT 62.050 168.420 62.350 169.880 ;
        RECT 61.060 168.120 62.740 168.420 ;
        RECT 55.700 167.980 56.620 168.020 ;
        RECT 59.660 167.980 60.580 168.020 ;
        RECT 55.540 167.680 56.620 167.980 ;
        RECT 59.500 167.680 60.580 167.980 ;
        RECT 55.700 167.100 56.620 167.140 ;
        RECT 59.660 167.100 60.580 167.140 ;
        RECT 55.540 166.800 56.620 167.100 ;
        RECT 59.500 166.800 60.580 167.100 ;
        RECT 53.380 166.360 54.460 166.660 ;
        RECT 53.770 164.900 54.070 166.360 ;
        RECT 55.540 165.920 56.620 166.220 ;
        RECT 59.500 165.920 60.580 166.220 ;
        RECT 55.930 165.340 56.230 165.920 ;
        RECT 59.890 165.340 60.190 165.920 ;
        RECT 55.540 165.040 60.580 165.340 ;
        RECT 53.380 164.600 54.460 164.900 ;
        RECT 53.770 163.140 54.070 164.600 ;
        RECT 55.540 164.160 56.620 164.460 ;
        RECT 55.930 163.620 56.230 164.160 ;
        RECT 55.700 163.580 56.620 163.620 ;
        RECT 55.540 163.280 56.620 163.580 ;
        RECT 53.380 162.840 54.460 163.140 ;
        RECT 53.770 161.380 54.070 162.840 ;
        RECT 55.540 162.400 56.620 162.700 ;
        RECT 55.930 161.820 56.230 162.400 ;
        RECT 58.900 161.820 59.200 165.040 ;
        RECT 59.660 164.460 60.580 164.500 ;
        RECT 59.500 164.160 60.580 164.460 ;
        RECT 59.890 163.620 60.190 164.160 ;
        RECT 59.660 163.580 60.580 163.620 ;
        RECT 59.500 163.280 60.580 163.580 ;
        RECT 59.500 162.400 60.580 162.700 ;
        RECT 59.890 161.820 60.190 162.400 ;
        RECT 61.060 161.820 61.360 168.120 ;
        RECT 61.740 168.080 62.660 168.120 ;
        RECT 61.660 166.360 62.740 166.660 ;
        RECT 62.050 164.900 62.350 166.360 ;
        RECT 61.660 164.600 62.740 164.900 ;
        RECT 62.050 163.140 62.350 164.600 ;
        RECT 61.660 162.840 62.740 163.140 ;
        RECT 55.540 161.520 61.360 161.820 ;
        RECT 62.050 161.380 62.350 162.840 ;
        RECT 53.380 161.080 55.060 161.380 ;
        RECT 61.660 161.080 62.740 161.380 ;
        RECT 54.760 160.060 55.060 161.080 ;
        RECT 55.700 160.940 56.620 160.980 ;
        RECT 59.660 160.940 60.580 160.980 ;
        RECT 55.540 160.640 56.620 160.940 ;
        RECT 59.500 160.640 60.580 160.940 ;
        RECT 54.760 159.760 60.580 160.060 ;
        RECT 53.380 159.620 54.300 159.660 ;
        RECT 61.820 159.620 62.740 159.660 ;
        RECT 52.780 159.320 54.460 159.620 ;
        RECT 61.660 159.320 62.740 159.620 ;
        RECT 52.780 154.340 53.080 159.320 ;
        RECT 53.770 157.860 54.070 159.320 ;
        RECT 55.540 158.880 56.620 159.180 ;
        RECT 59.500 158.880 60.580 159.180 ;
        RECT 55.930 158.300 56.230 158.880 ;
        RECT 59.890 158.300 60.190 158.880 ;
        RECT 55.540 158.000 56.620 158.300 ;
        RECT 59.500 158.000 60.580 158.300 ;
        RECT 53.380 157.560 54.460 157.860 ;
        RECT 61.060 157.560 62.740 157.860 ;
        RECT 53.770 156.100 54.070 157.560 ;
        RECT 55.540 157.120 56.620 157.420 ;
        RECT 59.500 157.120 60.580 157.420 ;
        RECT 55.930 156.540 56.230 157.120 ;
        RECT 59.890 156.540 60.190 157.120 ;
        RECT 55.540 156.240 56.620 156.540 ;
        RECT 59.500 156.240 60.580 156.540 ;
        RECT 53.380 155.800 54.460 156.100 ;
        RECT 55.700 155.660 56.620 155.700 ;
        RECT 59.660 155.660 60.580 155.700 ;
        RECT 55.540 155.360 56.620 155.660 ;
        RECT 59.500 155.360 60.580 155.660 ;
        RECT 59.660 154.780 60.580 154.820 ;
        RECT 55.540 154.480 60.580 154.780 ;
        RECT 52.780 154.040 54.460 154.340 ;
        RECT 52.780 142.020 53.080 154.040 ;
        RECT 53.770 152.580 54.070 154.040 ;
        RECT 55.540 153.600 56.620 153.900 ;
        RECT 59.500 153.600 60.580 153.900 ;
        RECT 55.930 153.020 56.230 153.600 ;
        RECT 59.890 153.020 60.190 153.600 ;
        RECT 55.540 152.720 56.620 153.020 ;
        RECT 59.500 152.720 60.580 153.020 ;
        RECT 61.060 152.580 61.360 157.560 ;
        RECT 61.660 156.100 62.580 156.140 ;
        RECT 61.660 155.800 63.340 156.100 ;
        RECT 61.820 154.340 62.740 154.380 ;
        RECT 61.660 154.040 62.740 154.340 ;
        RECT 53.380 152.280 54.460 152.580 ;
        RECT 61.060 152.280 62.740 152.580 ;
        RECT 53.770 150.820 54.070 152.280 ;
        RECT 55.540 151.840 56.620 152.140 ;
        RECT 59.500 151.840 60.580 152.140 ;
        RECT 55.930 151.260 56.230 151.840 ;
        RECT 59.890 151.260 60.190 151.840 ;
        RECT 55.540 150.960 56.620 151.260 ;
        RECT 59.500 150.960 60.580 151.260 ;
        RECT 53.380 150.520 54.460 150.820 ;
        RECT 55.700 150.380 56.620 150.420 ;
        RECT 59.660 150.380 60.580 150.420 ;
        RECT 55.540 150.080 56.620 150.380 ;
        RECT 59.500 150.080 60.580 150.380 ;
        RECT 61.060 149.500 61.360 152.280 ;
        RECT 61.660 150.820 62.580 150.860 ;
        RECT 61.660 150.520 62.740 150.820 ;
        RECT 55.540 149.200 61.360 149.500 ;
        RECT 53.380 148.760 54.460 149.060 ;
        RECT 61.660 148.760 62.740 149.060 ;
        RECT 55.700 148.620 56.620 148.660 ;
        RECT 59.660 148.620 60.580 148.660 ;
        RECT 55.540 148.320 56.620 148.620 ;
        RECT 59.500 148.320 60.580 148.620 ;
        RECT 61.060 148.460 61.960 148.760 ;
        RECT 55.700 147.740 56.620 147.780 ;
        RECT 61.060 147.740 61.360 148.460 ;
        RECT 55.540 147.440 56.620 147.740 ;
        RECT 56.920 147.440 61.360 147.740 ;
        RECT 53.380 147.000 55.240 147.300 ;
        RECT 53.380 145.240 54.460 145.540 ;
        RECT 53.380 143.480 54.460 143.780 ;
        RECT 52.780 141.720 54.460 142.020 ;
        RECT 54.940 141.580 55.240 147.000 ;
        RECT 55.540 146.560 56.620 146.860 ;
        RECT 55.930 145.980 56.230 146.560 ;
        RECT 55.540 145.680 56.620 145.980 ;
        RECT 55.540 144.800 56.620 145.100 ;
        RECT 55.930 144.220 56.230 144.800 ;
        RECT 55.540 143.920 56.620 144.220 ;
        RECT 55.700 143.340 56.620 143.380 ;
        RECT 56.920 143.340 57.220 147.440 ;
        RECT 61.660 147.000 62.740 147.300 ;
        RECT 59.660 146.860 60.580 146.900 ;
        RECT 59.500 146.560 60.580 146.860 ;
        RECT 59.660 145.980 60.580 146.020 ;
        RECT 59.500 145.680 60.580 145.980 ;
        RECT 61.660 145.540 62.580 145.580 ;
        RECT 61.660 145.240 62.740 145.540 ;
        RECT 55.540 143.040 57.220 143.340 ;
        RECT 58.900 144.800 60.580 145.100 ;
        RECT 58.900 144.220 59.200 144.800 ;
        RECT 58.900 143.920 60.580 144.220 ;
        RECT 55.700 142.460 56.620 142.500 ;
        RECT 55.540 142.160 56.620 142.460 ;
        RECT 58.900 142.460 59.200 143.920 ;
        RECT 63.040 143.780 63.340 155.800 ;
        RECT 61.660 143.480 63.340 143.780 ;
        RECT 59.660 143.340 60.580 143.380 ;
        RECT 59.500 143.040 60.580 143.340 ;
        RECT 58.900 142.160 60.580 142.460 ;
        RECT 61.820 142.020 62.740 142.060 ;
        RECT 61.660 141.720 62.740 142.020 ;
        RECT 54.940 141.280 60.580 141.580 ;
        RECT 55.700 140.700 56.620 140.740 ;
        RECT 59.660 140.700 60.580 140.740 ;
        RECT 54.940 140.400 56.620 140.700 ;
        RECT 59.500 140.400 61.360 140.700 ;
        RECT 54.940 140.260 55.240 140.400 ;
        RECT 48.280 139.960 55.240 140.260 ;
        RECT 42.940 139.820 43.860 139.860 ;
        RECT 46.900 139.820 47.820 139.860 ;
        RECT 48.280 139.820 48.580 139.960 ;
        RECT 42.160 139.520 44.020 139.820 ;
        RECT 46.900 139.520 48.580 139.820 ;
        RECT 51.220 139.010 52.300 139.960 ;
        RECT 54.940 139.820 55.240 139.960 ;
        RECT 61.060 140.260 61.360 140.400 ;
        RECT 63.820 140.260 64.900 210.360 ;
        RECT 67.360 210.220 67.660 210.360 ;
        RECT 73.480 210.660 73.780 210.800 ;
        RECT 76.420 210.660 77.500 211.610 ;
        RECT 80.900 211.100 81.820 211.140 ;
        RECT 84.860 211.100 85.780 211.140 ;
        RECT 80.140 210.800 81.820 211.100 ;
        RECT 84.700 210.800 86.560 211.100 ;
        RECT 80.140 210.660 80.440 210.800 ;
        RECT 73.480 210.360 80.440 210.660 ;
        RECT 68.140 210.220 69.060 210.260 ;
        RECT 72.100 210.220 73.020 210.260 ;
        RECT 73.480 210.220 73.780 210.360 ;
        RECT 67.360 209.920 69.220 210.220 ;
        RECT 72.100 209.920 73.780 210.220 ;
        RECT 72.100 209.340 73.020 209.570 ;
        RECT 68.140 209.040 73.180 209.340 ;
        RECT 65.980 208.600 67.660 208.900 ;
        RECT 74.260 208.600 75.340 208.900 ;
        RECT 65.980 207.140 66.900 207.180 ;
        RECT 65.980 206.840 67.060 207.140 ;
        RECT 67.360 206.700 67.660 208.600 ;
        RECT 68.140 208.460 69.060 208.500 ;
        RECT 72.100 208.460 73.020 208.500 ;
        RECT 68.140 208.160 69.220 208.460 ;
        RECT 72.100 208.160 73.180 208.460 ;
        RECT 68.140 207.580 69.060 207.620 ;
        RECT 68.140 207.280 69.220 207.580 ;
        RECT 69.520 207.280 73.180 207.580 ;
        RECT 69.520 206.700 69.820 207.280 ;
        RECT 74.260 206.840 75.340 207.140 ;
        RECT 67.360 206.400 69.820 206.700 ;
        RECT 72.100 206.400 73.180 206.700 ;
        RECT 69.520 205.820 69.820 206.400 ;
        RECT 72.490 205.820 72.790 206.400 ;
        RECT 68.140 205.520 69.820 205.820 ;
        RECT 72.100 205.520 73.180 205.820 ;
        RECT 65.980 205.080 67.060 205.380 ;
        RECT 74.260 205.080 75.340 205.380 ;
        RECT 66.760 204.780 67.660 205.080 ;
        RECT 67.360 204.060 67.660 204.780 ;
        RECT 68.140 204.940 69.060 204.980 ;
        RECT 72.100 204.940 73.020 204.980 ;
        RECT 68.140 204.640 69.220 204.940 ;
        RECT 72.100 204.640 73.180 204.940 ;
        RECT 67.360 203.760 73.180 204.060 ;
        RECT 65.980 203.320 67.060 203.620 ;
        RECT 74.260 203.320 75.340 203.620 ;
        RECT 66.760 203.020 67.660 203.320 ;
        RECT 67.360 202.300 67.660 203.020 ;
        RECT 68.140 203.180 69.060 203.220 ;
        RECT 72.100 203.180 73.020 203.220 ;
        RECT 68.140 202.880 69.220 203.180 ;
        RECT 72.100 202.880 73.180 203.180 ;
        RECT 72.100 202.300 73.020 202.340 ;
        RECT 67.360 202.000 69.820 202.300 ;
        RECT 72.100 202.000 73.180 202.300 ;
        RECT 65.980 201.860 66.900 201.900 ;
        RECT 65.980 201.560 67.060 201.860 ;
        RECT 69.520 201.420 69.820 202.000 ;
        RECT 74.260 201.560 75.340 201.860 ;
        RECT 68.140 201.120 69.220 201.420 ;
        RECT 69.520 201.120 73.180 201.420 ;
        RECT 68.530 200.540 68.830 201.120 ;
        RECT 69.520 200.540 69.820 201.120 ;
        RECT 68.140 200.240 69.220 200.540 ;
        RECT 69.520 200.240 73.180 200.540 ;
        RECT 65.980 199.800 67.060 200.100 ;
        RECT 74.260 199.800 75.340 200.100 ;
        RECT 66.370 198.340 66.670 199.800 ;
        RECT 68.140 199.660 69.060 199.700 ;
        RECT 72.100 199.660 73.020 199.700 ;
        RECT 68.140 199.360 69.220 199.660 ;
        RECT 72.100 199.360 73.180 199.660 ;
        RECT 68.140 198.480 73.180 198.780 ;
        RECT 65.980 198.040 67.660 198.340 ;
        RECT 74.260 198.040 75.340 198.340 ;
        RECT 67.360 197.020 67.660 198.040 ;
        RECT 68.140 197.900 69.060 197.940 ;
        RECT 72.100 197.900 73.020 197.940 ;
        RECT 68.140 197.600 69.220 197.900 ;
        RECT 72.100 197.600 73.180 197.900 ;
        RECT 67.360 196.720 73.180 197.020 ;
        RECT 74.260 196.580 75.180 196.620 ;
        RECT 65.980 196.280 67.060 196.580 ;
        RECT 74.260 196.280 75.340 196.580 ;
        RECT 68.140 196.140 69.060 196.180 ;
        RECT 72.100 196.140 73.020 196.180 ;
        RECT 68.140 195.840 69.220 196.140 ;
        RECT 72.100 195.840 73.180 196.140 ;
        RECT 68.140 195.260 69.060 195.300 ;
        RECT 68.140 194.960 73.180 195.260 ;
        RECT 65.980 194.520 67.060 194.820 ;
        RECT 66.370 193.060 66.670 194.520 ;
        RECT 68.140 194.080 69.220 194.380 ;
        RECT 68.530 193.500 68.830 194.080 ;
        RECT 68.140 193.200 69.220 193.500 ;
        RECT 65.980 192.760 67.060 193.060 ;
        RECT 66.370 191.340 66.670 192.760 ;
        RECT 68.140 192.620 69.060 192.660 ;
        RECT 68.140 192.320 69.220 192.620 ;
        RECT 68.530 191.780 68.830 192.320 ;
        RECT 68.140 191.740 69.060 191.780 ;
        RECT 68.140 191.440 69.220 191.740 ;
        RECT 65.980 191.300 66.900 191.340 ;
        RECT 65.980 191.000 67.060 191.300 ;
        RECT 66.370 189.540 66.670 191.000 ;
        RECT 68.140 190.560 69.220 190.860 ;
        RECT 68.530 189.980 68.830 190.560 ;
        RECT 68.140 189.680 69.220 189.980 ;
        RECT 65.980 189.240 67.060 189.540 ;
        RECT 68.140 189.100 69.060 189.140 ;
        RECT 69.520 189.100 69.820 194.960 ;
        RECT 74.260 194.520 75.340 194.820 ;
        RECT 72.100 194.080 73.180 194.380 ;
        RECT 72.490 193.500 72.790 194.080 ;
        RECT 72.100 193.200 73.180 193.500 ;
        RECT 74.650 193.100 74.950 194.520 ;
        RECT 74.260 193.060 75.180 193.100 ;
        RECT 74.260 192.760 75.340 193.060 ;
        RECT 72.100 192.620 73.020 192.660 ;
        RECT 72.100 192.320 73.180 192.620 ;
        RECT 72.490 191.780 72.790 192.320 ;
        RECT 72.100 191.740 73.020 191.780 ;
        RECT 72.100 191.440 73.180 191.740 ;
        RECT 74.260 191.000 75.340 191.300 ;
        RECT 72.100 190.560 73.180 190.860 ;
        RECT 72.490 189.980 72.790 190.560 ;
        RECT 72.100 189.680 73.180 189.980 ;
        RECT 74.650 189.540 74.950 191.000 ;
        RECT 73.480 189.240 75.340 189.540 ;
        RECT 68.140 188.800 69.220 189.100 ;
        RECT 69.520 188.800 73.180 189.100 ;
        RECT 68.140 188.220 69.060 188.260 ;
        RECT 72.100 188.220 73.020 188.260 ;
        RECT 68.140 187.920 69.220 188.220 ;
        RECT 72.100 187.920 73.180 188.220 ;
        RECT 65.980 187.480 67.060 187.780 ;
        RECT 66.370 186.020 66.670 187.480 ;
        RECT 68.140 187.040 69.220 187.340 ;
        RECT 72.100 187.040 73.180 187.340 ;
        RECT 68.530 186.460 68.830 187.040 ;
        RECT 72.490 186.460 72.790 187.040 ;
        RECT 68.140 186.160 73.180 186.460 ;
        RECT 65.980 185.720 67.060 186.020 ;
        RECT 66.370 184.260 66.670 185.720 ;
        RECT 68.140 185.580 69.060 185.620 ;
        RECT 68.140 185.280 69.220 185.580 ;
        RECT 68.530 184.740 68.830 185.280 ;
        RECT 68.140 184.700 69.060 184.740 ;
        RECT 68.140 184.400 69.220 184.700 ;
        RECT 65.980 183.960 67.060 184.260 ;
        RECT 66.370 182.500 66.670 183.960 ;
        RECT 68.140 183.520 69.220 183.820 ;
        RECT 68.530 182.940 68.830 183.520 ;
        RECT 69.520 182.940 69.820 186.160 ;
        RECT 72.100 185.280 73.180 185.580 ;
        RECT 72.490 184.740 72.790 185.280 ;
        RECT 72.100 184.700 73.020 184.740 ;
        RECT 72.100 184.400 73.180 184.700 ;
        RECT 72.100 183.520 73.180 183.820 ;
        RECT 71.310 182.940 71.650 183.210 ;
        RECT 72.490 182.940 72.790 183.520 ;
        RECT 73.480 182.940 73.780 189.240 ;
        RECT 74.260 187.480 75.340 187.780 ;
        RECT 74.650 186.020 74.950 187.480 ;
        RECT 74.260 185.720 75.340 186.020 ;
        RECT 74.650 184.260 74.950 185.720 ;
        RECT 74.260 183.960 75.340 184.260 ;
        RECT 68.140 182.640 73.780 182.940 ;
        RECT 65.980 182.200 67.660 182.500 ;
        RECT 71.310 182.290 71.650 182.640 ;
        RECT 74.650 182.500 74.950 183.960 ;
        RECT 74.260 182.200 75.340 182.500 ;
        RECT 65.980 180.440 67.060 180.740 ;
        RECT 66.370 178.980 66.670 180.440 ;
        RECT 65.980 178.680 67.060 178.980 ;
        RECT 66.370 177.220 66.670 178.680 ;
        RECT 65.980 176.920 67.060 177.220 ;
        RECT 66.370 175.500 66.670 176.920 ;
        RECT 67.360 175.900 67.660 182.200 ;
        RECT 68.140 182.060 69.060 182.100 ;
        RECT 72.100 182.060 73.020 182.100 ;
        RECT 68.140 181.760 69.220 182.060 ;
        RECT 72.100 181.760 73.180 182.060 ;
        RECT 68.140 181.180 69.060 181.220 ;
        RECT 72.100 181.180 73.020 181.220 ;
        RECT 68.140 180.880 69.220 181.180 ;
        RECT 72.100 180.880 73.180 181.180 ;
        RECT 74.260 180.440 75.340 180.740 ;
        RECT 68.140 180.000 69.220 180.300 ;
        RECT 72.100 180.000 73.180 180.300 ;
        RECT 68.530 179.420 68.830 180.000 ;
        RECT 72.490 179.420 72.790 180.000 ;
        RECT 68.140 179.120 73.180 179.420 ;
        RECT 68.140 178.540 69.060 178.580 ;
        RECT 68.140 178.240 69.220 178.540 ;
        RECT 68.530 177.700 68.830 178.240 ;
        RECT 68.140 177.660 69.060 177.700 ;
        RECT 68.140 177.360 69.220 177.660 ;
        RECT 68.140 176.480 69.220 176.780 ;
        RECT 68.530 175.900 68.830 176.480 ;
        RECT 69.520 175.900 69.820 179.120 ;
        RECT 74.650 178.980 74.950 180.440 ;
        RECT 74.260 178.680 75.340 178.980 ;
        RECT 72.100 178.240 73.180 178.540 ;
        RECT 72.490 177.700 72.790 178.240 ;
        RECT 72.100 177.660 73.020 177.700 ;
        RECT 72.100 177.360 73.180 177.660 ;
        RECT 74.650 177.220 74.950 178.680 ;
        RECT 74.260 176.920 75.340 177.220 ;
        RECT 72.100 176.480 73.180 176.780 ;
        RECT 70.435 175.900 70.775 176.170 ;
        RECT 72.490 175.900 72.790 176.480 ;
        RECT 67.360 175.600 73.180 175.900 ;
        RECT 65.980 175.460 66.900 175.500 ;
        RECT 65.980 175.160 67.060 175.460 ;
        RECT 70.435 175.250 70.775 175.600 ;
        RECT 74.650 175.460 74.950 176.920 ;
        RECT 74.260 175.160 75.340 175.460 ;
        RECT 68.140 175.020 69.060 175.060 ;
        RECT 72.100 175.020 73.020 175.060 ;
        RECT 68.140 174.720 69.220 175.020 ;
        RECT 72.100 174.720 73.180 175.020 ;
        RECT 68.140 174.140 69.060 174.180 ;
        RECT 72.100 174.140 73.020 174.180 ;
        RECT 68.140 173.840 69.220 174.140 ;
        RECT 72.100 173.840 73.180 174.140 ;
        RECT 65.980 173.400 67.060 173.700 ;
        RECT 74.260 173.400 75.340 173.700 ;
        RECT 66.370 171.940 66.670 173.400 ;
        RECT 68.140 172.960 69.220 173.260 ;
        RECT 72.100 172.960 73.180 173.260 ;
        RECT 68.530 172.380 68.830 172.960 ;
        RECT 72.490 172.380 72.790 172.960 ;
        RECT 68.140 172.080 73.180 172.380 ;
        RECT 65.980 171.640 67.060 171.940 ;
        RECT 66.370 170.180 66.670 171.640 ;
        RECT 68.140 171.500 69.060 171.540 ;
        RECT 68.140 171.200 69.220 171.500 ;
        RECT 68.530 170.660 68.830 171.200 ;
        RECT 68.140 170.620 69.060 170.660 ;
        RECT 68.140 170.320 69.220 170.620 ;
        RECT 65.980 169.880 67.060 170.180 ;
        RECT 66.370 168.420 66.670 169.880 ;
        RECT 68.140 169.440 69.220 169.740 ;
        RECT 68.530 168.860 68.830 169.440 ;
        RECT 69.520 169.130 69.820 172.080 ;
        RECT 74.650 171.940 74.950 173.400 ;
        RECT 74.260 171.640 75.340 171.940 ;
        RECT 72.100 171.200 73.180 171.500 ;
        RECT 72.490 170.660 72.790 171.200 ;
        RECT 72.100 170.620 73.020 170.660 ;
        RECT 72.100 170.320 73.180 170.620 ;
        RECT 74.650 170.180 74.950 171.640 ;
        RECT 74.260 169.880 75.340 170.180 ;
        RECT 72.100 169.440 73.180 169.740 ;
        RECT 69.520 168.860 69.975 169.130 ;
        RECT 72.490 168.900 72.790 169.440 ;
        RECT 72.100 168.860 73.020 168.900 ;
        RECT 68.140 168.560 73.180 168.860 ;
        RECT 65.980 168.120 67.660 168.420 ;
        RECT 69.635 168.210 69.975 168.560 ;
        RECT 74.650 168.420 74.950 169.880 ;
        RECT 74.260 168.120 75.340 168.420 ;
        RECT 66.060 168.080 66.980 168.120 ;
        RECT 65.980 166.360 67.060 166.660 ;
        RECT 66.370 164.900 66.670 166.360 ;
        RECT 65.980 164.600 67.060 164.900 ;
        RECT 66.370 163.140 66.670 164.600 ;
        RECT 65.980 162.840 67.060 163.140 ;
        RECT 66.370 161.380 66.670 162.840 ;
        RECT 67.360 161.820 67.660 168.120 ;
        RECT 68.140 167.980 69.060 168.020 ;
        RECT 72.100 167.980 73.020 168.020 ;
        RECT 68.140 167.680 69.220 167.980 ;
        RECT 72.100 167.680 73.180 167.980 ;
        RECT 68.140 167.100 69.060 167.140 ;
        RECT 72.100 167.100 73.020 167.140 ;
        RECT 68.140 166.800 69.220 167.100 ;
        RECT 72.100 166.800 73.180 167.100 ;
        RECT 74.260 166.360 75.340 166.660 ;
        RECT 68.140 165.920 69.220 166.220 ;
        RECT 72.100 165.920 73.180 166.220 ;
        RECT 68.530 165.340 68.830 165.920 ;
        RECT 72.490 165.340 72.790 165.920 ;
        RECT 68.140 165.040 73.180 165.340 ;
        RECT 68.140 164.460 69.060 164.500 ;
        RECT 68.140 164.160 69.220 164.460 ;
        RECT 68.530 163.620 68.830 164.160 ;
        RECT 68.140 163.580 69.060 163.620 ;
        RECT 68.140 163.280 69.220 163.580 ;
        RECT 68.140 162.400 69.220 162.700 ;
        RECT 68.530 161.820 68.830 162.400 ;
        RECT 69.520 161.820 69.820 165.040 ;
        RECT 74.650 164.900 74.950 166.360 ;
        RECT 74.260 164.600 75.340 164.900 ;
        RECT 72.100 164.160 73.180 164.460 ;
        RECT 72.490 163.620 72.790 164.160 ;
        RECT 72.100 163.580 73.020 163.620 ;
        RECT 72.100 163.280 73.180 163.580 ;
        RECT 74.650 163.140 74.950 164.600 ;
        RECT 74.260 162.840 75.340 163.140 ;
        RECT 72.100 162.400 73.180 162.700 ;
        RECT 72.490 161.820 72.790 162.400 ;
        RECT 67.360 161.520 73.180 161.820 ;
        RECT 74.650 161.380 74.950 162.840 ;
        RECT 65.980 161.080 67.060 161.380 ;
        RECT 73.660 161.080 75.340 161.380 ;
        RECT 68.140 160.940 69.060 160.980 ;
        RECT 72.100 160.940 73.020 160.980 ;
        RECT 68.140 160.640 69.220 160.940 ;
        RECT 72.100 160.640 73.180 160.940 ;
        RECT 73.660 160.060 73.960 161.080 ;
        RECT 68.140 159.760 73.960 160.060 ;
        RECT 65.980 159.620 66.900 159.660 ;
        RECT 74.260 159.620 75.180 159.660 ;
        RECT 65.980 159.320 67.060 159.620 ;
        RECT 74.260 159.320 75.940 159.620 ;
        RECT 68.140 158.880 69.220 159.180 ;
        RECT 72.100 158.880 73.180 159.180 ;
        RECT 68.530 158.300 68.830 158.880 ;
        RECT 72.490 158.300 72.790 158.880 ;
        RECT 68.140 158.000 69.220 158.300 ;
        RECT 72.100 158.000 73.180 158.300 ;
        RECT 74.650 157.860 74.950 159.320 ;
        RECT 65.980 157.560 67.660 157.860 ;
        RECT 74.260 157.560 75.340 157.860 ;
        RECT 65.980 156.100 66.900 156.140 ;
        RECT 65.380 155.800 67.060 156.100 ;
        RECT 65.380 143.780 65.680 155.800 ;
        RECT 65.980 154.340 66.900 154.380 ;
        RECT 65.980 154.040 67.060 154.340 ;
        RECT 67.360 152.580 67.660 157.560 ;
        RECT 68.140 157.120 69.220 157.420 ;
        RECT 72.100 157.120 73.180 157.420 ;
        RECT 68.530 156.540 68.830 157.120 ;
        RECT 72.490 156.540 72.790 157.120 ;
        RECT 68.140 156.240 69.220 156.540 ;
        RECT 72.100 156.240 73.180 156.540 ;
        RECT 74.650 156.100 74.950 157.560 ;
        RECT 74.260 155.800 75.340 156.100 ;
        RECT 68.140 155.660 69.060 155.700 ;
        RECT 72.100 155.660 73.020 155.700 ;
        RECT 68.140 155.360 69.220 155.660 ;
        RECT 72.100 155.360 73.180 155.660 ;
        RECT 68.140 154.780 69.060 154.820 ;
        RECT 68.140 154.480 73.180 154.780 ;
        RECT 75.640 154.340 75.940 159.320 ;
        RECT 74.260 154.040 75.940 154.340 ;
        RECT 68.140 153.600 69.220 153.900 ;
        RECT 72.100 153.600 73.180 153.900 ;
        RECT 68.530 153.020 68.830 153.600 ;
        RECT 72.490 153.020 72.790 153.600 ;
        RECT 68.140 152.720 69.220 153.020 ;
        RECT 72.100 152.720 73.180 153.020 ;
        RECT 74.650 152.580 74.950 154.040 ;
        RECT 65.980 152.280 67.660 152.580 ;
        RECT 74.260 152.280 75.340 152.580 ;
        RECT 66.140 150.820 67.060 150.860 ;
        RECT 65.980 150.520 67.060 150.820 ;
        RECT 67.360 149.500 67.660 152.280 ;
        RECT 68.140 151.840 69.220 152.140 ;
        RECT 72.100 151.840 73.180 152.140 ;
        RECT 68.530 151.260 68.830 151.840 ;
        RECT 72.490 151.260 72.790 151.840 ;
        RECT 68.140 150.960 69.220 151.260 ;
        RECT 72.100 150.960 73.180 151.260 ;
        RECT 74.650 150.820 74.950 152.280 ;
        RECT 74.260 150.520 75.340 150.820 ;
        RECT 68.140 150.380 69.060 150.420 ;
        RECT 72.100 150.380 73.020 150.420 ;
        RECT 68.140 150.080 69.220 150.380 ;
        RECT 72.100 150.080 73.180 150.380 ;
        RECT 67.360 149.200 73.180 149.500 ;
        RECT 65.980 148.760 67.060 149.060 ;
        RECT 74.260 148.760 75.340 149.060 ;
        RECT 66.760 148.460 67.660 148.760 ;
        RECT 67.360 147.740 67.660 148.460 ;
        RECT 68.140 148.620 69.060 148.660 ;
        RECT 72.100 148.620 73.020 148.660 ;
        RECT 68.140 148.320 69.220 148.620 ;
        RECT 72.100 148.320 73.180 148.620 ;
        RECT 72.100 147.740 73.020 147.780 ;
        RECT 67.360 147.440 71.800 147.740 ;
        RECT 72.100 147.440 73.180 147.740 ;
        RECT 65.980 147.000 67.060 147.300 ;
        RECT 68.140 146.860 69.060 146.900 ;
        RECT 68.140 146.560 69.220 146.860 ;
        RECT 68.140 145.980 69.060 146.020 ;
        RECT 68.140 145.680 69.220 145.980 ;
        RECT 66.140 145.540 67.060 145.580 ;
        RECT 65.980 145.240 67.060 145.540 ;
        RECT 68.140 144.800 69.820 145.100 ;
        RECT 69.520 144.220 69.820 144.800 ;
        RECT 68.140 143.920 69.820 144.220 ;
        RECT 65.380 143.480 67.060 143.780 ;
        RECT 68.140 143.340 69.060 143.380 ;
        RECT 68.140 143.040 69.220 143.340 ;
        RECT 69.520 142.460 69.820 143.920 ;
        RECT 71.500 143.340 71.800 147.440 ;
        RECT 73.480 147.000 75.340 147.300 ;
        RECT 72.100 146.560 73.180 146.860 ;
        RECT 72.490 145.980 72.790 146.560 ;
        RECT 72.100 145.680 73.180 145.980 ;
        RECT 72.100 144.800 73.180 145.100 ;
        RECT 72.490 144.220 72.790 144.800 ;
        RECT 72.100 143.920 73.180 144.220 ;
        RECT 72.100 143.340 73.020 143.380 ;
        RECT 71.500 143.040 73.180 143.340 ;
        RECT 68.140 142.160 69.820 142.460 ;
        RECT 72.100 142.460 73.020 142.500 ;
        RECT 72.100 142.160 73.180 142.460 ;
        RECT 65.980 142.020 66.900 142.060 ;
        RECT 65.980 141.720 67.060 142.020 ;
        RECT 73.480 141.580 73.780 147.000 ;
        RECT 74.260 145.240 75.340 145.540 ;
        RECT 74.260 143.480 75.340 143.780 ;
        RECT 75.640 142.020 75.940 154.040 ;
        RECT 74.260 141.720 75.940 142.020 ;
        RECT 68.140 141.280 73.780 141.580 ;
        RECT 68.140 140.700 69.060 140.740 ;
        RECT 72.100 140.700 73.020 140.740 ;
        RECT 67.360 140.400 69.220 140.700 ;
        RECT 72.100 140.400 73.780 140.700 ;
        RECT 67.360 140.260 67.660 140.400 ;
        RECT 61.060 139.960 67.660 140.260 ;
        RECT 55.700 139.820 56.620 139.860 ;
        RECT 59.660 139.820 60.580 139.860 ;
        RECT 61.060 139.820 61.360 139.960 ;
        RECT 54.940 139.520 56.620 139.820 ;
        RECT 59.500 139.520 61.360 139.820 ;
        RECT 63.820 139.010 64.900 139.960 ;
        RECT 67.360 139.820 67.660 139.960 ;
        RECT 73.480 140.260 73.780 140.400 ;
        RECT 76.420 140.260 77.500 210.360 ;
        RECT 80.140 210.220 80.440 210.360 ;
        RECT 86.260 210.660 86.560 210.800 ;
        RECT 89.020 210.660 90.100 211.610 ;
        RECT 93.340 211.100 94.260 211.140 ;
        RECT 97.300 211.100 98.220 211.140 ;
        RECT 92.560 210.800 94.420 211.100 ;
        RECT 97.300 210.800 98.980 211.100 ;
        RECT 92.560 210.660 92.860 210.800 ;
        RECT 86.260 210.360 92.860 210.660 ;
        RECT 80.900 210.220 81.820 210.260 ;
        RECT 84.860 210.220 85.780 210.260 ;
        RECT 86.260 210.220 86.560 210.360 ;
        RECT 80.140 209.920 81.820 210.220 ;
        RECT 84.700 209.920 86.560 210.220 ;
        RECT 80.740 209.340 81.660 209.380 ;
        RECT 80.740 209.040 85.780 209.340 ;
        RECT 78.580 208.600 79.660 208.900 ;
        RECT 86.260 208.600 87.940 208.900 ;
        RECT 80.900 208.460 81.820 208.500 ;
        RECT 84.860 208.460 85.780 208.500 ;
        RECT 80.740 208.160 81.820 208.460 ;
        RECT 84.700 208.160 85.780 208.460 ;
        RECT 84.860 207.580 85.780 207.620 ;
        RECT 80.740 207.280 84.400 207.580 ;
        RECT 84.700 207.280 85.780 207.580 ;
        RECT 78.580 206.840 79.660 207.140 ;
        RECT 84.100 206.700 84.400 207.280 ;
        RECT 86.260 206.700 86.560 208.600 ;
        RECT 86.860 207.140 87.780 207.180 ;
        RECT 86.860 206.840 87.940 207.140 ;
        RECT 80.740 206.400 81.820 206.700 ;
        RECT 84.100 206.400 86.560 206.700 ;
        RECT 81.130 205.820 81.430 206.400 ;
        RECT 84.100 205.820 84.400 206.400 ;
        RECT 80.740 205.520 81.820 205.820 ;
        RECT 84.100 205.520 85.780 205.820 ;
        RECT 78.580 205.080 79.660 205.380 ;
        RECT 86.860 205.080 87.940 205.380 ;
        RECT 80.900 204.940 81.820 204.980 ;
        RECT 84.860 204.940 85.780 204.980 ;
        RECT 80.740 204.640 81.820 204.940 ;
        RECT 84.700 204.640 85.780 204.940 ;
        RECT 86.260 204.780 87.160 205.080 ;
        RECT 86.260 204.060 86.560 204.780 ;
        RECT 80.740 203.760 86.560 204.060 ;
        RECT 78.580 203.320 79.660 203.620 ;
        RECT 86.860 203.320 87.940 203.620 ;
        RECT 80.900 203.180 81.820 203.220 ;
        RECT 84.860 203.180 85.780 203.220 ;
        RECT 80.740 202.880 81.820 203.180 ;
        RECT 84.700 202.880 85.780 203.180 ;
        RECT 86.260 203.020 87.160 203.320 ;
        RECT 80.900 202.300 81.820 202.340 ;
        RECT 86.260 202.300 86.560 203.020 ;
        RECT 80.740 202.000 81.820 202.300 ;
        RECT 84.100 202.000 86.560 202.300 ;
        RECT 78.580 201.560 79.660 201.860 ;
        RECT 84.100 201.420 84.400 202.000 ;
        RECT 87.020 201.860 87.940 201.900 ;
        RECT 86.860 201.560 87.940 201.860 ;
        RECT 80.740 201.120 84.400 201.420 ;
        RECT 84.700 201.120 85.780 201.420 ;
        RECT 84.100 200.540 84.400 201.120 ;
        RECT 85.090 200.540 85.390 201.120 ;
        RECT 80.740 200.240 84.400 200.540 ;
        RECT 84.700 200.240 85.780 200.540 ;
        RECT 78.580 199.800 79.660 200.100 ;
        RECT 86.860 199.800 87.940 200.100 ;
        RECT 80.900 199.660 81.820 199.700 ;
        RECT 84.860 199.660 85.780 199.700 ;
        RECT 80.740 199.360 81.820 199.660 ;
        RECT 84.700 199.360 85.780 199.660 ;
        RECT 80.740 198.480 85.780 198.780 ;
        RECT 87.250 198.340 87.550 199.800 ;
        RECT 78.580 198.040 79.660 198.340 ;
        RECT 86.260 198.040 87.940 198.340 ;
        RECT 80.900 197.900 81.820 197.940 ;
        RECT 84.860 197.900 85.780 197.940 ;
        RECT 80.740 197.600 81.820 197.900 ;
        RECT 84.700 197.600 85.780 197.900 ;
        RECT 86.260 197.020 86.560 198.040 ;
        RECT 80.740 196.720 86.560 197.020 ;
        RECT 78.740 196.580 79.660 196.620 ;
        RECT 78.580 196.280 79.660 196.580 ;
        RECT 86.860 196.280 87.940 196.580 ;
        RECT 80.900 196.140 81.820 196.180 ;
        RECT 84.860 196.140 85.780 196.180 ;
        RECT 80.740 195.840 81.820 196.140 ;
        RECT 84.700 195.840 85.780 196.140 ;
        RECT 84.860 195.260 85.780 195.300 ;
        RECT 80.740 194.960 85.780 195.260 ;
        RECT 78.580 194.520 79.660 194.820 ;
        RECT 78.970 193.100 79.270 194.520 ;
        RECT 80.740 194.080 81.820 194.380 ;
        RECT 81.130 193.500 81.430 194.080 ;
        RECT 80.740 193.200 81.820 193.500 ;
        RECT 78.740 193.060 79.660 193.100 ;
        RECT 78.580 192.760 79.660 193.060 ;
        RECT 80.900 192.620 81.820 192.660 ;
        RECT 80.740 192.320 81.820 192.620 ;
        RECT 81.130 191.780 81.430 192.320 ;
        RECT 80.900 191.740 81.820 191.780 ;
        RECT 80.740 191.440 81.820 191.740 ;
        RECT 78.580 191.000 79.660 191.300 ;
        RECT 78.970 189.540 79.270 191.000 ;
        RECT 80.740 190.560 81.820 190.860 ;
        RECT 81.130 189.980 81.430 190.560 ;
        RECT 80.740 189.680 81.820 189.980 ;
        RECT 78.580 189.240 80.440 189.540 ;
        RECT 78.580 187.480 79.660 187.780 ;
        RECT 78.970 186.020 79.270 187.480 ;
        RECT 78.580 185.720 79.660 186.020 ;
        RECT 78.970 184.260 79.270 185.720 ;
        RECT 78.580 183.960 79.660 184.260 ;
        RECT 78.970 182.500 79.270 183.960 ;
        RECT 80.140 182.940 80.440 189.240 ;
        RECT 84.100 189.100 84.400 194.960 ;
        RECT 86.860 194.520 87.940 194.820 ;
        RECT 84.700 194.080 85.780 194.380 ;
        RECT 85.090 193.500 85.390 194.080 ;
        RECT 84.700 193.200 85.780 193.500 ;
        RECT 87.250 193.060 87.550 194.520 ;
        RECT 86.860 192.760 87.940 193.060 ;
        RECT 84.860 192.620 85.780 192.660 ;
        RECT 84.700 192.320 85.780 192.620 ;
        RECT 85.090 191.780 85.390 192.320 ;
        RECT 84.860 191.740 85.780 191.780 ;
        RECT 84.700 191.440 85.780 191.740 ;
        RECT 87.250 191.340 87.550 192.760 ;
        RECT 86.860 191.300 87.780 191.340 ;
        RECT 86.860 191.000 87.940 191.300 ;
        RECT 84.700 190.560 85.780 190.860 ;
        RECT 85.090 189.980 85.390 190.560 ;
        RECT 84.700 189.680 85.780 189.980 ;
        RECT 87.250 189.540 87.550 191.000 ;
        RECT 86.860 189.240 87.940 189.540 ;
        RECT 84.860 189.100 85.780 189.140 ;
        RECT 80.740 188.800 84.400 189.100 ;
        RECT 84.700 188.800 85.780 189.100 ;
        RECT 80.900 188.220 81.820 188.260 ;
        RECT 84.860 188.220 85.780 188.260 ;
        RECT 80.740 187.920 81.820 188.220 ;
        RECT 84.700 187.920 85.780 188.220 ;
        RECT 86.860 187.480 87.940 187.780 ;
        RECT 80.740 187.040 81.820 187.340 ;
        RECT 84.700 187.040 85.780 187.340 ;
        RECT 81.130 186.460 81.430 187.040 ;
        RECT 85.090 186.460 85.390 187.040 ;
        RECT 80.740 186.160 85.780 186.460 ;
        RECT 80.740 185.280 81.820 185.580 ;
        RECT 81.130 184.740 81.430 185.280 ;
        RECT 80.900 184.700 81.820 184.740 ;
        RECT 80.740 184.400 81.820 184.700 ;
        RECT 80.740 183.520 81.820 183.820 ;
        RECT 81.130 182.940 81.430 183.520 ;
        RECT 82.270 182.940 82.610 183.210 ;
        RECT 84.100 182.940 84.400 186.160 ;
        RECT 87.250 186.020 87.550 187.480 ;
        RECT 86.860 185.720 87.940 186.020 ;
        RECT 84.860 185.580 85.780 185.620 ;
        RECT 84.700 185.280 85.780 185.580 ;
        RECT 85.090 184.740 85.390 185.280 ;
        RECT 84.860 184.700 85.780 184.740 ;
        RECT 84.700 184.400 85.780 184.700 ;
        RECT 87.250 184.260 87.550 185.720 ;
        RECT 86.860 183.960 87.940 184.260 ;
        RECT 84.700 183.520 85.780 183.820 ;
        RECT 85.090 182.940 85.390 183.520 ;
        RECT 80.140 182.640 85.780 182.940 ;
        RECT 78.580 182.200 79.660 182.500 ;
        RECT 82.270 182.290 82.610 182.640 ;
        RECT 87.250 182.500 87.550 183.960 ;
        RECT 86.260 182.200 87.940 182.500 ;
        RECT 80.900 182.060 81.820 182.100 ;
        RECT 84.860 182.060 85.780 182.100 ;
        RECT 80.740 181.760 81.820 182.060 ;
        RECT 84.700 181.760 85.780 182.060 ;
        RECT 80.900 181.180 81.820 181.220 ;
        RECT 84.860 181.180 85.780 181.220 ;
        RECT 80.740 180.880 81.820 181.180 ;
        RECT 84.700 180.880 85.780 181.180 ;
        RECT 78.580 180.440 79.660 180.740 ;
        RECT 78.970 178.980 79.270 180.440 ;
        RECT 80.740 180.000 81.820 180.300 ;
        RECT 84.700 180.000 85.780 180.300 ;
        RECT 81.130 179.420 81.430 180.000 ;
        RECT 85.090 179.420 85.390 180.000 ;
        RECT 80.740 179.120 85.780 179.420 ;
        RECT 78.580 178.680 79.660 178.980 ;
        RECT 78.970 177.220 79.270 178.680 ;
        RECT 80.740 178.240 81.820 178.540 ;
        RECT 81.130 177.700 81.430 178.240 ;
        RECT 80.900 177.660 81.820 177.700 ;
        RECT 80.740 177.360 81.820 177.660 ;
        RECT 78.580 176.920 79.660 177.220 ;
        RECT 78.970 175.460 79.270 176.920 ;
        RECT 80.740 176.480 81.820 176.780 ;
        RECT 81.130 175.900 81.430 176.480 ;
        RECT 83.145 175.900 83.485 176.170 ;
        RECT 84.100 175.900 84.400 179.120 ;
        RECT 84.860 178.540 85.780 178.580 ;
        RECT 84.700 178.240 85.780 178.540 ;
        RECT 85.090 177.700 85.390 178.240 ;
        RECT 84.860 177.660 85.780 177.700 ;
        RECT 84.700 177.360 85.780 177.660 ;
        RECT 84.700 176.480 85.780 176.780 ;
        RECT 85.090 175.900 85.390 176.480 ;
        RECT 86.260 175.900 86.560 182.200 ;
        RECT 86.860 180.440 87.940 180.740 ;
        RECT 87.250 178.980 87.550 180.440 ;
        RECT 86.860 178.680 87.940 178.980 ;
        RECT 87.250 177.220 87.550 178.680 ;
        RECT 86.860 176.920 87.940 177.220 ;
        RECT 80.740 175.600 86.560 175.900 ;
        RECT 78.580 175.160 79.660 175.460 ;
        RECT 83.145 175.250 83.485 175.600 ;
        RECT 87.250 175.500 87.550 176.920 ;
        RECT 87.020 175.460 87.940 175.500 ;
        RECT 86.860 175.160 87.940 175.460 ;
        RECT 80.900 175.020 81.820 175.060 ;
        RECT 84.860 175.020 85.780 175.060 ;
        RECT 80.740 174.720 81.820 175.020 ;
        RECT 84.700 174.720 85.780 175.020 ;
        RECT 80.900 174.140 81.820 174.180 ;
        RECT 84.860 174.140 85.780 174.180 ;
        RECT 80.740 173.840 81.820 174.140 ;
        RECT 84.700 173.840 85.780 174.140 ;
        RECT 78.580 173.400 79.660 173.700 ;
        RECT 86.860 173.400 87.940 173.700 ;
        RECT 78.970 171.940 79.270 173.400 ;
        RECT 80.740 172.960 81.820 173.260 ;
        RECT 84.700 172.960 85.780 173.260 ;
        RECT 81.130 172.380 81.430 172.960 ;
        RECT 85.090 172.380 85.390 172.960 ;
        RECT 80.740 172.080 85.780 172.380 ;
        RECT 78.580 171.640 79.660 171.940 ;
        RECT 78.970 170.180 79.270 171.640 ;
        RECT 80.740 171.200 81.820 171.500 ;
        RECT 81.130 170.660 81.430 171.200 ;
        RECT 80.900 170.620 81.820 170.660 ;
        RECT 80.740 170.320 81.820 170.620 ;
        RECT 78.580 169.880 79.660 170.180 ;
        RECT 78.970 168.420 79.270 169.880 ;
        RECT 80.740 169.440 81.820 169.740 ;
        RECT 81.130 168.900 81.430 169.440 ;
        RECT 84.100 169.130 84.400 172.080 ;
        RECT 87.250 171.940 87.550 173.400 ;
        RECT 86.860 171.640 87.940 171.940 ;
        RECT 84.860 171.500 85.780 171.540 ;
        RECT 84.700 171.200 85.780 171.500 ;
        RECT 85.090 170.660 85.390 171.200 ;
        RECT 84.860 170.620 85.780 170.660 ;
        RECT 84.700 170.320 85.780 170.620 ;
        RECT 87.250 170.180 87.550 171.640 ;
        RECT 86.860 169.880 87.940 170.180 ;
        RECT 84.700 169.440 85.780 169.740 ;
        RECT 80.900 168.860 81.820 168.900 ;
        RECT 83.945 168.860 84.400 169.130 ;
        RECT 85.090 168.860 85.390 169.440 ;
        RECT 80.740 168.560 85.780 168.860 ;
        RECT 78.580 168.120 79.660 168.420 ;
        RECT 83.945 168.210 84.285 168.560 ;
        RECT 87.250 168.420 87.550 169.880 ;
        RECT 86.260 168.120 87.940 168.420 ;
        RECT 80.900 167.980 81.820 168.020 ;
        RECT 84.860 167.980 85.780 168.020 ;
        RECT 80.740 167.680 81.820 167.980 ;
        RECT 84.700 167.680 85.780 167.980 ;
        RECT 80.900 167.100 81.820 167.140 ;
        RECT 84.860 167.100 85.780 167.140 ;
        RECT 80.740 166.800 81.820 167.100 ;
        RECT 84.700 166.800 85.780 167.100 ;
        RECT 78.580 166.360 79.660 166.660 ;
        RECT 78.970 164.900 79.270 166.360 ;
        RECT 80.740 165.920 81.820 166.220 ;
        RECT 84.700 165.920 85.780 166.220 ;
        RECT 81.130 165.340 81.430 165.920 ;
        RECT 85.090 165.340 85.390 165.920 ;
        RECT 80.740 165.040 85.780 165.340 ;
        RECT 78.580 164.600 79.660 164.900 ;
        RECT 78.970 163.140 79.270 164.600 ;
        RECT 80.740 164.160 81.820 164.460 ;
        RECT 81.130 163.620 81.430 164.160 ;
        RECT 80.900 163.580 81.820 163.620 ;
        RECT 80.740 163.280 81.820 163.580 ;
        RECT 78.580 162.840 79.660 163.140 ;
        RECT 78.970 161.380 79.270 162.840 ;
        RECT 80.740 162.400 81.820 162.700 ;
        RECT 81.130 161.820 81.430 162.400 ;
        RECT 84.100 161.820 84.400 165.040 ;
        RECT 84.860 164.460 85.780 164.500 ;
        RECT 84.700 164.160 85.780 164.460 ;
        RECT 85.090 163.620 85.390 164.160 ;
        RECT 84.860 163.580 85.780 163.620 ;
        RECT 84.700 163.280 85.780 163.580 ;
        RECT 84.700 162.400 85.780 162.700 ;
        RECT 85.090 161.820 85.390 162.400 ;
        RECT 86.260 161.820 86.560 168.120 ;
        RECT 86.940 168.080 87.860 168.120 ;
        RECT 86.860 166.360 87.940 166.660 ;
        RECT 87.250 164.900 87.550 166.360 ;
        RECT 86.860 164.600 87.940 164.900 ;
        RECT 87.250 163.140 87.550 164.600 ;
        RECT 86.860 162.840 87.940 163.140 ;
        RECT 80.740 161.520 86.560 161.820 ;
        RECT 87.250 161.380 87.550 162.840 ;
        RECT 78.580 161.080 80.260 161.380 ;
        RECT 86.860 161.080 87.940 161.380 ;
        RECT 79.960 160.060 80.260 161.080 ;
        RECT 80.900 160.940 81.820 160.980 ;
        RECT 84.860 160.940 85.780 160.980 ;
        RECT 80.740 160.640 81.820 160.940 ;
        RECT 84.700 160.640 85.780 160.940 ;
        RECT 79.960 159.760 85.780 160.060 ;
        RECT 78.580 159.620 79.500 159.660 ;
        RECT 87.020 159.620 87.940 159.660 ;
        RECT 77.980 159.320 79.660 159.620 ;
        RECT 86.860 159.320 87.940 159.620 ;
        RECT 77.980 154.340 78.280 159.320 ;
        RECT 78.970 157.860 79.270 159.320 ;
        RECT 80.740 158.880 81.820 159.180 ;
        RECT 84.700 158.880 85.780 159.180 ;
        RECT 81.130 158.300 81.430 158.880 ;
        RECT 85.090 158.300 85.390 158.880 ;
        RECT 80.740 158.000 81.820 158.300 ;
        RECT 84.700 158.000 85.780 158.300 ;
        RECT 78.580 157.560 79.660 157.860 ;
        RECT 86.260 157.560 87.940 157.860 ;
        RECT 78.970 156.100 79.270 157.560 ;
        RECT 80.740 157.120 81.820 157.420 ;
        RECT 84.700 157.120 85.780 157.420 ;
        RECT 81.130 156.540 81.430 157.120 ;
        RECT 85.090 156.540 85.390 157.120 ;
        RECT 80.740 156.240 81.820 156.540 ;
        RECT 84.700 156.240 85.780 156.540 ;
        RECT 78.580 155.800 79.660 156.100 ;
        RECT 80.900 155.660 81.820 155.700 ;
        RECT 84.860 155.660 85.780 155.700 ;
        RECT 80.740 155.360 81.820 155.660 ;
        RECT 84.700 155.360 85.780 155.660 ;
        RECT 84.860 154.780 85.780 154.820 ;
        RECT 80.740 154.480 85.780 154.780 ;
        RECT 77.980 154.040 79.660 154.340 ;
        RECT 77.980 142.020 78.280 154.040 ;
        RECT 78.970 152.580 79.270 154.040 ;
        RECT 80.740 153.600 81.820 153.900 ;
        RECT 84.700 153.600 85.780 153.900 ;
        RECT 81.130 153.020 81.430 153.600 ;
        RECT 85.090 153.020 85.390 153.600 ;
        RECT 80.740 152.720 81.820 153.020 ;
        RECT 84.700 152.720 85.780 153.020 ;
        RECT 86.260 152.580 86.560 157.560 ;
        RECT 86.860 156.100 87.780 156.140 ;
        RECT 86.860 155.800 88.540 156.100 ;
        RECT 87.020 154.340 87.940 154.380 ;
        RECT 86.860 154.040 87.940 154.340 ;
        RECT 78.580 152.280 79.660 152.580 ;
        RECT 86.260 152.280 87.940 152.580 ;
        RECT 78.970 150.820 79.270 152.280 ;
        RECT 80.740 151.840 81.820 152.140 ;
        RECT 84.700 151.840 85.780 152.140 ;
        RECT 81.130 151.260 81.430 151.840 ;
        RECT 85.090 151.260 85.390 151.840 ;
        RECT 80.740 150.960 81.820 151.260 ;
        RECT 84.700 150.960 85.780 151.260 ;
        RECT 78.580 150.520 79.660 150.820 ;
        RECT 80.900 150.380 81.820 150.420 ;
        RECT 84.860 150.380 85.780 150.420 ;
        RECT 80.740 150.080 81.820 150.380 ;
        RECT 84.700 150.080 85.780 150.380 ;
        RECT 86.260 149.500 86.560 152.280 ;
        RECT 86.860 150.820 87.780 150.860 ;
        RECT 86.860 150.520 87.940 150.820 ;
        RECT 80.740 149.200 86.560 149.500 ;
        RECT 78.580 148.760 79.660 149.060 ;
        RECT 86.860 148.760 87.940 149.060 ;
        RECT 80.900 148.620 81.820 148.660 ;
        RECT 84.860 148.620 85.780 148.660 ;
        RECT 80.740 148.320 81.820 148.620 ;
        RECT 84.700 148.320 85.780 148.620 ;
        RECT 86.260 148.460 87.160 148.760 ;
        RECT 80.900 147.740 81.820 147.780 ;
        RECT 86.260 147.740 86.560 148.460 ;
        RECT 80.740 147.440 81.820 147.740 ;
        RECT 82.120 147.440 86.560 147.740 ;
        RECT 78.580 147.000 80.440 147.300 ;
        RECT 78.580 145.240 79.660 145.540 ;
        RECT 78.580 143.480 79.660 143.780 ;
        RECT 77.980 141.720 79.660 142.020 ;
        RECT 80.140 141.580 80.440 147.000 ;
        RECT 80.740 146.560 81.820 146.860 ;
        RECT 81.130 145.980 81.430 146.560 ;
        RECT 80.740 145.680 81.820 145.980 ;
        RECT 80.740 144.800 81.820 145.100 ;
        RECT 81.130 144.220 81.430 144.800 ;
        RECT 80.740 143.920 81.820 144.220 ;
        RECT 80.900 143.340 81.820 143.380 ;
        RECT 82.120 143.340 82.420 147.440 ;
        RECT 86.860 147.000 87.940 147.300 ;
        RECT 84.860 146.860 85.780 146.900 ;
        RECT 84.700 146.560 85.780 146.860 ;
        RECT 84.860 145.980 85.780 146.020 ;
        RECT 84.700 145.680 85.780 145.980 ;
        RECT 86.860 145.540 87.780 145.580 ;
        RECT 86.860 145.240 87.940 145.540 ;
        RECT 80.740 143.040 82.420 143.340 ;
        RECT 84.100 144.800 85.780 145.100 ;
        RECT 84.100 144.220 84.400 144.800 ;
        RECT 84.100 143.920 85.780 144.220 ;
        RECT 80.900 142.460 81.820 142.500 ;
        RECT 80.740 142.160 81.820 142.460 ;
        RECT 84.100 142.460 84.400 143.920 ;
        RECT 88.240 143.780 88.540 155.800 ;
        RECT 86.860 143.480 88.540 143.780 ;
        RECT 84.860 143.340 85.780 143.380 ;
        RECT 84.700 143.040 85.780 143.340 ;
        RECT 84.100 142.160 85.780 142.460 ;
        RECT 87.020 142.020 87.940 142.060 ;
        RECT 86.860 141.720 87.940 142.020 ;
        RECT 80.140 141.280 85.780 141.580 ;
        RECT 80.900 140.700 81.820 140.740 ;
        RECT 84.860 140.700 85.780 140.740 ;
        RECT 80.140 140.400 81.820 140.700 ;
        RECT 84.700 140.400 86.560 140.700 ;
        RECT 80.140 140.260 80.440 140.400 ;
        RECT 73.480 139.960 80.440 140.260 ;
        RECT 68.140 139.820 69.060 139.860 ;
        RECT 72.100 139.820 73.020 139.860 ;
        RECT 73.480 139.820 73.780 139.960 ;
        RECT 67.360 139.520 69.220 139.820 ;
        RECT 72.100 139.520 73.780 139.820 ;
        RECT 76.420 139.010 77.500 139.960 ;
        RECT 80.140 139.820 80.440 139.960 ;
        RECT 86.260 140.260 86.560 140.400 ;
        RECT 89.020 140.260 90.100 210.360 ;
        RECT 92.560 210.220 92.860 210.360 ;
        RECT 98.680 210.660 98.980 210.800 ;
        RECT 101.620 210.660 102.700 211.610 ;
        RECT 106.100 211.100 107.020 211.140 ;
        RECT 110.060 211.100 110.980 211.140 ;
        RECT 105.340 210.800 107.020 211.100 ;
        RECT 109.900 210.800 111.760 211.100 ;
        RECT 105.340 210.660 105.640 210.800 ;
        RECT 98.680 210.360 105.640 210.660 ;
        RECT 93.340 210.220 94.260 210.260 ;
        RECT 97.300 210.220 98.220 210.260 ;
        RECT 98.680 210.220 98.980 210.360 ;
        RECT 92.560 209.920 94.420 210.220 ;
        RECT 97.300 209.920 98.980 210.220 ;
        RECT 97.300 209.340 98.220 209.570 ;
        RECT 93.340 209.040 98.380 209.340 ;
        RECT 91.180 208.600 92.860 208.900 ;
        RECT 99.460 208.600 100.540 208.900 ;
        RECT 91.180 207.140 92.100 207.180 ;
        RECT 91.180 206.840 92.260 207.140 ;
        RECT 92.560 206.700 92.860 208.600 ;
        RECT 93.340 208.460 94.260 208.500 ;
        RECT 97.300 208.460 98.220 208.500 ;
        RECT 93.340 208.160 94.420 208.460 ;
        RECT 97.300 208.160 98.380 208.460 ;
        RECT 93.340 207.580 94.260 207.620 ;
        RECT 93.340 207.280 94.420 207.580 ;
        RECT 94.720 207.280 98.380 207.580 ;
        RECT 94.720 206.700 95.020 207.280 ;
        RECT 99.460 206.840 100.540 207.140 ;
        RECT 92.560 206.400 95.020 206.700 ;
        RECT 97.300 206.400 98.380 206.700 ;
        RECT 94.720 205.820 95.020 206.400 ;
        RECT 97.690 205.820 97.990 206.400 ;
        RECT 93.340 205.520 95.020 205.820 ;
        RECT 97.300 205.520 98.380 205.820 ;
        RECT 91.180 205.080 92.260 205.380 ;
        RECT 99.460 205.080 100.540 205.380 ;
        RECT 91.960 204.780 92.860 205.080 ;
        RECT 92.560 204.060 92.860 204.780 ;
        RECT 93.340 204.940 94.260 204.980 ;
        RECT 97.300 204.940 98.220 204.980 ;
        RECT 93.340 204.640 94.420 204.940 ;
        RECT 97.300 204.640 98.380 204.940 ;
        RECT 92.560 203.760 98.380 204.060 ;
        RECT 91.180 203.320 92.260 203.620 ;
        RECT 99.460 203.320 100.540 203.620 ;
        RECT 91.960 203.020 92.860 203.320 ;
        RECT 92.560 202.300 92.860 203.020 ;
        RECT 93.340 203.180 94.260 203.220 ;
        RECT 97.300 203.180 98.220 203.220 ;
        RECT 93.340 202.880 94.420 203.180 ;
        RECT 97.300 202.880 98.380 203.180 ;
        RECT 97.300 202.300 98.220 202.340 ;
        RECT 92.560 202.000 95.020 202.300 ;
        RECT 97.300 202.000 98.380 202.300 ;
        RECT 91.180 201.860 92.100 201.900 ;
        RECT 91.180 201.560 92.260 201.860 ;
        RECT 94.720 201.420 95.020 202.000 ;
        RECT 99.460 201.560 100.540 201.860 ;
        RECT 93.340 201.120 94.420 201.420 ;
        RECT 94.720 201.120 98.380 201.420 ;
        RECT 93.730 200.540 94.030 201.120 ;
        RECT 94.720 200.540 95.020 201.120 ;
        RECT 93.340 200.240 94.420 200.540 ;
        RECT 94.720 200.240 98.380 200.540 ;
        RECT 91.180 199.800 92.260 200.100 ;
        RECT 99.460 199.800 100.540 200.100 ;
        RECT 91.570 198.340 91.870 199.800 ;
        RECT 93.340 199.660 94.260 199.700 ;
        RECT 97.300 199.660 98.220 199.700 ;
        RECT 93.340 199.360 94.420 199.660 ;
        RECT 97.300 199.360 98.380 199.660 ;
        RECT 93.340 198.480 98.380 198.780 ;
        RECT 91.180 198.040 92.860 198.340 ;
        RECT 99.460 198.040 100.540 198.340 ;
        RECT 92.560 197.020 92.860 198.040 ;
        RECT 93.340 197.900 94.260 197.940 ;
        RECT 97.300 197.900 98.220 197.940 ;
        RECT 93.340 197.600 94.420 197.900 ;
        RECT 97.300 197.600 98.380 197.900 ;
        RECT 92.560 196.720 98.380 197.020 ;
        RECT 99.460 196.580 100.380 196.620 ;
        RECT 91.180 196.280 92.260 196.580 ;
        RECT 99.460 196.280 100.540 196.580 ;
        RECT 93.340 196.140 94.260 196.180 ;
        RECT 97.300 196.140 98.220 196.180 ;
        RECT 93.340 195.840 94.420 196.140 ;
        RECT 97.300 195.840 98.380 196.140 ;
        RECT 93.340 195.260 94.260 195.300 ;
        RECT 93.340 194.960 98.380 195.260 ;
        RECT 91.180 194.520 92.260 194.820 ;
        RECT 91.570 193.060 91.870 194.520 ;
        RECT 93.340 194.080 94.420 194.380 ;
        RECT 93.730 193.500 94.030 194.080 ;
        RECT 93.340 193.200 94.420 193.500 ;
        RECT 91.180 192.760 92.260 193.060 ;
        RECT 91.570 191.340 91.870 192.760 ;
        RECT 93.340 192.620 94.260 192.660 ;
        RECT 93.340 192.320 94.420 192.620 ;
        RECT 93.730 191.780 94.030 192.320 ;
        RECT 93.340 191.740 94.260 191.780 ;
        RECT 93.340 191.440 94.420 191.740 ;
        RECT 91.180 191.300 92.100 191.340 ;
        RECT 91.180 191.000 92.260 191.300 ;
        RECT 91.570 189.540 91.870 191.000 ;
        RECT 93.340 190.560 94.420 190.860 ;
        RECT 93.730 189.980 94.030 190.560 ;
        RECT 93.340 189.680 94.420 189.980 ;
        RECT 91.180 189.240 92.260 189.540 ;
        RECT 93.340 189.100 94.260 189.140 ;
        RECT 94.720 189.100 95.020 194.960 ;
        RECT 99.460 194.520 100.540 194.820 ;
        RECT 97.300 194.080 98.380 194.380 ;
        RECT 97.690 193.500 97.990 194.080 ;
        RECT 97.300 193.200 98.380 193.500 ;
        RECT 99.850 193.100 100.150 194.520 ;
        RECT 99.460 193.060 100.380 193.100 ;
        RECT 99.460 192.760 100.540 193.060 ;
        RECT 97.300 192.620 98.220 192.660 ;
        RECT 97.300 192.320 98.380 192.620 ;
        RECT 97.690 191.780 97.990 192.320 ;
        RECT 97.300 191.740 98.220 191.780 ;
        RECT 97.300 191.440 98.380 191.740 ;
        RECT 99.460 191.000 100.540 191.300 ;
        RECT 97.300 190.560 98.380 190.860 ;
        RECT 97.690 189.980 97.990 190.560 ;
        RECT 97.300 189.680 98.380 189.980 ;
        RECT 99.850 189.540 100.150 191.000 ;
        RECT 98.680 189.240 100.540 189.540 ;
        RECT 93.340 188.800 94.420 189.100 ;
        RECT 94.720 188.800 98.380 189.100 ;
        RECT 93.340 188.220 94.260 188.260 ;
        RECT 97.300 188.220 98.220 188.260 ;
        RECT 93.340 187.920 94.420 188.220 ;
        RECT 97.300 187.920 98.380 188.220 ;
        RECT 91.180 187.480 92.260 187.780 ;
        RECT 91.570 186.020 91.870 187.480 ;
        RECT 93.340 187.040 94.420 187.340 ;
        RECT 97.300 187.040 98.380 187.340 ;
        RECT 93.730 186.460 94.030 187.040 ;
        RECT 97.690 186.460 97.990 187.040 ;
        RECT 93.340 186.160 98.380 186.460 ;
        RECT 91.180 185.720 92.260 186.020 ;
        RECT 91.570 184.260 91.870 185.720 ;
        RECT 93.340 185.580 94.260 185.620 ;
        RECT 93.340 185.280 94.420 185.580 ;
        RECT 93.730 184.740 94.030 185.280 ;
        RECT 93.340 184.700 94.260 184.740 ;
        RECT 93.340 184.400 94.420 184.700 ;
        RECT 91.180 183.960 92.260 184.260 ;
        RECT 91.570 182.500 91.870 183.960 ;
        RECT 93.340 183.520 94.420 183.820 ;
        RECT 93.730 182.940 94.030 183.520 ;
        RECT 94.720 182.940 95.020 186.160 ;
        RECT 97.300 185.280 98.380 185.580 ;
        RECT 97.690 184.740 97.990 185.280 ;
        RECT 97.300 184.700 98.220 184.740 ;
        RECT 97.300 184.400 98.380 184.700 ;
        RECT 97.300 183.520 98.380 183.820 ;
        RECT 96.510 182.940 96.850 183.210 ;
        RECT 97.690 182.940 97.990 183.520 ;
        RECT 98.680 182.940 98.980 189.240 ;
        RECT 99.460 187.480 100.540 187.780 ;
        RECT 99.850 186.020 100.150 187.480 ;
        RECT 99.460 185.720 100.540 186.020 ;
        RECT 99.850 184.260 100.150 185.720 ;
        RECT 99.460 183.960 100.540 184.260 ;
        RECT 93.340 182.640 98.980 182.940 ;
        RECT 91.180 182.200 92.860 182.500 ;
        RECT 96.510 182.290 96.850 182.640 ;
        RECT 99.850 182.500 100.150 183.960 ;
        RECT 99.460 182.200 100.540 182.500 ;
        RECT 91.180 180.440 92.260 180.740 ;
        RECT 91.570 178.980 91.870 180.440 ;
        RECT 91.180 178.680 92.260 178.980 ;
        RECT 91.570 177.220 91.870 178.680 ;
        RECT 91.180 176.920 92.260 177.220 ;
        RECT 91.570 175.500 91.870 176.920 ;
        RECT 92.560 175.900 92.860 182.200 ;
        RECT 93.340 182.060 94.260 182.100 ;
        RECT 97.300 182.060 98.220 182.100 ;
        RECT 93.340 181.760 94.420 182.060 ;
        RECT 97.300 181.760 98.380 182.060 ;
        RECT 93.340 181.180 94.260 181.220 ;
        RECT 97.300 181.180 98.220 181.220 ;
        RECT 93.340 180.880 94.420 181.180 ;
        RECT 97.300 180.880 98.380 181.180 ;
        RECT 99.460 180.440 100.540 180.740 ;
        RECT 93.340 180.000 94.420 180.300 ;
        RECT 97.300 180.000 98.380 180.300 ;
        RECT 93.730 179.420 94.030 180.000 ;
        RECT 97.690 179.420 97.990 180.000 ;
        RECT 93.340 179.120 98.380 179.420 ;
        RECT 93.340 178.540 94.260 178.580 ;
        RECT 93.340 178.240 94.420 178.540 ;
        RECT 93.730 177.700 94.030 178.240 ;
        RECT 93.340 177.660 94.260 177.700 ;
        RECT 93.340 177.360 94.420 177.660 ;
        RECT 93.340 176.480 94.420 176.780 ;
        RECT 93.730 175.900 94.030 176.480 ;
        RECT 94.720 175.900 95.020 179.120 ;
        RECT 99.850 178.980 100.150 180.440 ;
        RECT 99.460 178.680 100.540 178.980 ;
        RECT 97.300 178.240 98.380 178.540 ;
        RECT 97.690 177.700 97.990 178.240 ;
        RECT 97.300 177.660 98.220 177.700 ;
        RECT 97.300 177.360 98.380 177.660 ;
        RECT 99.850 177.220 100.150 178.680 ;
        RECT 99.460 176.920 100.540 177.220 ;
        RECT 97.300 176.480 98.380 176.780 ;
        RECT 95.635 175.900 95.975 176.170 ;
        RECT 97.690 175.900 97.990 176.480 ;
        RECT 92.560 175.600 98.380 175.900 ;
        RECT 91.180 175.460 92.100 175.500 ;
        RECT 91.180 175.160 92.260 175.460 ;
        RECT 95.635 175.250 95.975 175.600 ;
        RECT 99.850 175.460 100.150 176.920 ;
        RECT 99.460 175.160 100.540 175.460 ;
        RECT 93.340 175.020 94.260 175.060 ;
        RECT 97.300 175.020 98.220 175.060 ;
        RECT 93.340 174.720 94.420 175.020 ;
        RECT 97.300 174.720 98.380 175.020 ;
        RECT 93.340 174.140 94.260 174.180 ;
        RECT 97.300 174.140 98.220 174.180 ;
        RECT 93.340 173.840 94.420 174.140 ;
        RECT 97.300 173.840 98.380 174.140 ;
        RECT 91.180 173.400 92.260 173.700 ;
        RECT 99.460 173.400 100.540 173.700 ;
        RECT 91.570 171.940 91.870 173.400 ;
        RECT 93.340 172.960 94.420 173.260 ;
        RECT 97.300 172.960 98.380 173.260 ;
        RECT 93.730 172.380 94.030 172.960 ;
        RECT 97.690 172.380 97.990 172.960 ;
        RECT 93.340 172.080 98.380 172.380 ;
        RECT 91.180 171.640 92.260 171.940 ;
        RECT 91.570 170.180 91.870 171.640 ;
        RECT 93.340 171.500 94.260 171.540 ;
        RECT 93.340 171.200 94.420 171.500 ;
        RECT 93.730 170.660 94.030 171.200 ;
        RECT 93.340 170.620 94.260 170.660 ;
        RECT 93.340 170.320 94.420 170.620 ;
        RECT 91.180 169.880 92.260 170.180 ;
        RECT 91.570 168.420 91.870 169.880 ;
        RECT 93.340 169.440 94.420 169.740 ;
        RECT 93.730 168.860 94.030 169.440 ;
        RECT 94.720 169.130 95.020 172.080 ;
        RECT 99.850 171.940 100.150 173.400 ;
        RECT 99.460 171.640 100.540 171.940 ;
        RECT 97.300 171.200 98.380 171.500 ;
        RECT 97.690 170.660 97.990 171.200 ;
        RECT 97.300 170.620 98.220 170.660 ;
        RECT 97.300 170.320 98.380 170.620 ;
        RECT 99.850 170.180 100.150 171.640 ;
        RECT 99.460 169.880 100.540 170.180 ;
        RECT 97.300 169.440 98.380 169.740 ;
        RECT 94.720 168.860 95.175 169.130 ;
        RECT 97.690 168.900 97.990 169.440 ;
        RECT 97.300 168.860 98.220 168.900 ;
        RECT 93.340 168.560 98.380 168.860 ;
        RECT 91.180 168.120 92.860 168.420 ;
        RECT 94.835 168.210 95.175 168.560 ;
        RECT 99.850 168.420 100.150 169.880 ;
        RECT 99.460 168.120 100.540 168.420 ;
        RECT 91.260 168.080 92.180 168.120 ;
        RECT 91.180 166.360 92.260 166.660 ;
        RECT 91.570 164.900 91.870 166.360 ;
        RECT 91.180 164.600 92.260 164.900 ;
        RECT 91.570 163.140 91.870 164.600 ;
        RECT 91.180 162.840 92.260 163.140 ;
        RECT 91.570 161.380 91.870 162.840 ;
        RECT 92.560 161.820 92.860 168.120 ;
        RECT 93.340 167.980 94.260 168.020 ;
        RECT 97.300 167.980 98.220 168.020 ;
        RECT 93.340 167.680 94.420 167.980 ;
        RECT 97.300 167.680 98.380 167.980 ;
        RECT 93.340 167.100 94.260 167.140 ;
        RECT 97.300 167.100 98.220 167.140 ;
        RECT 93.340 166.800 94.420 167.100 ;
        RECT 97.300 166.800 98.380 167.100 ;
        RECT 99.460 166.360 100.540 166.660 ;
        RECT 93.340 165.920 94.420 166.220 ;
        RECT 97.300 165.920 98.380 166.220 ;
        RECT 93.730 165.340 94.030 165.920 ;
        RECT 97.690 165.340 97.990 165.920 ;
        RECT 93.340 165.040 98.380 165.340 ;
        RECT 93.340 164.460 94.260 164.500 ;
        RECT 93.340 164.160 94.420 164.460 ;
        RECT 93.730 163.620 94.030 164.160 ;
        RECT 93.340 163.580 94.260 163.620 ;
        RECT 93.340 163.280 94.420 163.580 ;
        RECT 93.340 162.400 94.420 162.700 ;
        RECT 93.730 161.820 94.030 162.400 ;
        RECT 94.720 161.820 95.020 165.040 ;
        RECT 99.850 164.900 100.150 166.360 ;
        RECT 99.460 164.600 100.540 164.900 ;
        RECT 97.300 164.160 98.380 164.460 ;
        RECT 97.690 163.620 97.990 164.160 ;
        RECT 97.300 163.580 98.220 163.620 ;
        RECT 97.300 163.280 98.380 163.580 ;
        RECT 99.850 163.140 100.150 164.600 ;
        RECT 99.460 162.840 100.540 163.140 ;
        RECT 97.300 162.400 98.380 162.700 ;
        RECT 97.690 161.820 97.990 162.400 ;
        RECT 92.560 161.520 98.380 161.820 ;
        RECT 99.850 161.380 100.150 162.840 ;
        RECT 91.180 161.080 92.260 161.380 ;
        RECT 98.860 161.080 100.540 161.380 ;
        RECT 93.340 160.940 94.260 160.980 ;
        RECT 97.300 160.940 98.220 160.980 ;
        RECT 93.340 160.640 94.420 160.940 ;
        RECT 97.300 160.640 98.380 160.940 ;
        RECT 98.860 160.060 99.160 161.080 ;
        RECT 93.340 159.760 99.160 160.060 ;
        RECT 91.180 159.620 92.100 159.660 ;
        RECT 99.460 159.620 100.380 159.660 ;
        RECT 91.180 159.320 92.260 159.620 ;
        RECT 99.460 159.320 101.140 159.620 ;
        RECT 93.340 158.880 94.420 159.180 ;
        RECT 97.300 158.880 98.380 159.180 ;
        RECT 93.730 158.300 94.030 158.880 ;
        RECT 97.690 158.300 97.990 158.880 ;
        RECT 93.340 158.000 94.420 158.300 ;
        RECT 97.300 158.000 98.380 158.300 ;
        RECT 99.850 157.860 100.150 159.320 ;
        RECT 91.180 157.560 92.860 157.860 ;
        RECT 99.460 157.560 100.540 157.860 ;
        RECT 91.180 156.100 92.100 156.140 ;
        RECT 90.580 155.800 92.260 156.100 ;
        RECT 90.580 143.780 90.880 155.800 ;
        RECT 91.180 154.340 92.100 154.380 ;
        RECT 91.180 154.040 92.260 154.340 ;
        RECT 92.560 152.580 92.860 157.560 ;
        RECT 93.340 157.120 94.420 157.420 ;
        RECT 97.300 157.120 98.380 157.420 ;
        RECT 93.730 156.540 94.030 157.120 ;
        RECT 97.690 156.540 97.990 157.120 ;
        RECT 93.340 156.240 94.420 156.540 ;
        RECT 97.300 156.240 98.380 156.540 ;
        RECT 99.850 156.100 100.150 157.560 ;
        RECT 99.460 155.800 100.540 156.100 ;
        RECT 93.340 155.660 94.260 155.700 ;
        RECT 97.300 155.660 98.220 155.700 ;
        RECT 93.340 155.360 94.420 155.660 ;
        RECT 97.300 155.360 98.380 155.660 ;
        RECT 93.340 154.780 94.260 154.820 ;
        RECT 93.340 154.480 98.380 154.780 ;
        RECT 100.840 154.340 101.140 159.320 ;
        RECT 99.460 154.040 101.140 154.340 ;
        RECT 93.340 153.600 94.420 153.900 ;
        RECT 97.300 153.600 98.380 153.900 ;
        RECT 93.730 153.020 94.030 153.600 ;
        RECT 97.690 153.020 97.990 153.600 ;
        RECT 93.340 152.720 94.420 153.020 ;
        RECT 97.300 152.720 98.380 153.020 ;
        RECT 99.850 152.580 100.150 154.040 ;
        RECT 91.180 152.280 92.860 152.580 ;
        RECT 99.460 152.280 100.540 152.580 ;
        RECT 91.340 150.820 92.260 150.860 ;
        RECT 91.180 150.520 92.260 150.820 ;
        RECT 92.560 149.500 92.860 152.280 ;
        RECT 93.340 151.840 94.420 152.140 ;
        RECT 97.300 151.840 98.380 152.140 ;
        RECT 93.730 151.260 94.030 151.840 ;
        RECT 97.690 151.260 97.990 151.840 ;
        RECT 93.340 150.960 94.420 151.260 ;
        RECT 97.300 150.960 98.380 151.260 ;
        RECT 99.850 150.820 100.150 152.280 ;
        RECT 99.460 150.520 100.540 150.820 ;
        RECT 93.340 150.380 94.260 150.420 ;
        RECT 97.300 150.380 98.220 150.420 ;
        RECT 93.340 150.080 94.420 150.380 ;
        RECT 97.300 150.080 98.380 150.380 ;
        RECT 92.560 149.200 98.380 149.500 ;
        RECT 91.180 148.760 92.260 149.060 ;
        RECT 99.460 148.760 100.540 149.060 ;
        RECT 91.960 148.460 92.860 148.760 ;
        RECT 92.560 147.740 92.860 148.460 ;
        RECT 93.340 148.620 94.260 148.660 ;
        RECT 97.300 148.620 98.220 148.660 ;
        RECT 93.340 148.320 94.420 148.620 ;
        RECT 97.300 148.320 98.380 148.620 ;
        RECT 97.300 147.740 98.220 147.780 ;
        RECT 92.560 147.440 97.000 147.740 ;
        RECT 97.300 147.440 98.380 147.740 ;
        RECT 91.180 147.000 92.260 147.300 ;
        RECT 93.340 146.860 94.260 146.900 ;
        RECT 93.340 146.560 94.420 146.860 ;
        RECT 93.340 145.980 94.260 146.020 ;
        RECT 93.340 145.680 94.420 145.980 ;
        RECT 91.340 145.540 92.260 145.580 ;
        RECT 91.180 145.240 92.260 145.540 ;
        RECT 93.340 144.800 95.020 145.100 ;
        RECT 94.720 144.220 95.020 144.800 ;
        RECT 93.340 143.920 95.020 144.220 ;
        RECT 90.580 143.480 92.260 143.780 ;
        RECT 93.340 143.340 94.260 143.380 ;
        RECT 93.340 143.040 94.420 143.340 ;
        RECT 94.720 142.460 95.020 143.920 ;
        RECT 96.700 143.340 97.000 147.440 ;
        RECT 98.680 147.000 100.540 147.300 ;
        RECT 97.300 146.560 98.380 146.860 ;
        RECT 97.690 145.980 97.990 146.560 ;
        RECT 97.300 145.680 98.380 145.980 ;
        RECT 97.300 144.800 98.380 145.100 ;
        RECT 97.690 144.220 97.990 144.800 ;
        RECT 97.300 143.920 98.380 144.220 ;
        RECT 97.300 143.340 98.220 143.380 ;
        RECT 96.700 143.040 98.380 143.340 ;
        RECT 93.340 142.160 95.020 142.460 ;
        RECT 97.300 142.460 98.220 142.500 ;
        RECT 97.300 142.160 98.380 142.460 ;
        RECT 91.180 142.020 92.100 142.060 ;
        RECT 91.180 141.720 92.260 142.020 ;
        RECT 98.680 141.580 98.980 147.000 ;
        RECT 99.460 145.240 100.540 145.540 ;
        RECT 99.460 143.480 100.540 143.780 ;
        RECT 100.840 142.020 101.140 154.040 ;
        RECT 99.460 141.720 101.140 142.020 ;
        RECT 93.340 141.280 98.980 141.580 ;
        RECT 93.340 140.700 94.260 140.740 ;
        RECT 97.300 140.700 98.220 140.740 ;
        RECT 92.560 140.400 94.420 140.700 ;
        RECT 97.300 140.400 98.980 140.700 ;
        RECT 92.560 140.260 92.860 140.400 ;
        RECT 86.260 139.960 92.860 140.260 ;
        RECT 80.900 139.820 81.820 139.860 ;
        RECT 84.860 139.820 85.780 139.860 ;
        RECT 86.260 139.820 86.560 139.960 ;
        RECT 80.140 139.520 81.820 139.820 ;
        RECT 84.700 139.520 86.560 139.820 ;
        RECT 89.020 139.010 90.100 139.960 ;
        RECT 92.560 139.820 92.860 139.960 ;
        RECT 98.680 140.260 98.980 140.400 ;
        RECT 101.620 140.260 102.700 210.360 ;
        RECT 105.340 210.220 105.640 210.360 ;
        RECT 111.460 210.660 111.760 210.800 ;
        RECT 114.220 210.660 115.300 211.610 ;
        RECT 111.460 210.360 115.300 210.660 ;
        RECT 106.100 210.220 107.020 210.260 ;
        RECT 110.060 210.220 110.980 210.260 ;
        RECT 111.460 210.220 111.760 210.360 ;
        RECT 105.340 209.920 107.020 210.220 ;
        RECT 109.900 209.920 111.760 210.220 ;
        RECT 105.940 209.340 106.860 209.380 ;
        RECT 105.940 209.040 110.980 209.340 ;
        RECT 114.220 208.900 115.300 210.360 ;
        RECT 118.540 209.340 119.460 209.380 ;
        RECT 122.500 209.340 123.420 209.380 ;
        RECT 117.760 209.040 119.620 209.340 ;
        RECT 122.500 209.040 124.180 209.340 ;
        RECT 117.760 208.900 118.060 209.040 ;
        RECT 103.780 208.600 104.860 208.900 ;
        RECT 111.460 208.600 113.140 208.900 ;
        RECT 114.220 208.600 118.060 208.900 ;
        RECT 106.100 208.460 107.020 208.500 ;
        RECT 110.060 208.460 110.980 208.500 ;
        RECT 105.940 208.160 107.020 208.460 ;
        RECT 109.900 208.160 110.980 208.460 ;
        RECT 110.060 207.580 110.980 207.620 ;
        RECT 105.940 207.280 109.600 207.580 ;
        RECT 109.900 207.280 110.980 207.580 ;
        RECT 103.780 206.840 104.860 207.140 ;
        RECT 109.300 206.700 109.600 207.280 ;
        RECT 111.460 206.700 111.760 208.600 ;
        RECT 112.060 207.140 112.980 207.180 ;
        RECT 112.060 206.840 113.140 207.140 ;
        RECT 105.940 206.400 107.020 206.700 ;
        RECT 109.300 206.400 111.760 206.700 ;
        RECT 106.330 205.820 106.630 206.400 ;
        RECT 109.300 205.820 109.600 206.400 ;
        RECT 105.940 205.520 107.020 205.820 ;
        RECT 109.300 205.520 110.980 205.820 ;
        RECT 103.780 205.080 104.860 205.380 ;
        RECT 112.060 205.080 113.140 205.380 ;
        RECT 106.100 204.940 107.020 204.980 ;
        RECT 110.060 204.940 110.980 204.980 ;
        RECT 105.940 204.640 107.020 204.940 ;
        RECT 109.900 204.640 110.980 204.940 ;
        RECT 111.460 204.780 112.360 205.080 ;
        RECT 111.460 204.060 111.760 204.780 ;
        RECT 105.940 203.760 111.760 204.060 ;
        RECT 103.780 203.320 104.860 203.620 ;
        RECT 112.060 203.320 113.140 203.620 ;
        RECT 106.100 203.180 107.020 203.220 ;
        RECT 110.060 203.180 110.980 203.220 ;
        RECT 105.940 202.880 107.020 203.180 ;
        RECT 109.900 202.880 110.980 203.180 ;
        RECT 111.460 203.020 112.360 203.320 ;
        RECT 106.100 202.300 107.020 202.340 ;
        RECT 111.460 202.300 111.760 203.020 ;
        RECT 105.940 202.000 107.020 202.300 ;
        RECT 109.300 202.000 111.760 202.300 ;
        RECT 103.780 201.560 104.860 201.860 ;
        RECT 109.300 201.420 109.600 202.000 ;
        RECT 112.220 201.860 113.140 201.900 ;
        RECT 112.060 201.560 113.140 201.860 ;
        RECT 105.940 201.120 109.600 201.420 ;
        RECT 109.900 201.120 110.980 201.420 ;
        RECT 109.300 200.540 109.600 201.120 ;
        RECT 110.290 200.540 110.590 201.120 ;
        RECT 105.940 200.240 109.600 200.540 ;
        RECT 109.900 200.240 110.980 200.540 ;
        RECT 103.780 199.800 104.860 200.100 ;
        RECT 112.060 199.800 113.140 200.100 ;
        RECT 106.100 199.660 107.020 199.700 ;
        RECT 110.060 199.660 110.980 199.700 ;
        RECT 105.940 199.360 107.020 199.660 ;
        RECT 109.900 199.360 110.980 199.660 ;
        RECT 109.980 198.780 110.900 198.820 ;
        RECT 105.940 198.480 110.980 198.780 ;
        RECT 112.450 198.340 112.750 199.800 ;
        RECT 103.780 198.040 104.860 198.340 ;
        RECT 111.460 198.040 113.140 198.340 ;
        RECT 106.100 197.900 107.020 197.940 ;
        RECT 110.060 197.900 110.980 197.940 ;
        RECT 105.940 197.600 107.020 197.900 ;
        RECT 109.900 197.600 110.980 197.900 ;
        RECT 111.460 197.020 111.760 198.040 ;
        RECT 105.940 196.720 111.760 197.020 ;
        RECT 103.940 196.580 104.860 196.620 ;
        RECT 103.780 196.280 104.860 196.580 ;
        RECT 112.060 196.280 113.140 196.580 ;
        RECT 106.100 196.140 107.020 196.180 ;
        RECT 110.060 196.140 110.980 196.180 ;
        RECT 105.940 195.840 107.020 196.140 ;
        RECT 109.900 195.840 110.980 196.140 ;
        RECT 110.060 195.260 110.980 195.300 ;
        RECT 105.940 194.960 110.980 195.260 ;
        RECT 103.780 194.520 104.860 194.820 ;
        RECT 104.170 193.100 104.470 194.520 ;
        RECT 105.940 194.080 107.020 194.380 ;
        RECT 106.330 193.500 106.630 194.080 ;
        RECT 105.940 193.200 107.020 193.500 ;
        RECT 103.940 193.060 104.860 193.100 ;
        RECT 103.780 192.760 104.860 193.060 ;
        RECT 106.100 192.620 107.020 192.660 ;
        RECT 105.940 192.320 107.020 192.620 ;
        RECT 106.330 191.780 106.630 192.320 ;
        RECT 106.100 191.740 107.020 191.780 ;
        RECT 105.940 191.440 107.020 191.740 ;
        RECT 103.780 191.000 104.860 191.300 ;
        RECT 104.170 189.540 104.470 191.000 ;
        RECT 105.940 190.560 107.020 190.860 ;
        RECT 106.330 189.980 106.630 190.560 ;
        RECT 105.940 189.680 107.020 189.980 ;
        RECT 103.780 189.240 105.640 189.540 ;
        RECT 103.780 187.480 104.860 187.780 ;
        RECT 104.170 186.020 104.470 187.480 ;
        RECT 103.780 185.720 104.860 186.020 ;
        RECT 104.170 184.260 104.470 185.720 ;
        RECT 103.780 183.960 104.860 184.260 ;
        RECT 104.170 182.500 104.470 183.960 ;
        RECT 105.340 182.940 105.640 189.240 ;
        RECT 109.300 189.100 109.600 194.960 ;
        RECT 112.060 194.820 112.980 194.860 ;
        RECT 112.060 194.520 113.140 194.820 ;
        RECT 109.900 194.080 110.980 194.380 ;
        RECT 110.290 193.500 110.590 194.080 ;
        RECT 109.900 193.200 110.980 193.500 ;
        RECT 112.450 193.060 112.750 194.520 ;
        RECT 112.060 192.760 113.140 193.060 ;
        RECT 110.060 192.620 110.980 192.660 ;
        RECT 109.900 192.320 110.980 192.620 ;
        RECT 110.290 191.780 110.590 192.320 ;
        RECT 110.060 191.740 110.980 191.780 ;
        RECT 109.900 191.440 110.980 191.740 ;
        RECT 112.450 191.340 112.750 192.760 ;
        RECT 112.060 191.300 112.980 191.340 ;
        RECT 112.060 191.000 113.140 191.300 ;
        RECT 109.900 190.560 110.980 190.860 ;
        RECT 110.290 189.980 110.590 190.560 ;
        RECT 109.900 189.680 110.980 189.980 ;
        RECT 112.450 189.540 112.750 191.000 ;
        RECT 112.060 189.240 113.140 189.540 ;
        RECT 110.060 189.100 110.980 189.140 ;
        RECT 105.940 188.800 109.600 189.100 ;
        RECT 109.900 188.800 110.980 189.100 ;
        RECT 106.100 188.220 107.020 188.260 ;
        RECT 110.060 188.220 110.980 188.260 ;
        RECT 105.940 187.920 107.020 188.220 ;
        RECT 109.900 187.920 110.980 188.220 ;
        RECT 112.060 187.480 113.140 187.780 ;
        RECT 105.940 187.040 107.020 187.340 ;
        RECT 109.900 187.040 110.980 187.340 ;
        RECT 106.330 186.460 106.630 187.040 ;
        RECT 110.290 186.460 110.590 187.040 ;
        RECT 105.940 186.160 110.980 186.460 ;
        RECT 105.940 185.280 107.020 185.580 ;
        RECT 106.330 184.740 106.630 185.280 ;
        RECT 106.100 184.700 107.020 184.740 ;
        RECT 105.940 184.400 107.020 184.700 ;
        RECT 105.940 183.520 107.020 183.820 ;
        RECT 106.330 182.940 106.630 183.520 ;
        RECT 107.470 182.940 107.810 183.210 ;
        RECT 109.300 182.940 109.600 186.160 ;
        RECT 112.450 186.020 112.750 187.480 ;
        RECT 112.060 185.720 113.140 186.020 ;
        RECT 110.060 185.580 110.980 185.620 ;
        RECT 109.900 185.280 110.980 185.580 ;
        RECT 110.290 184.740 110.590 185.280 ;
        RECT 110.060 184.700 110.980 184.740 ;
        RECT 109.900 184.400 110.980 184.700 ;
        RECT 112.450 184.260 112.750 185.720 ;
        RECT 112.060 183.960 113.140 184.260 ;
        RECT 109.900 183.520 110.980 183.820 ;
        RECT 110.290 182.940 110.590 183.520 ;
        RECT 105.340 182.640 110.980 182.940 ;
        RECT 103.780 182.200 104.860 182.500 ;
        RECT 107.470 182.290 107.810 182.640 ;
        RECT 112.450 182.500 112.750 183.960 ;
        RECT 111.460 182.200 113.140 182.500 ;
        RECT 106.100 182.060 107.020 182.100 ;
        RECT 110.060 182.060 110.980 182.100 ;
        RECT 105.940 181.760 107.020 182.060 ;
        RECT 109.900 181.760 110.980 182.060 ;
        RECT 106.100 181.180 107.020 181.220 ;
        RECT 110.060 181.180 110.980 181.220 ;
        RECT 105.940 180.880 107.020 181.180 ;
        RECT 109.900 180.880 110.980 181.180 ;
        RECT 103.780 180.440 104.860 180.740 ;
        RECT 104.170 178.980 104.470 180.440 ;
        RECT 105.940 180.000 107.020 180.300 ;
        RECT 109.900 180.000 110.980 180.300 ;
        RECT 106.330 179.420 106.630 180.000 ;
        RECT 110.290 179.420 110.590 180.000 ;
        RECT 105.940 179.120 110.980 179.420 ;
        RECT 103.780 178.680 104.860 178.980 ;
        RECT 104.170 177.220 104.470 178.680 ;
        RECT 105.940 178.240 107.020 178.540 ;
        RECT 106.330 177.700 106.630 178.240 ;
        RECT 106.100 177.660 107.020 177.700 ;
        RECT 105.940 177.360 107.020 177.660 ;
        RECT 103.780 176.920 104.860 177.220 ;
        RECT 104.170 175.460 104.470 176.920 ;
        RECT 105.940 176.480 107.020 176.780 ;
        RECT 106.330 175.900 106.630 176.480 ;
        RECT 108.345 175.900 108.685 176.170 ;
        RECT 109.300 175.900 109.600 179.120 ;
        RECT 110.060 178.540 110.980 178.580 ;
        RECT 109.900 178.240 110.980 178.540 ;
        RECT 110.290 177.700 110.590 178.240 ;
        RECT 110.060 177.660 110.980 177.700 ;
        RECT 109.900 177.360 110.980 177.660 ;
        RECT 109.900 176.480 110.980 176.780 ;
        RECT 110.290 175.900 110.590 176.480 ;
        RECT 111.460 175.900 111.760 182.200 ;
        RECT 112.060 180.440 113.140 180.740 ;
        RECT 112.450 178.980 112.750 180.440 ;
        RECT 112.060 178.680 113.140 178.980 ;
        RECT 112.450 177.220 112.750 178.680 ;
        RECT 112.060 176.920 113.140 177.220 ;
        RECT 105.940 175.600 111.760 175.900 ;
        RECT 103.780 175.160 104.860 175.460 ;
        RECT 108.345 175.250 108.685 175.600 ;
        RECT 112.450 175.500 112.750 176.920 ;
        RECT 112.220 175.460 113.140 175.500 ;
        RECT 112.060 175.160 113.140 175.460 ;
        RECT 106.100 175.020 107.020 175.060 ;
        RECT 110.060 175.020 110.980 175.060 ;
        RECT 105.940 174.720 107.020 175.020 ;
        RECT 109.900 174.720 110.980 175.020 ;
        RECT 106.100 174.140 107.020 174.180 ;
        RECT 110.060 174.140 110.980 174.180 ;
        RECT 105.940 173.840 107.020 174.140 ;
        RECT 109.900 173.840 110.980 174.140 ;
        RECT 103.780 173.400 104.860 173.700 ;
        RECT 112.060 173.400 113.140 173.700 ;
        RECT 104.170 171.940 104.470 173.400 ;
        RECT 105.940 172.960 107.020 173.260 ;
        RECT 109.900 172.960 110.980 173.260 ;
        RECT 106.330 172.380 106.630 172.960 ;
        RECT 110.290 172.380 110.590 172.960 ;
        RECT 105.940 172.080 110.980 172.380 ;
        RECT 103.780 171.640 104.860 171.940 ;
        RECT 104.170 170.180 104.470 171.640 ;
        RECT 105.940 171.200 107.020 171.500 ;
        RECT 106.330 170.660 106.630 171.200 ;
        RECT 106.100 170.620 107.020 170.660 ;
        RECT 105.940 170.320 107.020 170.620 ;
        RECT 103.780 169.880 104.860 170.180 ;
        RECT 104.170 168.420 104.470 169.880 ;
        RECT 105.940 169.440 107.020 169.740 ;
        RECT 106.330 168.900 106.630 169.440 ;
        RECT 109.300 169.130 109.600 172.080 ;
        RECT 112.450 171.940 112.750 173.400 ;
        RECT 112.060 171.640 113.140 171.940 ;
        RECT 110.060 171.500 110.980 171.540 ;
        RECT 109.900 171.200 110.980 171.500 ;
        RECT 110.290 170.660 110.590 171.200 ;
        RECT 110.060 170.620 110.980 170.660 ;
        RECT 109.900 170.320 110.980 170.620 ;
        RECT 112.450 170.180 112.750 171.640 ;
        RECT 112.060 169.880 113.140 170.180 ;
        RECT 109.900 169.440 110.980 169.740 ;
        RECT 106.100 168.860 107.020 168.900 ;
        RECT 109.145 168.860 109.600 169.130 ;
        RECT 110.290 168.860 110.590 169.440 ;
        RECT 105.940 168.560 110.980 168.860 ;
        RECT 103.780 168.120 104.860 168.420 ;
        RECT 109.145 168.210 109.485 168.560 ;
        RECT 112.450 168.420 112.750 169.880 ;
        RECT 111.460 168.120 113.140 168.420 ;
        RECT 106.100 167.980 107.020 168.020 ;
        RECT 110.060 167.980 110.980 168.020 ;
        RECT 105.940 167.680 107.020 167.980 ;
        RECT 109.900 167.680 110.980 167.980 ;
        RECT 106.100 167.100 107.020 167.140 ;
        RECT 110.060 167.100 110.980 167.140 ;
        RECT 105.940 166.800 107.020 167.100 ;
        RECT 109.900 166.800 110.980 167.100 ;
        RECT 103.780 166.360 104.860 166.660 ;
        RECT 104.170 164.900 104.470 166.360 ;
        RECT 105.940 165.920 107.020 166.220 ;
        RECT 109.900 165.920 110.980 166.220 ;
        RECT 106.330 165.340 106.630 165.920 ;
        RECT 110.290 165.340 110.590 165.920 ;
        RECT 105.940 165.040 110.980 165.340 ;
        RECT 103.780 164.600 104.860 164.900 ;
        RECT 104.170 163.140 104.470 164.600 ;
        RECT 105.940 164.160 107.020 164.460 ;
        RECT 106.330 163.620 106.630 164.160 ;
        RECT 106.100 163.580 107.020 163.620 ;
        RECT 105.940 163.280 107.020 163.580 ;
        RECT 103.780 162.840 104.860 163.140 ;
        RECT 104.170 161.380 104.470 162.840 ;
        RECT 105.940 162.400 107.020 162.700 ;
        RECT 106.330 161.820 106.630 162.400 ;
        RECT 109.300 161.820 109.600 165.040 ;
        RECT 110.060 164.460 110.980 164.500 ;
        RECT 109.900 164.160 110.980 164.460 ;
        RECT 110.290 163.620 110.590 164.160 ;
        RECT 110.060 163.580 110.980 163.620 ;
        RECT 109.900 163.280 110.980 163.580 ;
        RECT 109.900 162.400 110.980 162.700 ;
        RECT 110.290 161.820 110.590 162.400 ;
        RECT 111.460 161.820 111.760 168.120 ;
        RECT 112.140 168.080 113.060 168.120 ;
        RECT 112.060 166.360 113.140 166.660 ;
        RECT 112.450 164.900 112.750 166.360 ;
        RECT 112.060 164.600 113.140 164.900 ;
        RECT 112.450 163.140 112.750 164.600 ;
        RECT 112.060 162.840 113.140 163.140 ;
        RECT 105.940 161.520 111.760 161.820 ;
        RECT 112.450 161.380 112.750 162.840 ;
        RECT 103.780 161.080 105.460 161.380 ;
        RECT 112.060 161.080 113.140 161.380 ;
        RECT 105.160 160.060 105.460 161.080 ;
        RECT 106.100 160.940 107.020 160.980 ;
        RECT 110.060 160.940 110.980 160.980 ;
        RECT 105.940 160.640 107.020 160.940 ;
        RECT 109.900 160.640 110.980 160.940 ;
        RECT 105.160 159.760 110.980 160.060 ;
        RECT 103.780 159.620 104.700 159.660 ;
        RECT 112.220 159.620 113.140 159.660 ;
        RECT 103.180 159.320 104.860 159.620 ;
        RECT 112.060 159.320 113.140 159.620 ;
        RECT 103.180 154.340 103.480 159.320 ;
        RECT 104.170 157.860 104.470 159.320 ;
        RECT 105.940 158.880 107.020 159.180 ;
        RECT 109.900 158.880 110.980 159.180 ;
        RECT 106.330 158.300 106.630 158.880 ;
        RECT 110.290 158.300 110.590 158.880 ;
        RECT 105.940 158.000 107.020 158.300 ;
        RECT 109.900 158.000 110.980 158.300 ;
        RECT 103.780 157.560 104.860 157.860 ;
        RECT 111.460 157.560 113.140 157.860 ;
        RECT 104.170 156.100 104.470 157.560 ;
        RECT 105.940 157.120 107.020 157.420 ;
        RECT 109.900 157.120 110.980 157.420 ;
        RECT 106.330 156.540 106.630 157.120 ;
        RECT 110.290 156.540 110.590 157.120 ;
        RECT 105.940 156.240 107.020 156.540 ;
        RECT 109.900 156.240 110.980 156.540 ;
        RECT 103.780 155.800 104.860 156.100 ;
        RECT 106.100 155.660 107.020 155.700 ;
        RECT 110.060 155.660 110.980 155.700 ;
        RECT 105.940 155.360 107.020 155.660 ;
        RECT 109.900 155.360 110.980 155.660 ;
        RECT 110.060 154.780 110.980 154.820 ;
        RECT 105.940 154.480 110.980 154.780 ;
        RECT 103.180 154.040 104.860 154.340 ;
        RECT 103.180 142.020 103.480 154.040 ;
        RECT 104.170 152.580 104.470 154.040 ;
        RECT 105.940 153.600 107.020 153.900 ;
        RECT 109.900 153.600 110.980 153.900 ;
        RECT 106.330 153.020 106.630 153.600 ;
        RECT 110.290 153.020 110.590 153.600 ;
        RECT 105.940 152.720 107.020 153.020 ;
        RECT 109.900 152.720 110.980 153.020 ;
        RECT 111.460 152.580 111.760 157.560 ;
        RECT 112.060 156.100 112.980 156.140 ;
        RECT 112.060 155.800 113.740 156.100 ;
        RECT 112.220 154.340 113.140 154.380 ;
        RECT 112.060 154.040 113.140 154.340 ;
        RECT 103.780 152.280 104.860 152.580 ;
        RECT 111.460 152.280 113.140 152.580 ;
        RECT 104.170 150.820 104.470 152.280 ;
        RECT 105.940 151.840 107.020 152.140 ;
        RECT 109.900 151.840 110.980 152.140 ;
        RECT 106.330 151.260 106.630 151.840 ;
        RECT 110.290 151.260 110.590 151.840 ;
        RECT 105.940 150.960 107.020 151.260 ;
        RECT 109.900 150.960 110.980 151.260 ;
        RECT 103.780 150.520 104.860 150.820 ;
        RECT 106.100 150.380 107.020 150.420 ;
        RECT 110.060 150.380 110.980 150.420 ;
        RECT 105.940 150.080 107.020 150.380 ;
        RECT 109.900 150.080 110.980 150.380 ;
        RECT 111.460 149.500 111.760 152.280 ;
        RECT 112.060 150.820 112.980 150.860 ;
        RECT 112.060 150.520 113.140 150.820 ;
        RECT 105.940 149.200 111.760 149.500 ;
        RECT 103.780 148.760 104.860 149.060 ;
        RECT 112.060 148.760 113.140 149.060 ;
        RECT 106.100 148.620 107.020 148.660 ;
        RECT 110.060 148.620 110.980 148.660 ;
        RECT 105.940 148.320 107.020 148.620 ;
        RECT 109.900 148.320 110.980 148.620 ;
        RECT 111.460 148.460 112.360 148.760 ;
        RECT 106.100 147.740 107.020 147.780 ;
        RECT 111.460 147.740 111.760 148.460 ;
        RECT 105.940 147.440 107.020 147.740 ;
        RECT 107.320 147.440 111.760 147.740 ;
        RECT 103.780 147.000 105.640 147.300 ;
        RECT 103.780 145.240 104.860 145.540 ;
        RECT 103.780 143.480 104.860 143.780 ;
        RECT 103.180 141.720 104.860 142.020 ;
        RECT 105.340 141.580 105.640 147.000 ;
        RECT 105.940 146.560 107.020 146.860 ;
        RECT 106.330 145.980 106.630 146.560 ;
        RECT 105.940 145.680 107.020 145.980 ;
        RECT 105.940 144.800 107.020 145.100 ;
        RECT 106.330 144.220 106.630 144.800 ;
        RECT 105.940 143.920 107.020 144.220 ;
        RECT 106.100 143.340 107.020 143.380 ;
        RECT 107.320 143.340 107.620 147.440 ;
        RECT 112.060 147.000 113.140 147.300 ;
        RECT 110.060 146.860 110.980 146.900 ;
        RECT 109.900 146.560 110.980 146.860 ;
        RECT 110.060 145.980 110.980 146.020 ;
        RECT 109.900 145.680 110.980 145.980 ;
        RECT 112.060 145.540 112.980 145.580 ;
        RECT 112.060 145.240 113.140 145.540 ;
        RECT 105.940 143.040 107.620 143.340 ;
        RECT 109.300 144.800 110.980 145.100 ;
        RECT 109.300 144.220 109.600 144.800 ;
        RECT 109.300 143.920 110.980 144.220 ;
        RECT 106.100 142.460 107.020 142.500 ;
        RECT 105.940 142.160 107.020 142.460 ;
        RECT 109.300 142.460 109.600 143.920 ;
        RECT 113.440 143.780 113.740 155.800 ;
        RECT 112.060 143.480 113.740 143.780 ;
        RECT 110.060 143.340 110.980 143.380 ;
        RECT 109.900 143.040 110.980 143.340 ;
        RECT 109.300 142.160 110.980 142.460 ;
        RECT 112.220 142.020 113.140 142.060 ;
        RECT 112.060 141.720 113.140 142.020 ;
        RECT 105.340 141.280 110.980 141.580 ;
        RECT 106.100 140.700 107.020 140.740 ;
        RECT 110.060 140.700 110.980 140.740 ;
        RECT 105.340 140.400 107.020 140.700 ;
        RECT 109.900 140.400 111.760 140.700 ;
        RECT 105.340 140.260 105.640 140.400 ;
        RECT 98.680 139.960 105.640 140.260 ;
        RECT 93.340 139.820 94.260 139.860 ;
        RECT 97.300 139.820 98.220 139.860 ;
        RECT 98.680 139.820 98.980 139.960 ;
        RECT 92.560 139.520 94.420 139.820 ;
        RECT 97.300 139.520 98.980 139.820 ;
        RECT 101.620 139.010 102.700 139.960 ;
        RECT 105.340 139.820 105.640 139.960 ;
        RECT 111.460 140.260 111.760 140.400 ;
        RECT 114.220 140.260 115.300 208.600 ;
        RECT 117.760 208.460 118.060 208.600 ;
        RECT 123.880 208.900 124.180 209.040 ;
        RECT 126.820 208.900 127.900 209.850 ;
        RECT 123.880 208.600 127.900 208.900 ;
        RECT 118.540 208.460 119.460 208.500 ;
        RECT 122.500 208.460 123.420 208.500 ;
        RECT 123.880 208.460 124.180 208.600 ;
        RECT 117.760 208.160 119.620 208.460 ;
        RECT 122.500 208.160 124.180 208.460 ;
        RECT 116.380 207.140 117.300 207.370 ;
        RECT 118.540 207.280 124.180 207.580 ;
        RECT 116.380 206.840 117.460 207.140 ;
        RECT 118.540 206.700 119.460 206.740 ;
        RECT 122.500 206.700 123.420 206.740 ;
        RECT 118.540 206.400 119.620 206.700 ;
        RECT 122.500 206.400 123.580 206.700 ;
        RECT 118.540 205.820 119.460 205.860 ;
        RECT 118.540 205.520 119.620 205.820 ;
        RECT 119.920 205.520 123.580 205.820 ;
        RECT 116.380 205.080 117.460 205.380 ;
        RECT 119.920 204.940 120.220 205.520 ;
        RECT 117.940 204.640 120.220 204.940 ;
        RECT 122.500 204.640 123.580 204.940 ;
        RECT 116.380 203.320 117.460 203.620 ;
        RECT 116.380 201.560 117.460 201.860 ;
        RECT 117.940 200.100 118.240 204.640 ;
        RECT 119.920 204.060 120.220 204.640 ;
        RECT 122.890 204.060 123.190 204.640 ;
        RECT 118.540 203.760 120.220 204.060 ;
        RECT 122.500 203.760 123.580 204.060 ;
        RECT 118.540 203.180 119.460 203.220 ;
        RECT 122.500 203.180 123.420 203.220 ;
        RECT 118.540 202.880 119.620 203.180 ;
        RECT 122.500 202.880 123.580 203.180 ;
        RECT 118.540 202.300 119.460 202.340 ;
        RECT 122.500 202.300 123.420 202.340 ;
        RECT 118.540 202.000 120.220 202.300 ;
        RECT 122.500 202.000 123.580 202.300 ;
        RECT 119.920 201.420 120.220 202.000 ;
        RECT 123.880 201.860 124.180 207.280 ;
        RECT 124.660 206.840 125.740 207.140 ;
        RECT 124.740 205.380 125.660 205.420 ;
        RECT 124.660 205.080 125.740 205.380 ;
        RECT 124.660 203.620 125.580 203.660 ;
        RECT 124.660 203.320 125.740 203.620 ;
        RECT 123.880 201.560 125.740 201.860 ;
        RECT 118.540 201.120 119.620 201.420 ;
        RECT 119.920 201.120 123.580 201.420 ;
        RECT 118.930 200.540 119.230 201.120 ;
        RECT 119.920 200.540 120.220 201.120 ;
        RECT 118.540 200.240 119.620 200.540 ;
        RECT 119.920 200.240 123.580 200.540 ;
        RECT 116.380 199.800 118.240 200.100 ;
        RECT 124.660 199.800 125.740 200.100 ;
        RECT 118.540 199.660 119.460 199.700 ;
        RECT 122.500 199.660 123.420 199.700 ;
        RECT 118.540 199.360 119.620 199.660 ;
        RECT 122.500 199.360 123.580 199.660 ;
        RECT 117.760 198.480 123.580 198.780 ;
        RECT 116.380 198.340 117.300 198.380 ;
        RECT 116.380 198.040 117.460 198.340 ;
        RECT 117.760 196.580 118.060 198.480 ;
        RECT 124.660 198.040 125.740 198.340 ;
        RECT 118.540 197.900 119.460 197.940 ;
        RECT 122.500 197.900 123.420 197.940 ;
        RECT 118.540 197.600 119.620 197.900 ;
        RECT 122.500 197.600 123.580 197.900 ;
        RECT 118.540 196.720 124.180 197.020 ;
        RECT 115.780 196.280 118.060 196.580 ;
        RECT 115.780 173.700 116.080 196.280 ;
        RECT 122.890 196.140 123.190 196.720 ;
        RECT 123.880 196.580 124.180 196.720 ;
        RECT 123.880 196.280 125.740 196.580 ;
        RECT 118.540 195.840 119.620 196.140 ;
        RECT 122.500 195.840 123.580 196.140 ;
        RECT 118.930 195.260 119.230 195.840 ;
        RECT 122.890 195.260 123.190 195.840 ;
        RECT 118.540 194.960 119.620 195.260 ;
        RECT 122.500 194.960 123.580 195.260 ;
        RECT 116.380 194.520 117.460 194.820 ;
        RECT 116.770 193.060 117.070 194.520 ;
        RECT 118.930 194.380 119.230 194.960 ;
        RECT 122.890 194.380 123.190 194.960 ;
        RECT 125.050 194.820 125.350 196.280 ;
        RECT 124.660 194.520 125.740 194.820 ;
        RECT 118.540 194.080 119.620 194.380 ;
        RECT 122.500 194.080 123.580 194.380 ;
        RECT 118.930 193.500 119.230 194.080 ;
        RECT 122.890 193.500 123.190 194.080 ;
        RECT 118.540 193.200 119.620 193.500 ;
        RECT 122.500 193.200 123.580 193.500 ;
        RECT 116.380 192.760 117.460 193.060 ;
        RECT 116.770 191.300 117.070 192.760 ;
        RECT 118.930 192.620 119.230 193.200 ;
        RECT 122.890 192.620 123.190 193.200 ;
        RECT 125.050 193.060 125.350 194.520 ;
        RECT 124.660 192.760 125.740 193.060 ;
        RECT 118.540 192.320 119.620 192.620 ;
        RECT 122.500 192.320 123.580 192.620 ;
        RECT 118.930 191.740 119.230 192.320 ;
        RECT 122.890 191.740 123.190 192.320 ;
        RECT 118.540 191.440 119.620 191.740 ;
        RECT 122.500 191.440 123.580 191.740 ;
        RECT 116.380 191.000 117.460 191.300 ;
        RECT 116.770 189.540 117.070 191.000 ;
        RECT 118.930 190.860 119.230 191.440 ;
        RECT 122.890 190.860 123.190 191.440 ;
        RECT 125.050 191.300 125.350 192.760 ;
        RECT 124.660 191.000 125.740 191.300 ;
        RECT 118.540 190.560 119.620 190.860 ;
        RECT 122.500 190.560 123.580 190.860 ;
        RECT 118.930 189.980 119.230 190.560 ;
        RECT 122.890 189.980 123.190 190.560 ;
        RECT 118.540 189.680 119.620 189.980 ;
        RECT 122.500 189.680 123.580 189.980 ;
        RECT 116.380 189.240 117.460 189.540 ;
        RECT 116.770 187.820 117.070 189.240 ;
        RECT 118.930 189.100 119.230 189.680 ;
        RECT 122.890 189.100 123.190 189.680 ;
        RECT 125.050 189.540 125.350 191.000 ;
        RECT 124.660 189.240 125.740 189.540 ;
        RECT 118.540 188.800 119.620 189.100 ;
        RECT 122.500 188.800 123.580 189.100 ;
        RECT 118.930 188.220 119.230 188.800 ;
        RECT 122.890 188.220 123.190 188.800 ;
        RECT 118.540 187.920 119.620 188.220 ;
        RECT 122.500 187.920 123.580 188.220 ;
        RECT 116.540 187.780 117.460 187.820 ;
        RECT 116.380 187.480 117.460 187.780 ;
        RECT 118.930 187.340 119.230 187.920 ;
        RECT 122.890 187.340 123.190 187.920 ;
        RECT 125.050 187.780 125.350 189.240 ;
        RECT 124.660 187.480 125.740 187.780 ;
        RECT 118.540 187.040 119.620 187.340 ;
        RECT 122.500 187.040 123.580 187.340 ;
        RECT 118.930 186.460 119.230 187.040 ;
        RECT 122.890 186.500 123.190 187.040 ;
        RECT 122.500 186.460 123.420 186.500 ;
        RECT 118.540 186.160 120.220 186.460 ;
        RECT 122.500 186.160 123.580 186.460 ;
        RECT 116.380 186.020 117.300 186.060 ;
        RECT 116.380 185.720 117.460 186.020 ;
        RECT 118.540 185.580 119.460 185.620 ;
        RECT 119.920 185.580 120.220 186.160 ;
        RECT 124.660 185.720 125.740 186.020 ;
        RECT 118.540 185.280 119.620 185.580 ;
        RECT 119.920 185.280 123.580 185.580 ;
        RECT 122.500 184.700 123.420 184.740 ;
        RECT 118.540 184.400 122.200 184.700 ;
        RECT 122.500 184.400 123.580 184.700 ;
        RECT 116.380 183.960 117.460 184.260 ;
        RECT 118.540 183.520 119.620 183.820 ;
        RECT 118.930 182.940 119.230 183.520 ;
        RECT 121.900 182.940 122.200 184.400 ;
        RECT 124.660 183.960 125.740 184.260 ;
        RECT 122.500 183.520 123.580 183.820 ;
        RECT 122.890 182.940 123.190 183.520 ;
        RECT 118.540 182.640 120.220 182.940 ;
        RECT 116.540 182.500 117.460 182.540 ;
        RECT 116.380 182.200 117.460 182.500 ;
        RECT 116.770 180.740 117.070 182.200 ;
        RECT 118.540 181.760 119.620 182.060 ;
        RECT 118.930 181.180 119.230 181.760 ;
        RECT 117.940 180.880 119.620 181.180 ;
        RECT 116.380 180.440 117.460 180.740 ;
        RECT 116.770 178.980 117.070 180.440 ;
        RECT 116.380 178.680 117.460 178.980 ;
        RECT 116.770 177.220 117.070 178.680 ;
        RECT 117.940 177.660 118.240 180.880 ;
        RECT 118.540 180.000 119.620 180.300 ;
        RECT 118.930 179.420 119.230 180.000 ;
        RECT 119.920 179.420 120.220 182.640 ;
        RECT 118.540 179.120 120.220 179.420 ;
        RECT 121.900 182.640 123.580 182.940 ;
        RECT 121.900 179.420 122.200 182.640 ;
        RECT 125.050 182.500 125.350 183.960 ;
        RECT 124.660 182.200 125.740 182.500 ;
        RECT 122.500 182.060 123.420 182.100 ;
        RECT 122.500 181.760 123.580 182.060 ;
        RECT 122.890 181.220 123.190 181.760 ;
        RECT 122.500 181.180 123.420 181.220 ;
        RECT 122.500 180.880 123.580 181.180 ;
        RECT 125.050 180.740 125.350 182.200 ;
        RECT 123.880 180.440 125.740 180.740 ;
        RECT 122.500 180.300 123.420 180.340 ;
        RECT 122.500 180.000 123.580 180.300 ;
        RECT 122.890 179.420 123.190 180.000 ;
        RECT 121.900 179.120 123.580 179.420 ;
        RECT 118.540 178.240 119.620 178.540 ;
        RECT 118.930 177.660 119.230 178.240 ;
        RECT 117.940 177.360 119.620 177.660 ;
        RECT 116.380 176.920 117.460 177.220 ;
        RECT 116.770 175.460 117.070 176.920 ;
        RECT 116.380 175.160 117.460 175.460 ;
        RECT 117.940 174.140 118.240 177.360 ;
        RECT 118.540 176.480 119.620 176.780 ;
        RECT 118.930 175.900 119.230 176.480 ;
        RECT 119.920 175.900 120.220 179.120 ;
        RECT 122.500 178.540 123.420 178.580 ;
        RECT 122.500 178.240 123.580 178.540 ;
        RECT 122.890 177.700 123.190 178.240 ;
        RECT 122.500 177.660 123.420 177.700 ;
        RECT 122.500 177.360 123.580 177.660 ;
        RECT 122.500 176.480 123.580 176.780 ;
        RECT 122.890 175.900 123.190 176.480 ;
        RECT 118.540 175.600 123.580 175.900 ;
        RECT 122.500 175.020 123.420 175.060 ;
        RECT 118.540 174.720 119.620 175.020 ;
        RECT 122.500 174.720 123.580 175.020 ;
        RECT 118.930 174.140 119.230 174.720 ;
        RECT 122.890 174.180 123.190 174.720 ;
        RECT 122.500 174.140 123.420 174.180 ;
        RECT 117.940 173.840 120.220 174.140 ;
        RECT 122.500 173.840 123.580 174.140 ;
        RECT 115.780 173.400 117.460 173.700 ;
        RECT 115.780 154.340 116.080 173.400 ;
        RECT 116.380 171.640 117.460 171.940 ;
        RECT 116.770 170.180 117.070 171.640 ;
        RECT 116.380 169.880 117.460 170.180 ;
        RECT 116.380 168.120 117.460 168.420 ;
        RECT 116.770 166.660 117.070 168.120 ;
        RECT 116.380 166.360 117.460 166.660 ;
        RECT 116.380 164.600 117.460 164.900 ;
        RECT 116.380 162.840 117.460 163.140 ;
        RECT 116.770 161.380 117.070 162.840 ;
        RECT 117.940 161.820 118.240 173.840 ;
        RECT 118.540 173.260 119.460 173.300 ;
        RECT 119.920 173.260 120.220 173.840 ;
        RECT 118.540 172.960 119.620 173.260 ;
        RECT 119.920 172.960 123.580 173.260 ;
        RECT 118.540 172.380 119.460 172.420 ;
        RECT 122.500 172.380 123.420 172.420 ;
        RECT 118.540 172.080 119.620 172.380 ;
        RECT 122.500 172.080 123.580 172.380 ;
        RECT 118.540 171.200 123.580 171.500 ;
        RECT 119.920 170.620 120.220 171.200 ;
        RECT 122.500 170.620 123.420 170.660 ;
        RECT 118.540 170.320 123.580 170.620 ;
        RECT 123.880 170.180 124.180 180.440 ;
        RECT 124.660 178.680 126.340 178.980 ;
        RECT 124.660 177.220 125.580 177.260 ;
        RECT 124.660 176.920 125.740 177.220 ;
        RECT 126.040 175.460 126.340 178.680 ;
        RECT 124.660 175.160 126.340 175.460 ;
        RECT 126.040 173.700 126.340 175.160 ;
        RECT 124.660 173.400 126.340 173.700 ;
        RECT 124.660 171.640 125.740 171.940 ;
        RECT 125.050 170.180 125.350 171.640 ;
        RECT 123.880 169.880 125.740 170.180 ;
        RECT 118.540 169.740 119.460 169.780 ;
        RECT 122.500 169.740 123.420 169.780 ;
        RECT 118.540 169.440 119.620 169.740 ;
        RECT 122.500 169.440 123.580 169.740 ;
        RECT 118.540 168.860 119.460 168.900 ;
        RECT 122.500 168.860 123.420 168.900 ;
        RECT 118.540 168.560 119.620 168.860 ;
        RECT 122.500 168.560 123.580 168.860 ;
        RECT 118.540 167.680 123.580 167.980 ;
        RECT 118.620 167.100 119.540 167.330 ;
        RECT 119.920 167.100 120.220 167.680 ;
        RECT 118.540 166.800 123.580 167.100 ;
        RECT 118.540 166.220 119.460 166.260 ;
        RECT 122.500 166.220 123.420 166.260 ;
        RECT 118.540 165.920 119.620 166.220 ;
        RECT 122.500 165.920 123.580 166.220 ;
        RECT 122.500 165.340 123.420 165.380 ;
        RECT 118.540 165.040 122.200 165.340 ;
        RECT 122.500 165.040 123.580 165.340 ;
        RECT 118.540 164.160 119.620 164.460 ;
        RECT 118.930 163.580 119.230 164.160 ;
        RECT 121.900 163.580 122.200 165.040 ;
        RECT 123.880 164.460 124.180 169.880 ;
        RECT 124.660 168.120 125.740 168.420 ;
        RECT 125.050 166.700 125.350 168.120 ;
        RECT 124.660 166.660 125.580 166.700 ;
        RECT 124.660 166.360 125.740 166.660 ;
        RECT 124.660 164.600 125.740 164.900 ;
        RECT 122.500 164.160 124.180 164.460 ;
        RECT 122.890 163.580 123.190 164.160 ;
        RECT 118.540 163.280 120.220 163.580 ;
        RECT 118.540 162.400 119.620 162.700 ;
        RECT 118.930 161.820 119.230 162.400 ;
        RECT 117.940 161.520 119.620 161.820 ;
        RECT 116.380 161.080 117.460 161.380 ;
        RECT 116.770 159.620 117.070 161.080 ;
        RECT 116.380 159.320 117.460 159.620 ;
        RECT 116.770 157.860 117.070 159.320 ;
        RECT 117.940 158.300 118.240 161.520 ;
        RECT 118.540 160.640 119.620 160.940 ;
        RECT 118.930 160.060 119.230 160.640 ;
        RECT 119.920 160.060 120.220 163.280 ;
        RECT 118.540 159.760 120.220 160.060 ;
        RECT 121.900 163.280 123.580 163.580 ;
        RECT 121.900 160.060 122.200 163.280 ;
        RECT 125.050 163.180 125.350 164.600 ;
        RECT 124.660 163.140 125.580 163.180 ;
        RECT 124.660 162.840 125.740 163.140 ;
        RECT 122.500 162.700 123.420 162.740 ;
        RECT 122.500 162.400 123.580 162.700 ;
        RECT 122.890 161.860 123.190 162.400 ;
        RECT 122.500 161.820 123.420 161.860 ;
        RECT 122.500 161.520 123.580 161.820 ;
        RECT 125.050 161.380 125.350 162.840 ;
        RECT 124.660 161.080 125.740 161.380 ;
        RECT 122.500 160.640 123.580 160.940 ;
        RECT 122.890 160.060 123.190 160.640 ;
        RECT 121.900 159.760 123.580 160.060 ;
        RECT 118.540 158.880 119.620 159.180 ;
        RECT 118.930 158.300 119.230 158.880 ;
        RECT 117.940 158.000 119.620 158.300 ;
        RECT 116.380 157.560 117.460 157.860 ;
        RECT 116.770 156.140 117.070 157.560 ;
        RECT 116.540 156.100 117.460 156.140 ;
        RECT 116.380 155.800 117.460 156.100 ;
        RECT 117.940 154.780 118.240 158.000 ;
        RECT 118.540 157.120 119.620 157.420 ;
        RECT 118.930 156.540 119.230 157.120 ;
        RECT 119.920 156.540 120.220 159.760 ;
        RECT 124.660 159.320 126.340 159.620 ;
        RECT 122.500 159.180 123.420 159.220 ;
        RECT 122.500 158.880 123.580 159.180 ;
        RECT 122.890 158.340 123.190 158.880 ;
        RECT 122.500 158.300 123.420 158.340 ;
        RECT 122.500 158.000 123.580 158.300 ;
        RECT 124.660 157.860 125.580 157.900 ;
        RECT 124.660 157.560 125.740 157.860 ;
        RECT 122.500 157.120 123.580 157.420 ;
        RECT 122.890 156.540 123.190 157.120 ;
        RECT 118.540 156.240 123.580 156.540 ;
        RECT 126.040 156.100 126.340 159.320 ;
        RECT 124.660 155.800 126.340 156.100 ;
        RECT 122.500 155.660 123.420 155.700 ;
        RECT 118.540 155.360 119.620 155.660 ;
        RECT 122.500 155.360 123.580 155.660 ;
        RECT 118.930 154.780 119.230 155.360 ;
        RECT 122.890 154.820 123.190 155.360 ;
        RECT 122.500 154.780 123.420 154.820 ;
        RECT 117.940 154.480 120.220 154.780 ;
        RECT 122.500 154.480 123.580 154.780 ;
        RECT 115.780 154.040 117.460 154.340 ;
        RECT 115.780 152.580 116.080 154.040 ;
        RECT 118.540 153.900 119.460 153.940 ;
        RECT 119.920 153.900 120.220 154.480 ;
        RECT 126.040 154.340 126.340 155.800 ;
        RECT 124.660 154.040 126.340 154.340 ;
        RECT 118.540 153.600 119.620 153.900 ;
        RECT 119.920 153.600 123.580 153.900 ;
        RECT 118.540 152.720 124.180 153.020 ;
        RECT 115.780 152.280 117.460 152.580 ;
        RECT 122.890 152.140 123.190 152.720 ;
        RECT 123.880 152.580 124.180 152.720 ;
        RECT 123.880 152.280 125.740 152.580 ;
        RECT 118.540 151.840 119.620 152.140 ;
        RECT 122.500 151.840 123.580 152.140 ;
        RECT 118.930 151.260 119.230 151.840 ;
        RECT 122.890 151.260 123.190 151.840 ;
        RECT 118.540 150.960 119.620 151.260 ;
        RECT 122.500 150.960 123.580 151.260 ;
        RECT 116.540 150.820 117.460 150.860 ;
        RECT 116.380 150.520 117.460 150.820 ;
        RECT 116.770 149.060 117.070 150.520 ;
        RECT 118.930 150.380 119.230 150.960 ;
        RECT 122.890 150.380 123.190 150.960 ;
        RECT 125.050 150.820 125.350 152.280 ;
        RECT 124.660 150.520 125.740 150.820 ;
        RECT 118.540 150.080 119.620 150.380 ;
        RECT 122.500 150.080 123.580 150.380 ;
        RECT 118.930 149.500 119.230 150.080 ;
        RECT 122.890 149.500 123.190 150.080 ;
        RECT 118.540 149.200 119.620 149.500 ;
        RECT 122.500 149.200 123.580 149.500 ;
        RECT 116.380 148.760 117.460 149.060 ;
        RECT 116.770 147.300 117.070 148.760 ;
        RECT 118.930 148.620 119.230 149.200 ;
        RECT 122.890 148.620 123.190 149.200 ;
        RECT 125.050 149.060 125.350 150.520 ;
        RECT 124.660 148.760 125.740 149.060 ;
        RECT 118.540 148.320 119.620 148.620 ;
        RECT 122.500 148.320 123.580 148.620 ;
        RECT 118.930 147.740 119.230 148.320 ;
        RECT 122.890 147.740 123.190 148.320 ;
        RECT 118.540 147.440 119.620 147.740 ;
        RECT 122.500 147.440 123.580 147.740 ;
        RECT 116.380 147.000 117.460 147.300 ;
        RECT 116.770 145.540 117.070 147.000 ;
        RECT 118.930 146.860 119.230 147.440 ;
        RECT 122.890 146.860 123.190 147.440 ;
        RECT 125.050 147.300 125.350 148.760 ;
        RECT 124.660 147.000 125.740 147.300 ;
        RECT 118.540 146.560 119.620 146.860 ;
        RECT 122.500 146.560 123.580 146.860 ;
        RECT 118.930 145.980 119.230 146.560 ;
        RECT 122.890 145.980 123.190 146.560 ;
        RECT 118.540 145.680 119.620 145.980 ;
        RECT 122.500 145.680 123.580 145.980 ;
        RECT 116.380 145.240 117.460 145.540 ;
        RECT 116.770 143.780 117.070 145.240 ;
        RECT 118.930 145.100 119.230 145.680 ;
        RECT 122.890 145.100 123.190 145.680 ;
        RECT 125.050 145.540 125.350 147.000 ;
        RECT 124.660 145.240 125.740 145.540 ;
        RECT 118.540 144.800 119.620 145.100 ;
        RECT 122.500 144.800 123.580 145.100 ;
        RECT 118.930 144.220 119.230 144.800 ;
        RECT 122.890 144.220 123.190 144.800 ;
        RECT 118.540 143.920 119.620 144.220 ;
        RECT 122.500 143.920 123.580 144.220 ;
        RECT 116.380 143.480 117.460 143.780 ;
        RECT 118.930 143.340 119.230 143.920 ;
        RECT 122.890 143.340 123.190 143.920 ;
        RECT 125.050 143.780 125.350 145.240 ;
        RECT 124.660 143.480 125.740 143.780 ;
        RECT 118.540 143.040 119.620 143.340 ;
        RECT 122.500 143.040 123.580 143.340 ;
        RECT 118.930 142.460 119.230 143.040 ;
        RECT 122.890 142.500 123.190 143.040 ;
        RECT 122.500 142.460 123.420 142.500 ;
        RECT 118.540 142.160 120.220 142.460 ;
        RECT 122.500 142.160 123.580 142.460 ;
        RECT 116.380 142.020 117.300 142.060 ;
        RECT 116.380 141.720 117.460 142.020 ;
        RECT 118.540 141.580 119.460 141.620 ;
        RECT 119.920 141.580 120.220 142.160 ;
        RECT 124.660 141.720 125.740 142.020 ;
        RECT 118.540 141.280 119.620 141.580 ;
        RECT 119.920 141.280 123.580 141.580 ;
        RECT 118.540 140.700 119.460 140.740 ;
        RECT 122.500 140.700 123.420 140.740 ;
        RECT 117.760 140.400 119.620 140.700 ;
        RECT 122.500 140.400 124.180 140.700 ;
        RECT 117.760 140.260 118.060 140.400 ;
        RECT 111.460 139.960 118.060 140.260 ;
        RECT 106.100 139.820 107.020 139.860 ;
        RECT 110.060 139.820 110.980 139.860 ;
        RECT 111.460 139.820 111.760 139.960 ;
        RECT 105.340 139.520 107.020 139.820 ;
        RECT 109.900 139.520 111.760 139.820 ;
        RECT 114.220 139.010 115.300 139.960 ;
        RECT 117.760 139.820 118.060 139.960 ;
        RECT 123.880 140.260 124.180 140.400 ;
        RECT 126.820 140.260 127.900 208.600 ;
        RECT 123.880 139.960 127.900 140.260 ;
        RECT 118.540 139.820 119.460 139.860 ;
        RECT 122.500 139.820 123.420 139.860 ;
        RECT 123.880 139.820 124.180 139.960 ;
        RECT 117.760 139.520 119.620 139.820 ;
        RECT 122.500 139.520 124.180 139.820 ;
        RECT 126.820 139.010 127.900 139.960 ;
        RECT 23.480 109.500 23.820 109.730 ;
        RECT 117.300 109.500 117.640 109.730 ;
        RECT 13.320 109.120 58.160 109.500 ;
        RECT 58.460 109.120 59.760 109.500 ;
        RECT 81.360 109.120 82.660 109.500 ;
        RECT 82.960 109.120 127.800 109.500 ;
        RECT 23.480 108.810 23.820 109.120 ;
        RECT 117.300 108.810 117.640 109.120 ;
        RECT 22.080 106.440 22.420 106.670 ;
        RECT 26.280 106.440 26.620 106.670 ;
        RECT 44.480 106.440 44.820 106.670 ;
        RECT 48.680 106.440 49.020 106.670 ;
        RECT 92.100 106.440 92.440 106.670 ;
        RECT 96.300 106.440 96.640 106.670 ;
        RECT 114.500 106.440 114.840 106.670 ;
        RECT 118.700 106.440 119.040 106.670 ;
        RECT 13.320 106.060 58.160 106.440 ;
        RECT 58.460 106.060 59.760 106.440 ;
        RECT 81.360 106.060 82.660 106.440 ;
        RECT 82.960 106.060 127.800 106.440 ;
        RECT 22.080 105.750 22.420 106.060 ;
        RECT 26.280 105.750 26.620 106.060 ;
        RECT 44.480 105.750 44.820 106.060 ;
        RECT 48.680 105.750 49.020 106.060 ;
        RECT 92.100 105.750 92.440 106.060 ;
        RECT 96.300 105.750 96.640 106.060 ;
        RECT 114.500 105.750 114.840 106.060 ;
        RECT 118.700 105.750 119.040 106.060 ;
        RECT 19.280 103.380 19.620 103.610 ;
        RECT 20.680 103.380 21.020 103.610 ;
        RECT 27.680 103.380 28.020 103.610 ;
        RECT 29.080 103.380 29.420 103.610 ;
        RECT 41.680 103.380 42.020 103.610 ;
        RECT 43.080 103.380 43.420 103.610 ;
        RECT 50.080 103.380 50.420 103.610 ;
        RECT 51.480 103.380 51.820 103.610 ;
        RECT 89.300 103.380 89.640 103.610 ;
        RECT 90.700 103.380 91.040 103.610 ;
        RECT 97.700 103.380 98.040 103.610 ;
        RECT 99.100 103.380 99.440 103.610 ;
        RECT 111.700 103.380 112.040 103.610 ;
        RECT 113.100 103.380 113.440 103.610 ;
        RECT 120.100 103.380 120.440 103.610 ;
        RECT 121.500 103.380 121.840 103.610 ;
        RECT 13.320 103.000 58.160 103.380 ;
        RECT 58.460 103.000 59.760 103.380 ;
        RECT 81.360 103.000 82.660 103.380 ;
        RECT 82.960 103.000 127.800 103.380 ;
        RECT 19.280 102.690 19.620 103.000 ;
        RECT 20.680 102.690 21.020 103.000 ;
        RECT 27.680 102.690 28.020 103.000 ;
        RECT 29.080 102.690 29.420 103.000 ;
        RECT 41.680 102.690 42.020 103.000 ;
        RECT 43.080 102.690 43.420 103.000 ;
        RECT 50.080 102.690 50.420 103.000 ;
        RECT 51.480 102.690 51.820 103.000 ;
        RECT 89.300 102.690 89.640 103.000 ;
        RECT 90.700 102.690 91.040 103.000 ;
        RECT 97.700 102.690 98.040 103.000 ;
        RECT 99.100 102.690 99.440 103.000 ;
        RECT 111.700 102.690 112.040 103.000 ;
        RECT 113.100 102.690 113.440 103.000 ;
        RECT 120.100 102.690 120.440 103.000 ;
        RECT 121.500 102.690 121.840 103.000 ;
        RECT 24.880 100.320 25.220 100.550 ;
        RECT 45.880 100.320 46.220 100.550 ;
        RECT 94.900 100.320 95.240 100.550 ;
        RECT 115.900 100.320 116.240 100.550 ;
        RECT 13.320 99.940 58.160 100.320 ;
        RECT 58.460 99.940 59.760 100.320 ;
        RECT 81.360 99.940 82.660 100.320 ;
        RECT 82.960 99.940 127.800 100.320 ;
        RECT 24.880 99.630 25.220 99.940 ;
        RECT 45.880 99.630 46.220 99.940 ;
        RECT 94.900 99.630 95.240 99.940 ;
        RECT 115.900 99.630 116.240 99.940 ;
        RECT 13.680 97.260 14.020 97.490 ;
        RECT 15.080 97.260 15.420 97.490 ;
        RECT 16.480 97.260 16.820 97.490 ;
        RECT 17.880 97.260 18.220 97.490 ;
        RECT 30.480 97.260 30.820 97.490 ;
        RECT 31.880 97.260 32.220 97.490 ;
        RECT 33.280 97.260 33.620 97.490 ;
        RECT 34.680 97.260 35.020 97.490 ;
        RECT 36.080 97.260 36.420 97.490 ;
        RECT 37.480 97.260 37.820 97.490 ;
        RECT 38.880 97.260 39.220 97.490 ;
        RECT 40.280 97.260 40.620 97.490 ;
        RECT 52.880 97.260 53.220 97.490 ;
        RECT 54.280 97.260 54.620 97.490 ;
        RECT 55.680 97.260 56.020 97.490 ;
        RECT 57.080 97.260 57.420 97.490 ;
        RECT 83.700 97.260 84.040 97.490 ;
        RECT 85.100 97.260 85.440 97.490 ;
        RECT 86.500 97.260 86.840 97.490 ;
        RECT 87.900 97.260 88.240 97.490 ;
        RECT 100.500 97.260 100.840 97.490 ;
        RECT 101.900 97.260 102.240 97.490 ;
        RECT 103.300 97.260 103.640 97.490 ;
        RECT 104.700 97.260 105.040 97.490 ;
        RECT 106.100 97.260 106.440 97.490 ;
        RECT 107.500 97.260 107.840 97.490 ;
        RECT 108.900 97.260 109.240 97.490 ;
        RECT 110.300 97.260 110.640 97.490 ;
        RECT 122.900 97.260 123.240 97.490 ;
        RECT 124.300 97.260 124.640 97.490 ;
        RECT 125.700 97.260 126.040 97.490 ;
        RECT 127.100 97.260 127.440 97.490 ;
        RECT 13.320 96.880 58.160 97.260 ;
        RECT 58.460 96.880 59.760 97.260 ;
        RECT 81.360 96.880 82.660 97.260 ;
        RECT 82.960 96.880 127.800 97.260 ;
        RECT 13.680 96.570 14.020 96.880 ;
        RECT 15.080 96.570 15.420 96.880 ;
        RECT 16.480 96.570 16.820 96.880 ;
        RECT 17.880 96.570 18.220 96.880 ;
        RECT 30.480 96.570 30.820 96.880 ;
        RECT 31.880 96.570 32.220 96.880 ;
        RECT 33.280 96.570 33.620 96.880 ;
        RECT 34.680 96.570 35.020 96.880 ;
        RECT 36.080 96.570 36.420 96.880 ;
        RECT 37.480 96.570 37.820 96.880 ;
        RECT 38.880 96.570 39.220 96.880 ;
        RECT 40.280 96.570 40.620 96.880 ;
        RECT 52.880 96.570 53.220 96.880 ;
        RECT 54.280 96.570 54.620 96.880 ;
        RECT 55.680 96.570 56.020 96.880 ;
        RECT 57.080 96.570 57.420 96.880 ;
        RECT 83.700 96.570 84.040 96.880 ;
        RECT 85.100 96.570 85.440 96.880 ;
        RECT 86.500 96.570 86.840 96.880 ;
        RECT 87.900 96.570 88.240 96.880 ;
        RECT 100.500 96.570 100.840 96.880 ;
        RECT 101.900 96.570 102.240 96.880 ;
        RECT 103.300 96.570 103.640 96.880 ;
        RECT 104.700 96.570 105.040 96.880 ;
        RECT 106.100 96.570 106.440 96.880 ;
        RECT 107.500 96.570 107.840 96.880 ;
        RECT 108.900 96.570 109.240 96.880 ;
        RECT 110.300 96.570 110.640 96.880 ;
        RECT 122.900 96.570 123.240 96.880 ;
        RECT 124.300 96.570 124.640 96.880 ;
        RECT 125.700 96.570 126.040 96.880 ;
        RECT 127.100 96.570 127.440 96.880 ;
        RECT 47.280 94.200 47.620 94.430 ;
        RECT 93.500 94.200 93.840 94.430 ;
        RECT 13.320 93.820 58.160 94.200 ;
        RECT 58.460 93.820 59.760 94.200 ;
        RECT 81.360 93.820 82.660 94.200 ;
        RECT 82.960 93.820 127.800 94.200 ;
        RECT 47.280 93.510 47.620 93.820 ;
        RECT 93.500 93.510 93.840 93.820 ;
        RECT 23.480 92.100 23.820 92.330 ;
        RECT 117.300 92.100 117.640 92.330 ;
        RECT 13.320 91.720 58.160 92.100 ;
        RECT 58.460 91.720 59.760 92.100 ;
        RECT 81.360 91.720 82.660 92.100 ;
        RECT 82.960 91.720 127.800 92.100 ;
        RECT 23.480 91.410 23.820 91.720 ;
        RECT 117.300 91.410 117.640 91.720 ;
        RECT 22.080 89.040 22.420 89.270 ;
        RECT 26.280 89.040 26.620 89.270 ;
        RECT 44.480 89.040 44.820 89.270 ;
        RECT 48.680 89.040 49.020 89.270 ;
        RECT 92.100 89.040 92.440 89.270 ;
        RECT 96.300 89.040 96.640 89.270 ;
        RECT 114.500 89.040 114.840 89.270 ;
        RECT 118.700 89.040 119.040 89.270 ;
        RECT 13.320 88.660 58.160 89.040 ;
        RECT 58.460 88.660 59.760 89.040 ;
        RECT 81.360 88.660 82.660 89.040 ;
        RECT 82.960 88.660 127.800 89.040 ;
        RECT 22.080 88.350 22.420 88.660 ;
        RECT 26.280 88.350 26.620 88.660 ;
        RECT 44.480 88.350 44.820 88.660 ;
        RECT 48.680 88.350 49.020 88.660 ;
        RECT 92.100 88.350 92.440 88.660 ;
        RECT 96.300 88.350 96.640 88.660 ;
        RECT 114.500 88.350 114.840 88.660 ;
        RECT 118.700 88.350 119.040 88.660 ;
        RECT 19.280 85.980 19.620 86.210 ;
        RECT 20.680 85.980 21.020 86.210 ;
        RECT 27.680 85.980 28.020 86.210 ;
        RECT 29.080 85.980 29.420 86.210 ;
        RECT 41.680 85.980 42.020 86.210 ;
        RECT 43.080 85.980 43.420 86.210 ;
        RECT 50.080 85.980 50.420 86.210 ;
        RECT 51.480 85.980 51.820 86.210 ;
        RECT 89.300 85.980 89.640 86.210 ;
        RECT 90.700 85.980 91.040 86.210 ;
        RECT 97.700 85.980 98.040 86.210 ;
        RECT 99.100 85.980 99.440 86.210 ;
        RECT 111.700 85.980 112.040 86.210 ;
        RECT 113.100 85.980 113.440 86.210 ;
        RECT 120.100 85.980 120.440 86.210 ;
        RECT 121.500 85.980 121.840 86.210 ;
        RECT 13.320 85.600 58.160 85.980 ;
        RECT 58.460 85.600 59.760 85.980 ;
        RECT 81.360 85.600 82.660 85.980 ;
        RECT 82.960 85.600 127.800 85.980 ;
        RECT 19.280 85.290 19.620 85.600 ;
        RECT 20.680 85.290 21.020 85.600 ;
        RECT 27.680 85.290 28.020 85.600 ;
        RECT 29.080 85.290 29.420 85.600 ;
        RECT 41.680 85.290 42.020 85.600 ;
        RECT 43.080 85.290 43.420 85.600 ;
        RECT 50.080 85.290 50.420 85.600 ;
        RECT 51.480 85.290 51.820 85.600 ;
        RECT 89.300 85.290 89.640 85.600 ;
        RECT 90.700 85.290 91.040 85.600 ;
        RECT 97.700 85.290 98.040 85.600 ;
        RECT 99.100 85.290 99.440 85.600 ;
        RECT 111.700 85.290 112.040 85.600 ;
        RECT 113.100 85.290 113.440 85.600 ;
        RECT 120.100 85.290 120.440 85.600 ;
        RECT 121.500 85.290 121.840 85.600 ;
        RECT 24.880 82.920 25.220 83.150 ;
        RECT 45.880 82.920 46.220 83.150 ;
        RECT 94.900 82.920 95.240 83.150 ;
        RECT 115.900 82.920 116.240 83.150 ;
        RECT 13.320 82.540 58.160 82.920 ;
        RECT 58.460 82.540 59.760 82.920 ;
        RECT 81.360 82.540 82.660 82.920 ;
        RECT 82.960 82.540 127.800 82.920 ;
        RECT 24.880 82.230 25.220 82.540 ;
        RECT 45.880 82.230 46.220 82.540 ;
        RECT 94.900 82.230 95.240 82.540 ;
        RECT 115.900 82.230 116.240 82.540 ;
        RECT 13.680 79.860 14.020 80.090 ;
        RECT 15.080 79.860 15.420 80.090 ;
        RECT 16.480 79.860 16.820 80.090 ;
        RECT 17.880 79.860 18.220 80.090 ;
        RECT 30.480 79.860 30.820 80.090 ;
        RECT 31.880 79.860 32.220 80.090 ;
        RECT 33.280 79.860 33.620 80.090 ;
        RECT 34.680 79.860 35.020 80.090 ;
        RECT 36.080 79.860 36.420 80.090 ;
        RECT 37.480 79.860 37.820 80.090 ;
        RECT 38.880 79.860 39.220 80.090 ;
        RECT 40.280 79.860 40.620 80.090 ;
        RECT 52.880 79.860 53.220 80.090 ;
        RECT 54.280 79.860 54.620 80.090 ;
        RECT 55.680 79.860 56.020 80.090 ;
        RECT 57.080 79.860 57.420 80.090 ;
        RECT 83.700 79.860 84.040 80.090 ;
        RECT 85.100 79.860 85.440 80.090 ;
        RECT 86.500 79.860 86.840 80.090 ;
        RECT 87.900 79.860 88.240 80.090 ;
        RECT 100.500 79.860 100.840 80.090 ;
        RECT 101.900 79.860 102.240 80.090 ;
        RECT 103.300 79.860 103.640 80.090 ;
        RECT 104.700 79.860 105.040 80.090 ;
        RECT 106.100 79.860 106.440 80.090 ;
        RECT 107.500 79.860 107.840 80.090 ;
        RECT 108.900 79.860 109.240 80.090 ;
        RECT 110.300 79.860 110.640 80.090 ;
        RECT 122.900 79.860 123.240 80.090 ;
        RECT 124.300 79.860 124.640 80.090 ;
        RECT 125.700 79.860 126.040 80.090 ;
        RECT 127.100 79.860 127.440 80.090 ;
        RECT 13.320 79.480 58.160 79.860 ;
        RECT 58.460 79.480 59.760 79.860 ;
        RECT 81.360 79.480 82.660 79.860 ;
        RECT 82.960 79.480 127.800 79.860 ;
        RECT 13.680 79.170 14.020 79.480 ;
        RECT 15.080 79.170 15.420 79.480 ;
        RECT 16.480 79.170 16.820 79.480 ;
        RECT 17.880 79.170 18.220 79.480 ;
        RECT 30.480 79.170 30.820 79.480 ;
        RECT 31.880 79.170 32.220 79.480 ;
        RECT 33.280 79.170 33.620 79.480 ;
        RECT 34.680 79.170 35.020 79.480 ;
        RECT 36.080 79.170 36.420 79.480 ;
        RECT 37.480 79.170 37.820 79.480 ;
        RECT 38.880 79.170 39.220 79.480 ;
        RECT 40.280 79.170 40.620 79.480 ;
        RECT 52.880 79.170 53.220 79.480 ;
        RECT 54.280 79.170 54.620 79.480 ;
        RECT 55.680 79.170 56.020 79.480 ;
        RECT 57.080 79.170 57.420 79.480 ;
        RECT 83.700 79.170 84.040 79.480 ;
        RECT 85.100 79.170 85.440 79.480 ;
        RECT 86.500 79.170 86.840 79.480 ;
        RECT 87.900 79.170 88.240 79.480 ;
        RECT 100.500 79.170 100.840 79.480 ;
        RECT 101.900 79.170 102.240 79.480 ;
        RECT 103.300 79.170 103.640 79.480 ;
        RECT 104.700 79.170 105.040 79.480 ;
        RECT 106.100 79.170 106.440 79.480 ;
        RECT 107.500 79.170 107.840 79.480 ;
        RECT 108.900 79.170 109.240 79.480 ;
        RECT 110.300 79.170 110.640 79.480 ;
        RECT 122.900 79.170 123.240 79.480 ;
        RECT 124.300 79.170 124.640 79.480 ;
        RECT 125.700 79.170 126.040 79.480 ;
        RECT 127.100 79.170 127.440 79.480 ;
        RECT 47.280 76.800 47.620 77.030 ;
        RECT 93.500 76.800 93.840 77.030 ;
        RECT 13.320 76.420 58.160 76.800 ;
        RECT 58.460 76.420 59.760 76.800 ;
        RECT 81.360 76.420 82.660 76.800 ;
        RECT 82.960 76.420 127.800 76.800 ;
        RECT 47.280 76.110 47.620 76.420 ;
        RECT 93.500 76.110 93.840 76.420 ;
        RECT 23.480 74.700 23.820 74.930 ;
        RECT 117.300 74.700 117.640 74.930 ;
        RECT 13.320 74.320 58.160 74.700 ;
        RECT 58.460 74.320 59.760 74.700 ;
        RECT 81.360 74.320 82.660 74.700 ;
        RECT 82.960 74.320 127.800 74.700 ;
        RECT 23.480 74.010 23.820 74.320 ;
        RECT 117.300 74.010 117.640 74.320 ;
        RECT 22.080 71.640 22.420 71.870 ;
        RECT 26.280 71.640 26.620 71.870 ;
        RECT 44.480 71.640 44.820 71.870 ;
        RECT 48.680 71.640 49.020 71.870 ;
        RECT 92.100 71.640 92.440 71.870 ;
        RECT 96.300 71.640 96.640 71.870 ;
        RECT 114.500 71.640 114.840 71.870 ;
        RECT 118.700 71.640 119.040 71.870 ;
        RECT 13.320 71.260 58.160 71.640 ;
        RECT 58.460 71.260 59.760 71.640 ;
        RECT 81.360 71.260 82.660 71.640 ;
        RECT 82.960 71.260 127.800 71.640 ;
        RECT 22.080 70.950 22.420 71.260 ;
        RECT 26.280 70.950 26.620 71.260 ;
        RECT 44.480 70.950 44.820 71.260 ;
        RECT 48.680 70.950 49.020 71.260 ;
        RECT 92.100 70.950 92.440 71.260 ;
        RECT 96.300 70.950 96.640 71.260 ;
        RECT 114.500 70.950 114.840 71.260 ;
        RECT 118.700 70.950 119.040 71.260 ;
        RECT 19.280 68.580 19.620 68.810 ;
        RECT 20.680 68.580 21.020 68.810 ;
        RECT 27.680 68.580 28.020 68.810 ;
        RECT 29.080 68.580 29.420 68.810 ;
        RECT 41.680 68.580 42.020 68.810 ;
        RECT 43.080 68.580 43.420 68.810 ;
        RECT 50.080 68.580 50.420 68.810 ;
        RECT 51.480 68.580 51.820 68.810 ;
        RECT 89.300 68.580 89.640 68.810 ;
        RECT 90.700 68.580 91.040 68.810 ;
        RECT 97.700 68.580 98.040 68.810 ;
        RECT 99.100 68.580 99.440 68.810 ;
        RECT 111.700 68.580 112.040 68.810 ;
        RECT 113.100 68.580 113.440 68.810 ;
        RECT 120.100 68.580 120.440 68.810 ;
        RECT 121.500 68.580 121.840 68.810 ;
        RECT 13.320 68.200 58.160 68.580 ;
        RECT 58.460 68.200 59.760 68.580 ;
        RECT 81.360 68.200 82.660 68.580 ;
        RECT 82.960 68.200 127.800 68.580 ;
        RECT 19.280 67.890 19.620 68.200 ;
        RECT 20.680 67.890 21.020 68.200 ;
        RECT 27.680 67.890 28.020 68.200 ;
        RECT 29.080 67.890 29.420 68.200 ;
        RECT 41.680 67.890 42.020 68.200 ;
        RECT 43.080 67.890 43.420 68.200 ;
        RECT 50.080 67.890 50.420 68.200 ;
        RECT 51.480 67.890 51.820 68.200 ;
        RECT 89.300 67.890 89.640 68.200 ;
        RECT 90.700 67.890 91.040 68.200 ;
        RECT 97.700 67.890 98.040 68.200 ;
        RECT 99.100 67.890 99.440 68.200 ;
        RECT 111.700 67.890 112.040 68.200 ;
        RECT 113.100 67.890 113.440 68.200 ;
        RECT 120.100 67.890 120.440 68.200 ;
        RECT 121.500 67.890 121.840 68.200 ;
        RECT 24.880 65.520 25.220 65.750 ;
        RECT 45.880 65.520 46.220 65.750 ;
        RECT 94.900 65.520 95.240 65.750 ;
        RECT 115.900 65.520 116.240 65.750 ;
        RECT 13.320 65.140 58.160 65.520 ;
        RECT 58.460 65.140 59.760 65.520 ;
        RECT 81.360 65.140 82.660 65.520 ;
        RECT 82.960 65.140 127.800 65.520 ;
        RECT 24.880 64.830 25.220 65.140 ;
        RECT 45.880 64.830 46.220 65.140 ;
        RECT 94.900 64.830 95.240 65.140 ;
        RECT 115.900 64.830 116.240 65.140 ;
        RECT 13.680 62.460 14.020 62.690 ;
        RECT 15.080 62.460 15.420 62.690 ;
        RECT 16.480 62.460 16.820 62.690 ;
        RECT 17.880 62.460 18.220 62.690 ;
        RECT 30.480 62.460 30.820 62.690 ;
        RECT 31.880 62.460 32.220 62.690 ;
        RECT 33.280 62.460 33.620 62.690 ;
        RECT 34.680 62.460 35.020 62.690 ;
        RECT 36.080 62.460 36.420 62.690 ;
        RECT 37.480 62.460 37.820 62.690 ;
        RECT 38.880 62.460 39.220 62.690 ;
        RECT 40.280 62.460 40.620 62.690 ;
        RECT 52.880 62.460 53.220 62.690 ;
        RECT 54.280 62.460 54.620 62.690 ;
        RECT 55.680 62.460 56.020 62.690 ;
        RECT 57.080 62.460 57.420 62.690 ;
        RECT 83.700 62.460 84.040 62.690 ;
        RECT 85.100 62.460 85.440 62.690 ;
        RECT 86.500 62.460 86.840 62.690 ;
        RECT 87.900 62.460 88.240 62.690 ;
        RECT 100.500 62.460 100.840 62.690 ;
        RECT 101.900 62.460 102.240 62.690 ;
        RECT 103.300 62.460 103.640 62.690 ;
        RECT 104.700 62.460 105.040 62.690 ;
        RECT 106.100 62.460 106.440 62.690 ;
        RECT 107.500 62.460 107.840 62.690 ;
        RECT 108.900 62.460 109.240 62.690 ;
        RECT 110.300 62.460 110.640 62.690 ;
        RECT 122.900 62.460 123.240 62.690 ;
        RECT 124.300 62.460 124.640 62.690 ;
        RECT 125.700 62.460 126.040 62.690 ;
        RECT 127.100 62.460 127.440 62.690 ;
        RECT 13.320 62.080 58.160 62.460 ;
        RECT 58.460 62.080 59.760 62.460 ;
        RECT 81.360 62.080 82.660 62.460 ;
        RECT 82.960 62.080 127.800 62.460 ;
        RECT 13.680 61.770 14.020 62.080 ;
        RECT 15.080 61.770 15.420 62.080 ;
        RECT 16.480 61.770 16.820 62.080 ;
        RECT 17.880 61.770 18.220 62.080 ;
        RECT 30.480 61.770 30.820 62.080 ;
        RECT 31.880 61.770 32.220 62.080 ;
        RECT 33.280 61.770 33.620 62.080 ;
        RECT 34.680 61.770 35.020 62.080 ;
        RECT 36.080 61.770 36.420 62.080 ;
        RECT 37.480 61.770 37.820 62.080 ;
        RECT 38.880 61.770 39.220 62.080 ;
        RECT 40.280 61.770 40.620 62.080 ;
        RECT 52.880 61.770 53.220 62.080 ;
        RECT 54.280 61.770 54.620 62.080 ;
        RECT 55.680 61.770 56.020 62.080 ;
        RECT 57.080 61.770 57.420 62.080 ;
        RECT 83.700 61.770 84.040 62.080 ;
        RECT 85.100 61.770 85.440 62.080 ;
        RECT 86.500 61.770 86.840 62.080 ;
        RECT 87.900 61.770 88.240 62.080 ;
        RECT 100.500 61.770 100.840 62.080 ;
        RECT 101.900 61.770 102.240 62.080 ;
        RECT 103.300 61.770 103.640 62.080 ;
        RECT 104.700 61.770 105.040 62.080 ;
        RECT 106.100 61.770 106.440 62.080 ;
        RECT 107.500 61.770 107.840 62.080 ;
        RECT 108.900 61.770 109.240 62.080 ;
        RECT 110.300 61.770 110.640 62.080 ;
        RECT 122.900 61.770 123.240 62.080 ;
        RECT 124.300 61.770 124.640 62.080 ;
        RECT 125.700 61.770 126.040 62.080 ;
        RECT 127.100 61.770 127.440 62.080 ;
        RECT 47.280 59.400 47.620 59.630 ;
        RECT 59.420 59.400 59.760 59.670 ;
        RECT 13.320 59.020 58.160 59.400 ;
        RECT 58.460 59.020 59.760 59.400 ;
        RECT 47.280 58.710 47.620 59.020 ;
        RECT 59.420 58.750 59.760 59.020 ;
        RECT 81.360 59.400 81.700 59.670 ;
        RECT 93.500 59.400 93.840 59.630 ;
        RECT 81.360 59.020 82.660 59.400 ;
        RECT 82.960 59.020 127.800 59.400 ;
        RECT 81.360 58.750 81.700 59.020 ;
        RECT 93.500 58.710 93.840 59.020 ;
        RECT 23.480 57.300 23.820 57.530 ;
        RECT 117.300 57.300 117.640 57.530 ;
        RECT 13.320 56.920 58.160 57.300 ;
        RECT 58.460 56.920 59.760 57.300 ;
        RECT 81.360 56.920 82.660 57.300 ;
        RECT 82.960 56.920 127.800 57.300 ;
        RECT 23.480 56.610 23.820 56.920 ;
        RECT 117.300 56.610 117.640 56.920 ;
        RECT 22.080 54.240 22.420 54.470 ;
        RECT 26.280 54.240 26.620 54.470 ;
        RECT 44.480 54.240 44.820 54.470 ;
        RECT 48.680 54.240 49.020 54.470 ;
        RECT 92.100 54.240 92.440 54.470 ;
        RECT 96.300 54.240 96.640 54.470 ;
        RECT 114.500 54.240 114.840 54.470 ;
        RECT 118.700 54.240 119.040 54.470 ;
        RECT 13.320 53.860 58.160 54.240 ;
        RECT 58.460 53.860 59.760 54.240 ;
        RECT 81.360 53.860 82.660 54.240 ;
        RECT 82.960 53.860 127.800 54.240 ;
        RECT 22.080 53.550 22.420 53.860 ;
        RECT 26.280 53.550 26.620 53.860 ;
        RECT 44.480 53.550 44.820 53.860 ;
        RECT 48.680 53.550 49.020 53.860 ;
        RECT 92.100 53.550 92.440 53.860 ;
        RECT 96.300 53.550 96.640 53.860 ;
        RECT 114.500 53.550 114.840 53.860 ;
        RECT 118.700 53.550 119.040 53.860 ;
        RECT 19.280 51.180 19.620 51.410 ;
        RECT 20.680 51.180 21.020 51.410 ;
        RECT 27.680 51.180 28.020 51.410 ;
        RECT 29.080 51.180 29.420 51.410 ;
        RECT 41.680 51.180 42.020 51.410 ;
        RECT 43.080 51.180 43.420 51.410 ;
        RECT 50.080 51.180 50.420 51.410 ;
        RECT 51.480 51.180 51.820 51.410 ;
        RECT 89.300 51.180 89.640 51.410 ;
        RECT 90.700 51.180 91.040 51.410 ;
        RECT 97.700 51.180 98.040 51.410 ;
        RECT 99.100 51.180 99.440 51.410 ;
        RECT 111.700 51.180 112.040 51.410 ;
        RECT 113.100 51.180 113.440 51.410 ;
        RECT 120.100 51.180 120.440 51.410 ;
        RECT 121.500 51.180 121.840 51.410 ;
        RECT 13.320 50.800 58.160 51.180 ;
        RECT 58.460 50.800 59.760 51.180 ;
        RECT 81.360 50.800 82.660 51.180 ;
        RECT 82.960 50.800 127.800 51.180 ;
        RECT 19.280 50.490 19.620 50.800 ;
        RECT 20.680 50.490 21.020 50.800 ;
        RECT 27.680 50.490 28.020 50.800 ;
        RECT 29.080 50.490 29.420 50.800 ;
        RECT 41.680 50.490 42.020 50.800 ;
        RECT 43.080 50.490 43.420 50.800 ;
        RECT 50.080 50.490 50.420 50.800 ;
        RECT 51.480 50.490 51.820 50.800 ;
        RECT 89.300 50.490 89.640 50.800 ;
        RECT 90.700 50.490 91.040 50.800 ;
        RECT 97.700 50.490 98.040 50.800 ;
        RECT 99.100 50.490 99.440 50.800 ;
        RECT 111.700 50.490 112.040 50.800 ;
        RECT 113.100 50.490 113.440 50.800 ;
        RECT 120.100 50.490 120.440 50.800 ;
        RECT 121.500 50.490 121.840 50.800 ;
        RECT 24.880 48.120 25.220 48.350 ;
        RECT 45.880 48.120 46.220 48.350 ;
        RECT 94.900 48.120 95.240 48.350 ;
        RECT 115.900 48.120 116.240 48.350 ;
        RECT 13.320 47.740 58.160 48.120 ;
        RECT 58.460 47.740 59.760 48.120 ;
        RECT 81.360 47.740 82.660 48.120 ;
        RECT 82.960 47.740 127.800 48.120 ;
        RECT 24.880 47.430 25.220 47.740 ;
        RECT 45.880 47.430 46.220 47.740 ;
        RECT 94.900 47.430 95.240 47.740 ;
        RECT 115.900 47.430 116.240 47.740 ;
        RECT 13.680 45.060 14.020 45.290 ;
        RECT 15.080 45.060 15.420 45.290 ;
        RECT 16.480 45.060 16.820 45.290 ;
        RECT 17.880 45.060 18.220 45.290 ;
        RECT 30.480 45.060 30.820 45.290 ;
        RECT 31.880 45.060 32.220 45.290 ;
        RECT 33.280 45.060 33.620 45.290 ;
        RECT 34.680 45.060 35.020 45.290 ;
        RECT 36.080 45.060 36.420 45.290 ;
        RECT 37.480 45.060 37.820 45.290 ;
        RECT 38.880 45.060 39.220 45.290 ;
        RECT 40.280 45.060 40.620 45.290 ;
        RECT 52.880 45.060 53.220 45.290 ;
        RECT 54.280 45.060 54.620 45.290 ;
        RECT 55.680 45.060 56.020 45.290 ;
        RECT 57.080 45.060 57.420 45.290 ;
        RECT 83.700 45.060 84.040 45.290 ;
        RECT 85.100 45.060 85.440 45.290 ;
        RECT 86.500 45.060 86.840 45.290 ;
        RECT 87.900 45.060 88.240 45.290 ;
        RECT 100.500 45.060 100.840 45.290 ;
        RECT 101.900 45.060 102.240 45.290 ;
        RECT 103.300 45.060 103.640 45.290 ;
        RECT 104.700 45.060 105.040 45.290 ;
        RECT 106.100 45.060 106.440 45.290 ;
        RECT 107.500 45.060 107.840 45.290 ;
        RECT 108.900 45.060 109.240 45.290 ;
        RECT 110.300 45.060 110.640 45.290 ;
        RECT 122.900 45.060 123.240 45.290 ;
        RECT 124.300 45.060 124.640 45.290 ;
        RECT 125.700 45.060 126.040 45.290 ;
        RECT 127.100 45.060 127.440 45.290 ;
        RECT 13.320 44.680 58.160 45.060 ;
        RECT 58.460 44.680 59.760 45.060 ;
        RECT 81.360 44.680 82.660 45.060 ;
        RECT 82.960 44.680 127.800 45.060 ;
        RECT 13.680 44.370 14.020 44.680 ;
        RECT 15.080 44.370 15.420 44.680 ;
        RECT 16.480 44.370 16.820 44.680 ;
        RECT 17.880 44.370 18.220 44.680 ;
        RECT 30.480 44.370 30.820 44.680 ;
        RECT 31.880 44.370 32.220 44.680 ;
        RECT 33.280 44.370 33.620 44.680 ;
        RECT 34.680 44.370 35.020 44.680 ;
        RECT 36.080 44.370 36.420 44.680 ;
        RECT 37.480 44.370 37.820 44.680 ;
        RECT 38.880 44.370 39.220 44.680 ;
        RECT 40.280 44.370 40.620 44.680 ;
        RECT 52.880 44.370 53.220 44.680 ;
        RECT 54.280 44.370 54.620 44.680 ;
        RECT 55.680 44.370 56.020 44.680 ;
        RECT 57.080 44.370 57.420 44.680 ;
        RECT 83.700 44.370 84.040 44.680 ;
        RECT 85.100 44.370 85.440 44.680 ;
        RECT 86.500 44.370 86.840 44.680 ;
        RECT 87.900 44.370 88.240 44.680 ;
        RECT 100.500 44.370 100.840 44.680 ;
        RECT 101.900 44.370 102.240 44.680 ;
        RECT 103.300 44.370 103.640 44.680 ;
        RECT 104.700 44.370 105.040 44.680 ;
        RECT 106.100 44.370 106.440 44.680 ;
        RECT 107.500 44.370 107.840 44.680 ;
        RECT 108.900 44.370 109.240 44.680 ;
        RECT 110.300 44.370 110.640 44.680 ;
        RECT 122.900 44.370 123.240 44.680 ;
        RECT 124.300 44.370 124.640 44.680 ;
        RECT 125.700 44.370 126.040 44.680 ;
        RECT 127.100 44.370 127.440 44.680 ;
        RECT 47.280 42.000 47.620 42.230 ;
        RECT 93.500 42.000 93.840 42.230 ;
        RECT 13.320 41.620 58.160 42.000 ;
        RECT 58.460 41.620 59.760 42.000 ;
        RECT 81.360 41.620 82.660 42.000 ;
        RECT 82.960 41.620 127.800 42.000 ;
        RECT 47.280 41.310 47.620 41.620 ;
        RECT 93.500 41.310 93.840 41.620 ;
        RECT 13.600 38.540 49.240 38.980 ;
        RECT 13.600 37.660 48.520 38.100 ;
        RECT 13.600 36.340 13.960 37.660 ;
        RECT 48.880 37.220 49.240 38.540 ;
        RECT 14.320 36.780 49.240 37.220 ;
        RECT 13.600 35.900 48.520 36.340 ;
        RECT 13.600 34.580 13.960 35.900 ;
        RECT 48.880 35.460 49.240 36.780 ;
        RECT 14.320 35.020 49.240 35.460 ;
        RECT 92.080 38.540 127.720 38.980 ;
        RECT 92.080 37.220 92.440 38.540 ;
        RECT 92.800 37.660 127.720 38.100 ;
        RECT 92.080 36.780 127.000 37.220 ;
        RECT 92.080 35.460 92.440 36.780 ;
        RECT 127.360 36.340 127.720 37.660 ;
        RECT 92.800 35.900 127.720 36.340 ;
        RECT 92.080 35.020 127.000 35.460 ;
        RECT 127.360 34.580 127.720 35.900 ;
        RECT 13.600 34.140 49.240 34.580 ;
        RECT 92.080 34.140 127.720 34.580 ;
        RECT 13.600 33.260 49.240 33.700 ;
        RECT 13.600 32.380 48.520 32.820 ;
        RECT 13.600 31.060 13.960 32.380 ;
        RECT 48.880 31.940 49.240 33.260 ;
        RECT 92.080 33.260 127.720 33.700 ;
        RECT 14.320 31.500 49.240 31.940 ;
        RECT 13.600 30.620 48.520 31.060 ;
        RECT 13.600 29.300 13.960 30.620 ;
        RECT 48.880 30.180 49.240 31.500 ;
        RECT 14.320 29.740 49.240 30.180 ;
        RECT 50.320 31.870 51.400 32.820 ;
        RECT 54.800 32.310 55.720 32.350 ;
        RECT 58.760 32.310 59.680 32.350 ;
        RECT 54.040 32.010 55.720 32.310 ;
        RECT 58.600 32.010 60.460 32.310 ;
        RECT 54.040 31.870 54.340 32.010 ;
        RECT 50.320 31.570 54.340 31.870 ;
        RECT 13.600 28.860 49.240 29.300 ;
        RECT 13.600 27.980 49.240 28.420 ;
        RECT 13.600 27.100 48.520 27.540 ;
        RECT 13.600 25.780 13.960 27.100 ;
        RECT 48.880 26.660 49.240 27.980 ;
        RECT 14.320 26.220 49.240 26.660 ;
        RECT 13.600 25.340 48.520 25.780 ;
        RECT 13.600 24.020 13.960 25.340 ;
        RECT 48.880 24.900 49.240 26.220 ;
        RECT 14.320 24.460 49.240 24.900 ;
        RECT 50.320 28.350 51.400 31.570 ;
        RECT 54.040 31.430 54.340 31.570 ;
        RECT 60.160 31.870 60.460 32.010 ;
        RECT 62.920 31.870 64.000 32.820 ;
        RECT 60.160 31.570 64.000 31.870 ;
        RECT 54.800 31.430 55.720 31.470 ;
        RECT 58.760 31.430 59.680 31.470 ;
        RECT 60.160 31.430 60.460 31.570 ;
        RECT 54.040 31.130 55.720 31.430 ;
        RECT 58.600 31.130 60.460 31.430 ;
        RECT 58.760 30.550 59.680 30.590 ;
        RECT 54.040 30.250 55.720 30.550 ;
        RECT 58.600 30.250 59.680 30.550 ;
        RECT 54.040 30.110 54.340 30.250 ;
        RECT 52.480 29.810 54.340 30.110 ;
        RECT 60.760 29.810 61.840 30.110 ;
        RECT 54.800 29.670 55.720 29.710 ;
        RECT 58.760 29.670 59.680 29.710 ;
        RECT 54.640 29.370 55.720 29.670 ;
        RECT 58.600 29.370 59.680 29.670 ;
        RECT 54.800 28.790 55.720 28.830 ;
        RECT 58.760 28.790 59.680 28.830 ;
        RECT 54.040 28.490 55.720 28.790 ;
        RECT 58.600 28.490 60.460 28.790 ;
        RECT 54.040 28.350 54.340 28.490 ;
        RECT 50.320 28.050 54.340 28.350 ;
        RECT 13.600 23.580 49.240 24.020 ;
        RECT 13.600 22.700 49.240 23.140 ;
        RECT 13.600 21.820 48.520 22.260 ;
        RECT 13.600 20.500 13.960 21.820 ;
        RECT 48.880 21.380 49.240 22.700 ;
        RECT 14.320 20.940 49.240 21.380 ;
        RECT 13.600 20.060 48.520 20.500 ;
        RECT 13.600 18.740 13.960 20.060 ;
        RECT 48.880 19.620 49.240 20.940 ;
        RECT 14.320 19.180 49.240 19.620 ;
        RECT 13.600 18.300 49.240 18.740 ;
        RECT 13.600 17.420 49.240 17.860 ;
        RECT 13.600 16.540 48.520 16.980 ;
        RECT 13.600 15.220 13.960 16.540 ;
        RECT 48.880 16.100 49.240 17.420 ;
        RECT 14.320 15.660 49.240 16.100 ;
        RECT 13.600 14.780 48.520 15.220 ;
        RECT 13.600 13.460 13.960 14.780 ;
        RECT 48.880 14.340 49.240 15.660 ;
        RECT 14.320 13.900 49.240 14.340 ;
        RECT 50.320 14.270 51.400 28.050 ;
        RECT 54.040 27.910 54.340 28.050 ;
        RECT 60.160 28.350 60.460 28.490 ;
        RECT 62.920 28.350 64.000 31.570 ;
        RECT 60.160 28.050 64.000 28.350 ;
        RECT 54.800 27.910 55.720 27.950 ;
        RECT 58.760 27.910 59.680 27.950 ;
        RECT 60.160 27.910 60.460 28.050 ;
        RECT 54.040 27.610 55.720 27.910 ;
        RECT 58.600 27.610 60.460 27.910 ;
        RECT 54.800 27.030 55.720 27.240 ;
        RECT 54.640 26.730 55.720 27.030 ;
        RECT 58.600 26.730 60.460 27.030 ;
        RECT 60.160 26.590 60.460 26.730 ;
        RECT 52.480 26.290 53.560 26.590 ;
        RECT 60.160 26.290 61.840 26.590 ;
        RECT 54.800 26.150 55.720 26.190 ;
        RECT 58.760 26.150 59.680 26.190 ;
        RECT 54.640 25.850 55.720 26.150 ;
        RECT 58.600 25.850 59.680 26.150 ;
        RECT 54.800 25.270 55.720 25.310 ;
        RECT 58.680 25.270 59.600 25.310 ;
        RECT 54.640 24.970 55.720 25.270 ;
        RECT 58.000 24.970 59.680 25.270 ;
        RECT 52.480 24.530 54.340 24.830 ;
        RECT 52.480 22.770 53.560 23.070 ;
        RECT 54.040 22.630 54.340 24.530 ;
        RECT 54.640 24.090 55.720 24.390 ;
        RECT 55.030 23.550 55.330 24.090 ;
        RECT 54.800 23.510 55.720 23.550 ;
        RECT 54.640 23.210 55.720 23.510 ;
        RECT 58.000 22.630 58.300 24.970 ;
        RECT 60.920 24.830 61.840 24.870 ;
        RECT 60.760 24.530 61.840 24.830 ;
        RECT 58.600 24.090 59.680 24.390 ;
        RECT 58.990 23.510 59.290 24.090 ;
        RECT 58.600 23.210 59.680 23.510 ;
        RECT 60.920 23.070 61.840 23.110 ;
        RECT 60.760 22.770 61.840 23.070 ;
        RECT 58.760 22.630 59.680 22.670 ;
        RECT 54.040 22.330 58.300 22.630 ;
        RECT 58.600 22.330 59.680 22.630 ;
        RECT 58.760 21.750 59.680 21.790 ;
        RECT 54.640 21.450 59.680 21.750 ;
        RECT 51.880 21.010 53.560 21.310 ;
        RECT 60.160 21.010 61.840 21.310 ;
        RECT 51.880 17.790 52.180 21.010 ;
        RECT 54.800 20.870 55.720 20.910 ;
        RECT 54.640 20.570 59.680 20.870 ;
        RECT 55.030 19.990 55.330 20.570 ;
        RECT 58.990 19.990 59.290 20.570 ;
        RECT 54.640 19.690 55.720 19.990 ;
        RECT 58.600 19.690 59.680 19.990 ;
        RECT 52.640 19.550 53.560 19.590 ;
        RECT 52.480 19.250 53.560 19.550 ;
        RECT 54.800 19.110 55.720 19.150 ;
        RECT 58.760 19.110 59.680 19.150 ;
        RECT 54.640 18.810 55.720 19.110 ;
        RECT 58.600 18.810 59.680 19.110 ;
        RECT 55.030 18.270 55.330 18.810 ;
        RECT 58.990 18.270 59.290 18.810 ;
        RECT 54.800 18.230 55.720 18.270 ;
        RECT 58.760 18.230 59.680 18.270 ;
        RECT 54.640 17.930 55.720 18.230 ;
        RECT 58.600 17.930 59.680 18.230 ;
        RECT 52.640 17.790 53.560 17.830 ;
        RECT 51.880 17.490 53.560 17.790 ;
        RECT 60.160 17.350 60.460 21.010 ;
        RECT 60.760 19.250 61.840 19.550 ;
        RECT 61.150 17.790 61.450 19.250 ;
        RECT 60.760 17.490 61.840 17.790 ;
        RECT 54.640 17.050 60.460 17.350 ;
        RECT 54.800 16.470 55.720 16.510 ;
        RECT 58.760 16.470 59.680 16.700 ;
        RECT 54.640 16.170 59.680 16.470 ;
        RECT 60.840 16.030 61.760 16.070 ;
        RECT 52.480 15.730 53.560 16.030 ;
        RECT 60.760 15.730 61.840 16.030 ;
        RECT 54.800 15.590 55.720 15.630 ;
        RECT 58.760 15.590 59.680 15.630 ;
        RECT 54.640 15.290 55.720 15.590 ;
        RECT 58.600 15.290 59.680 15.590 ;
        RECT 54.800 14.710 55.720 14.750 ;
        RECT 58.760 14.710 59.680 14.750 ;
        RECT 54.040 14.410 55.720 14.710 ;
        RECT 58.600 14.410 60.460 14.710 ;
        RECT 54.040 14.270 54.340 14.410 ;
        RECT 50.320 13.970 54.340 14.270 ;
        RECT 13.600 13.020 49.240 13.460 ;
        RECT 50.320 13.020 51.400 13.970 ;
        RECT 54.040 13.830 54.340 13.970 ;
        RECT 60.160 14.270 60.460 14.410 ;
        RECT 62.920 14.270 64.000 28.050 ;
        RECT 77.320 31.870 78.400 32.820 ;
        RECT 81.640 32.310 82.560 32.350 ;
        RECT 85.600 32.310 86.520 32.350 ;
        RECT 80.860 32.010 82.720 32.310 ;
        RECT 85.600 32.010 87.280 32.310 ;
        RECT 80.860 31.870 81.160 32.010 ;
        RECT 77.320 31.570 81.160 31.870 ;
        RECT 77.320 28.350 78.400 31.570 ;
        RECT 80.860 31.430 81.160 31.570 ;
        RECT 86.980 31.870 87.280 32.010 ;
        RECT 89.920 31.870 91.000 32.820 ;
        RECT 86.980 31.570 91.000 31.870 ;
        RECT 81.640 31.430 82.560 31.470 ;
        RECT 85.600 31.430 86.520 31.470 ;
        RECT 86.980 31.430 87.280 31.570 ;
        RECT 80.860 31.130 82.720 31.430 ;
        RECT 85.600 31.130 87.280 31.430 ;
        RECT 81.640 30.550 82.560 30.590 ;
        RECT 81.640 30.250 82.720 30.550 ;
        RECT 85.600 30.250 87.280 30.550 ;
        RECT 86.980 30.110 87.280 30.250 ;
        RECT 79.480 29.810 80.560 30.110 ;
        RECT 86.980 29.810 88.840 30.110 ;
        RECT 81.640 29.670 82.560 29.710 ;
        RECT 85.600 29.670 86.520 29.710 ;
        RECT 81.640 29.370 82.720 29.670 ;
        RECT 85.600 29.370 86.680 29.670 ;
        RECT 81.640 28.790 82.560 28.830 ;
        RECT 85.600 28.790 86.520 28.830 ;
        RECT 80.860 28.490 82.720 28.790 ;
        RECT 85.600 28.490 87.280 28.790 ;
        RECT 80.860 28.350 81.160 28.490 ;
        RECT 77.320 28.050 81.160 28.350 ;
        RECT 65.800 26.730 67.480 27.030 ;
        RECT 65.800 26.150 66.720 26.190 ;
        RECT 65.200 25.850 66.880 26.150 ;
        RECT 65.200 24.390 65.500 25.850 ;
        RECT 67.180 25.270 67.480 26.730 ;
        RECT 68.120 26.590 69.040 26.630 ;
        RECT 67.960 26.290 69.040 26.590 ;
        RECT 65.800 24.970 67.480 25.270 ;
        RECT 65.200 24.090 66.880 24.390 ;
        RECT 65.200 22.630 65.500 24.090 ;
        RECT 67.180 23.510 67.480 24.970 ;
        RECT 68.350 24.830 68.650 26.290 ;
        RECT 67.960 24.530 69.040 24.830 ;
        RECT 65.800 23.210 67.480 23.510 ;
        RECT 65.200 22.330 66.880 22.630 ;
        RECT 65.200 20.870 65.500 22.330 ;
        RECT 67.180 21.750 67.480 23.210 ;
        RECT 68.350 23.070 68.650 24.530 ;
        RECT 67.960 22.770 69.040 23.070 ;
        RECT 65.800 21.450 67.480 21.750 ;
        RECT 65.200 20.570 66.880 20.870 ;
        RECT 67.180 19.990 67.480 21.450 ;
        RECT 68.350 21.310 68.650 22.770 ;
        RECT 67.960 21.010 69.040 21.310 ;
        RECT 65.800 19.690 67.480 19.990 ;
        RECT 65.800 19.110 66.720 19.150 ;
        RECT 60.160 13.970 64.000 14.270 ;
        RECT 54.800 13.830 55.720 13.870 ;
        RECT 58.760 13.830 59.680 13.870 ;
        RECT 60.160 13.830 60.460 13.970 ;
        RECT 54.040 13.530 55.720 13.830 ;
        RECT 58.600 13.530 60.460 13.830 ;
        RECT 62.920 13.020 64.000 13.970 ;
        RECT 65.200 18.810 66.880 19.110 ;
        RECT 65.200 17.350 65.500 18.810 ;
        RECT 65.960 18.230 66.880 18.270 ;
        RECT 67.180 18.230 67.480 19.690 ;
        RECT 67.960 19.250 69.040 19.550 ;
        RECT 65.800 17.930 67.480 18.230 ;
        RECT 65.200 17.050 66.880 17.350 ;
        RECT 65.200 15.590 65.500 17.050 ;
        RECT 67.180 16.470 67.480 17.930 ;
        RECT 68.350 17.830 68.650 19.250 ;
        RECT 68.040 17.790 68.960 17.830 ;
        RECT 67.960 17.490 69.040 17.790 ;
        RECT 65.800 16.170 67.480 16.470 ;
        RECT 65.200 15.290 66.880 15.590 ;
        RECT 65.200 13.830 65.500 15.290 ;
        RECT 67.180 14.710 67.480 16.170 ;
        RECT 68.350 16.030 68.650 17.490 ;
        RECT 67.960 15.730 69.040 16.030 ;
        RECT 65.800 14.410 67.480 14.710 ;
        RECT 65.880 14.370 66.800 14.410 ;
        RECT 68.350 14.270 68.650 15.730 ;
        RECT 67.960 13.970 69.040 14.270 ;
        RECT 65.200 13.530 66.880 13.830 ;
        RECT 70.120 13.020 71.200 27.540 ;
        RECT 73.840 26.730 75.520 27.030 ;
        RECT 72.280 26.590 73.200 26.630 ;
        RECT 72.280 26.290 73.360 26.590 ;
        RECT 72.670 24.830 72.970 26.290 ;
        RECT 73.840 25.270 74.140 26.730 ;
        RECT 74.440 26.150 75.360 26.190 ;
        RECT 74.440 25.850 76.120 26.150 ;
        RECT 73.840 24.970 75.520 25.270 ;
        RECT 72.280 24.530 73.360 24.830 ;
        RECT 72.670 23.070 72.970 24.530 ;
        RECT 73.840 23.510 74.140 24.970 ;
        RECT 75.820 24.390 76.120 25.850 ;
        RECT 74.440 24.090 76.120 24.390 ;
        RECT 73.840 23.210 75.520 23.510 ;
        RECT 72.280 22.770 73.360 23.070 ;
        RECT 72.670 21.310 72.970 22.770 ;
        RECT 73.840 21.750 74.140 23.210 ;
        RECT 75.820 22.630 76.120 24.090 ;
        RECT 74.440 22.330 76.120 22.630 ;
        RECT 73.840 21.450 75.520 21.750 ;
        RECT 72.280 21.010 73.360 21.310 ;
        RECT 73.840 19.990 74.140 21.450 ;
        RECT 75.820 20.870 76.120 22.330 ;
        RECT 74.440 20.570 76.120 20.870 ;
        RECT 73.840 19.690 75.520 19.990 ;
        RECT 72.280 19.250 73.360 19.550 ;
        RECT 72.670 17.830 72.970 19.250 ;
        RECT 73.840 18.230 74.140 19.690 ;
        RECT 74.440 19.110 75.360 19.150 ;
        RECT 74.440 18.810 76.120 19.110 ;
        RECT 74.440 18.230 75.360 18.270 ;
        RECT 73.840 17.930 75.520 18.230 ;
        RECT 72.360 17.790 73.280 17.830 ;
        RECT 72.280 17.490 73.360 17.790 ;
        RECT 72.670 16.030 72.970 17.490 ;
        RECT 73.840 16.470 74.140 17.930 ;
        RECT 75.820 17.350 76.120 18.810 ;
        RECT 74.440 17.050 76.120 17.350 ;
        RECT 73.840 16.170 75.520 16.470 ;
        RECT 72.280 15.730 73.360 16.030 ;
        RECT 72.670 14.270 72.970 15.730 ;
        RECT 73.840 14.710 74.140 16.170 ;
        RECT 75.820 15.590 76.120 17.050 ;
        RECT 74.440 15.290 76.120 15.590 ;
        RECT 73.840 14.410 75.520 14.710 ;
        RECT 74.520 14.370 75.440 14.410 ;
        RECT 72.280 13.970 73.360 14.270 ;
        RECT 75.820 13.830 76.120 15.290 ;
        RECT 74.440 13.530 76.120 13.830 ;
        RECT 77.320 14.270 78.400 28.050 ;
        RECT 80.860 27.910 81.160 28.050 ;
        RECT 86.980 28.350 87.280 28.490 ;
        RECT 89.920 28.350 91.000 31.570 ;
        RECT 92.080 31.940 92.440 33.260 ;
        RECT 92.800 32.380 127.720 32.820 ;
        RECT 92.080 31.500 127.000 31.940 ;
        RECT 92.080 30.180 92.440 31.500 ;
        RECT 127.360 31.060 127.720 32.380 ;
        RECT 92.800 30.620 127.720 31.060 ;
        RECT 92.080 29.740 127.000 30.180 ;
        RECT 127.360 29.300 127.720 30.620 ;
        RECT 92.080 28.860 127.720 29.300 ;
        RECT 86.980 28.050 91.000 28.350 ;
        RECT 81.640 27.910 82.560 27.950 ;
        RECT 85.600 27.910 86.520 27.950 ;
        RECT 86.980 27.910 87.280 28.050 ;
        RECT 80.860 27.610 82.720 27.910 ;
        RECT 85.600 27.610 87.280 27.910 ;
        RECT 85.600 27.030 86.520 27.240 ;
        RECT 80.860 26.730 82.720 27.030 ;
        RECT 85.600 26.730 86.680 27.030 ;
        RECT 80.860 26.590 81.160 26.730 ;
        RECT 79.480 26.290 81.160 26.590 ;
        RECT 87.760 26.290 88.840 26.590 ;
        RECT 81.640 26.150 82.560 26.190 ;
        RECT 85.600 26.150 86.520 26.190 ;
        RECT 81.640 25.850 82.720 26.150 ;
        RECT 85.600 25.850 86.680 26.150 ;
        RECT 81.720 25.270 82.640 25.310 ;
        RECT 85.600 25.270 86.520 25.310 ;
        RECT 81.640 24.970 83.320 25.270 ;
        RECT 85.600 24.970 86.680 25.270 ;
        RECT 79.480 24.830 80.400 24.870 ;
        RECT 79.480 24.530 80.560 24.830 ;
        RECT 81.640 24.090 82.720 24.390 ;
        RECT 82.030 23.510 82.330 24.090 ;
        RECT 81.640 23.210 82.720 23.510 ;
        RECT 79.480 23.070 80.400 23.110 ;
        RECT 79.480 22.770 80.560 23.070 ;
        RECT 81.640 22.630 82.560 22.670 ;
        RECT 83.020 22.630 83.320 24.970 ;
        RECT 86.980 24.530 88.840 24.830 ;
        RECT 85.600 24.090 86.680 24.390 ;
        RECT 85.990 23.550 86.290 24.090 ;
        RECT 85.600 23.510 86.520 23.550 ;
        RECT 85.600 23.210 86.680 23.510 ;
        RECT 86.980 22.630 87.280 24.530 ;
        RECT 87.760 22.770 88.840 23.070 ;
        RECT 81.640 22.330 82.720 22.630 ;
        RECT 83.020 22.330 87.280 22.630 ;
        RECT 81.640 21.750 82.560 21.790 ;
        RECT 81.640 21.450 86.680 21.750 ;
        RECT 79.480 21.010 81.160 21.310 ;
        RECT 87.760 21.010 89.440 21.310 ;
        RECT 79.480 19.250 80.560 19.550 ;
        RECT 79.870 17.790 80.170 19.250 ;
        RECT 79.480 17.490 80.560 17.790 ;
        RECT 80.860 17.350 81.160 21.010 ;
        RECT 85.600 20.870 86.520 20.910 ;
        RECT 81.640 20.570 86.680 20.870 ;
        RECT 82.030 19.990 82.330 20.570 ;
        RECT 85.990 19.990 86.290 20.570 ;
        RECT 81.640 19.690 82.720 19.990 ;
        RECT 85.600 19.690 86.680 19.990 ;
        RECT 87.760 19.550 88.680 19.590 ;
        RECT 87.760 19.250 88.840 19.550 ;
        RECT 81.640 19.110 82.560 19.150 ;
        RECT 85.600 19.110 86.520 19.150 ;
        RECT 81.640 18.810 82.720 19.110 ;
        RECT 85.600 18.810 86.680 19.110 ;
        RECT 82.030 18.270 82.330 18.810 ;
        RECT 85.990 18.270 86.290 18.810 ;
        RECT 81.640 18.230 82.560 18.270 ;
        RECT 85.600 18.230 86.520 18.270 ;
        RECT 81.640 17.930 82.720 18.230 ;
        RECT 85.600 17.930 86.680 18.230 ;
        RECT 87.760 17.790 88.680 17.830 ;
        RECT 89.140 17.790 89.440 21.010 ;
        RECT 87.760 17.490 89.440 17.790 ;
        RECT 80.860 17.050 86.680 17.350 ;
        RECT 81.640 16.470 82.560 16.700 ;
        RECT 85.600 16.470 86.520 16.510 ;
        RECT 81.640 16.170 86.680 16.470 ;
        RECT 79.560 16.030 80.480 16.070 ;
        RECT 79.480 15.730 80.560 16.030 ;
        RECT 87.760 15.730 88.840 16.030 ;
        RECT 81.640 15.590 82.560 15.630 ;
        RECT 85.600 15.590 86.520 15.630 ;
        RECT 81.640 15.290 82.720 15.590 ;
        RECT 85.600 15.290 86.680 15.590 ;
        RECT 81.640 14.710 82.560 14.750 ;
        RECT 85.600 14.710 86.520 14.750 ;
        RECT 80.860 14.410 82.720 14.710 ;
        RECT 85.600 14.410 87.280 14.710 ;
        RECT 80.860 14.270 81.160 14.410 ;
        RECT 77.320 13.970 81.160 14.270 ;
        RECT 77.320 13.020 78.400 13.970 ;
        RECT 80.860 13.830 81.160 13.970 ;
        RECT 86.980 14.270 87.280 14.410 ;
        RECT 89.920 14.270 91.000 28.050 ;
        RECT 92.080 27.980 127.720 28.420 ;
        RECT 92.080 26.660 92.440 27.980 ;
        RECT 92.800 27.100 127.720 27.540 ;
        RECT 92.080 26.220 127.000 26.660 ;
        RECT 92.080 24.900 92.440 26.220 ;
        RECT 127.360 25.780 127.720 27.100 ;
        RECT 92.800 25.340 127.720 25.780 ;
        RECT 92.080 24.460 127.000 24.900 ;
        RECT 127.360 24.020 127.720 25.340 ;
        RECT 92.080 23.580 127.720 24.020 ;
        RECT 92.080 22.700 127.720 23.140 ;
        RECT 92.080 21.380 92.440 22.700 ;
        RECT 92.800 21.820 127.720 22.260 ;
        RECT 92.080 20.940 127.000 21.380 ;
        RECT 92.080 19.620 92.440 20.940 ;
        RECT 127.360 20.500 127.720 21.820 ;
        RECT 92.800 20.060 127.720 20.500 ;
        RECT 92.080 19.180 127.000 19.620 ;
        RECT 127.360 18.740 127.720 20.060 ;
        RECT 92.080 18.300 127.720 18.740 ;
        RECT 86.980 13.970 91.000 14.270 ;
        RECT 81.640 13.830 82.560 13.870 ;
        RECT 85.600 13.830 86.520 13.870 ;
        RECT 86.980 13.830 87.280 13.970 ;
        RECT 80.860 13.530 82.720 13.830 ;
        RECT 85.600 13.530 87.280 13.830 ;
        RECT 89.920 13.020 91.000 13.970 ;
        RECT 92.080 17.420 127.720 17.860 ;
        RECT 92.080 16.100 92.440 17.420 ;
        RECT 92.800 16.540 127.720 16.980 ;
        RECT 92.080 15.660 127.000 16.100 ;
        RECT 92.080 14.340 92.440 15.660 ;
        RECT 127.360 15.220 127.720 16.540 ;
        RECT 92.800 14.780 127.720 15.220 ;
        RECT 92.080 13.900 127.000 14.340 ;
        RECT 127.360 13.460 127.720 14.780 ;
        RECT 92.080 13.020 127.720 13.460 ;
        RECT 130.920 10.640 131.920 213.990 ;
        RECT 8.640 9.640 131.920 10.640 ;
        RECT 134.520 7.040 135.520 217.590 ;
        RECT 5.040 6.040 135.520 7.040 ;
        RECT 60.840 5.320 61.760 5.360 ;
        RECT 79.560 5.320 80.480 5.360 ;
        RECT 136.240 5.320 136.540 222.190 ;
        RECT 5.040 5.020 136.540 5.320 ;
        RECT 139.360 221.930 140.440 222.880 ;
        RECT 143.680 222.370 144.600 222.410 ;
        RECT 147.640 222.370 148.560 222.410 ;
        RECT 142.900 222.070 144.760 222.370 ;
        RECT 147.640 222.070 149.320 222.370 ;
        RECT 142.900 221.930 143.200 222.070 ;
        RECT 139.360 221.630 143.200 221.930 ;
        RECT 61.600 4.300 62.520 4.340 ;
        RECT 78.720 4.300 79.640 4.340 ;
        RECT 4.020 4.000 136.540 4.300 ;
        RECT 139.360 3.690 140.440 221.630 ;
        RECT 142.900 221.490 143.200 221.630 ;
        RECT 149.020 221.930 149.320 222.070 ;
        RECT 151.960 221.930 153.040 222.880 ;
        RECT 149.020 221.630 153.040 221.930 ;
        RECT 143.680 221.490 144.600 221.530 ;
        RECT 147.640 221.490 148.560 221.530 ;
        RECT 149.020 221.490 149.320 221.630 ;
        RECT 142.900 221.190 144.760 221.490 ;
        RECT 147.640 221.190 149.320 221.490 ;
        RECT 147.640 220.610 148.560 220.650 ;
        RECT 143.680 220.310 148.720 220.610 ;
        RECT 141.520 219.870 143.200 220.170 ;
        RECT 149.800 219.870 150.880 220.170 ;
        RECT 142.900 218.850 143.200 219.870 ;
        RECT 143.680 219.730 144.600 219.770 ;
        RECT 147.640 219.730 148.560 219.770 ;
        RECT 143.680 219.430 144.760 219.730 ;
        RECT 147.640 219.430 148.720 219.730 ;
        RECT 143.680 218.850 144.600 218.890 ;
        RECT 142.900 218.550 148.720 218.850 ;
        RECT 141.520 218.410 142.440 218.450 ;
        RECT 141.520 218.110 142.600 218.410 ;
        RECT 149.020 218.110 150.880 218.410 ;
        RECT 143.680 217.670 144.760 217.970 ;
        RECT 147.640 217.670 148.720 217.970 ;
        RECT 144.070 217.090 144.370 217.670 ;
        RECT 148.030 217.090 148.330 217.670 ;
        RECT 143.680 216.790 148.720 217.090 ;
        RECT 141.520 216.350 142.600 216.650 ;
        RECT 143.680 215.910 144.760 216.210 ;
        RECT 144.070 215.330 144.370 215.910 ;
        RECT 143.680 215.030 144.760 215.330 ;
        RECT 141.520 214.890 142.440 214.930 ;
        RECT 141.520 214.590 142.600 214.890 ;
        RECT 143.680 214.450 144.600 214.490 ;
        RECT 147.040 214.450 147.340 216.790 ;
        RECT 147.640 216.210 148.560 216.250 ;
        RECT 147.640 215.910 148.720 216.210 ;
        RECT 147.640 215.330 148.560 215.370 ;
        RECT 147.640 215.030 148.720 215.330 ;
        RECT 143.680 214.150 144.760 214.450 ;
        RECT 147.040 214.150 148.720 214.450 ;
        RECT 143.680 213.570 144.600 213.610 ;
        RECT 143.680 213.270 148.720 213.570 ;
        RECT 141.520 212.830 142.600 213.130 ;
        RECT 142.300 212.530 143.200 212.830 ;
        RECT 141.520 211.070 142.600 211.370 ;
        RECT 141.520 209.610 142.440 209.650 ;
        RECT 141.520 209.310 142.600 209.610 ;
        RECT 142.900 207.850 143.200 212.530 ;
        RECT 143.680 212.390 144.760 212.690 ;
        RECT 147.640 212.390 148.720 212.690 ;
        RECT 144.070 211.810 144.370 212.390 ;
        RECT 148.030 211.810 148.330 212.390 ;
        RECT 143.680 211.510 144.760 211.810 ;
        RECT 147.640 211.510 148.720 211.810 ;
        RECT 143.680 210.930 144.600 210.970 ;
        RECT 147.640 210.930 148.560 210.970 ;
        RECT 143.680 210.630 144.760 210.930 ;
        RECT 147.640 210.630 148.720 210.930 ;
        RECT 147.640 210.050 148.560 210.090 ;
        RECT 143.680 209.750 148.720 210.050 ;
        RECT 143.680 209.170 144.600 209.210 ;
        RECT 147.640 209.170 148.560 209.210 ;
        RECT 143.680 208.870 144.760 209.170 ;
        RECT 147.640 208.870 148.720 209.170 ;
        RECT 143.680 208.290 144.600 208.330 ;
        RECT 143.680 207.990 148.720 208.290 ;
        RECT 141.520 207.550 143.200 207.850 ;
        RECT 141.520 205.790 142.600 206.090 ;
        RECT 141.520 204.330 142.440 204.370 ;
        RECT 141.520 204.030 142.600 204.330 ;
        RECT 141.520 202.270 142.600 202.570 ;
        RECT 142.900 201.250 143.200 207.550 ;
        RECT 143.680 207.110 144.760 207.410 ;
        RECT 144.070 206.530 144.370 207.110 ;
        RECT 143.680 206.230 144.760 206.530 ;
        RECT 143.680 205.650 144.600 205.690 ;
        RECT 143.680 205.350 144.760 205.650 ;
        RECT 145.060 204.770 145.360 207.990 ;
        RECT 147.640 207.110 148.720 207.410 ;
        RECT 148.030 206.530 148.330 207.110 ;
        RECT 147.640 206.230 148.720 206.530 ;
        RECT 147.640 205.650 148.560 205.690 ;
        RECT 147.640 205.350 148.720 205.650 ;
        RECT 143.680 204.470 148.720 204.770 ;
        RECT 149.020 204.330 149.320 218.110 ;
        RECT 149.800 216.650 150.720 216.690 ;
        RECT 149.800 216.350 150.880 216.650 ;
        RECT 149.800 214.590 150.880 214.890 ;
        RECT 149.800 213.130 150.720 213.170 ;
        RECT 149.800 212.830 150.880 213.130 ;
        RECT 149.800 211.370 150.720 211.410 ;
        RECT 149.800 211.070 150.880 211.370 ;
        RECT 149.800 209.310 150.880 209.610 ;
        RECT 149.800 207.850 150.720 207.890 ;
        RECT 149.800 207.550 150.880 207.850 ;
        RECT 149.800 206.090 150.720 206.130 ;
        RECT 149.800 205.790 150.880 206.090 ;
        RECT 149.020 204.030 150.880 204.330 ;
        RECT 143.680 203.590 144.760 203.890 ;
        RECT 147.640 203.590 148.720 203.890 ;
        RECT 144.070 203.010 144.370 203.590 ;
        RECT 148.030 203.010 148.330 203.590 ;
        RECT 143.680 202.710 144.760 203.010 ;
        RECT 147.640 202.710 148.720 203.010 ;
        RECT 143.680 202.130 144.600 202.170 ;
        RECT 147.640 202.130 148.560 202.170 ;
        RECT 143.680 201.830 144.760 202.130 ;
        RECT 147.640 201.830 148.720 202.130 ;
        RECT 149.020 201.250 149.320 204.030 ;
        RECT 149.800 202.270 150.880 202.570 ;
        RECT 142.900 200.950 149.320 201.250 ;
        RECT 141.520 200.510 142.600 200.810 ;
        RECT 149.800 200.510 150.880 200.810 ;
        RECT 143.680 200.370 144.600 200.410 ;
        RECT 147.640 200.370 148.560 200.410 ;
        RECT 143.680 200.070 144.760 200.370 ;
        RECT 147.640 200.070 148.720 200.370 ;
        RECT 149.020 200.210 150.100 200.510 ;
        RECT 143.680 199.490 144.600 199.530 ;
        RECT 147.640 199.490 148.560 199.530 ;
        RECT 143.680 199.190 145.360 199.490 ;
        RECT 147.640 199.190 148.720 199.490 ;
        RECT 141.520 199.050 142.440 199.090 ;
        RECT 141.520 198.750 142.600 199.050 ;
        RECT 145.060 198.610 145.360 199.190 ;
        RECT 143.680 198.310 144.760 198.610 ;
        RECT 145.060 198.310 148.720 198.610 ;
        RECT 144.070 197.730 144.370 198.310 ;
        RECT 145.060 197.730 145.360 198.310 ;
        RECT 147.640 197.730 148.560 197.770 ;
        RECT 149.020 197.730 149.320 200.210 ;
        RECT 149.800 198.750 150.880 199.050 ;
        RECT 143.680 197.430 144.760 197.730 ;
        RECT 145.060 197.430 149.320 197.730 ;
        RECT 141.520 196.990 142.600 197.290 ;
        RECT 149.800 196.990 150.880 197.290 ;
        RECT 143.680 196.850 144.600 196.890 ;
        RECT 147.640 196.850 148.560 196.890 ;
        RECT 143.680 196.550 144.760 196.850 ;
        RECT 147.640 196.550 148.720 196.850 ;
        RECT 147.640 195.970 148.560 196.010 ;
        RECT 143.680 195.670 148.720 195.970 ;
        RECT 141.520 195.230 143.200 195.530 ;
        RECT 149.800 195.230 150.880 195.530 ;
        RECT 142.900 194.210 143.200 195.230 ;
        RECT 143.680 195.090 144.600 195.130 ;
        RECT 147.640 195.090 148.560 195.130 ;
        RECT 143.680 194.790 144.760 195.090 ;
        RECT 147.640 194.790 148.720 195.090 ;
        RECT 143.680 194.210 144.600 194.250 ;
        RECT 142.900 193.910 148.720 194.210 ;
        RECT 141.520 193.770 142.440 193.810 ;
        RECT 141.520 193.470 142.600 193.770 ;
        RECT 149.020 193.470 150.880 193.770 ;
        RECT 143.680 193.030 144.760 193.330 ;
        RECT 147.640 193.030 148.720 193.330 ;
        RECT 144.070 192.450 144.370 193.030 ;
        RECT 148.030 192.450 148.330 193.030 ;
        RECT 143.680 192.150 148.720 192.450 ;
        RECT 141.520 191.710 142.600 192.010 ;
        RECT 143.680 191.270 144.760 191.570 ;
        RECT 144.070 190.690 144.370 191.270 ;
        RECT 143.680 190.390 144.760 190.690 ;
        RECT 141.520 190.250 142.440 190.290 ;
        RECT 141.520 189.950 142.600 190.250 ;
        RECT 143.680 189.810 144.600 189.850 ;
        RECT 147.040 189.810 147.340 192.150 ;
        RECT 147.640 191.570 148.560 191.610 ;
        RECT 147.640 191.270 148.720 191.570 ;
        RECT 147.640 190.690 148.560 190.730 ;
        RECT 147.640 190.390 148.720 190.690 ;
        RECT 143.680 189.510 144.760 189.810 ;
        RECT 147.040 189.510 148.720 189.810 ;
        RECT 143.680 188.930 144.600 188.970 ;
        RECT 143.680 188.630 148.720 188.930 ;
        RECT 141.520 188.190 142.600 188.490 ;
        RECT 142.300 187.890 143.200 188.190 ;
        RECT 141.520 186.430 142.600 186.730 ;
        RECT 141.520 184.970 142.440 185.010 ;
        RECT 141.520 184.670 142.600 184.970 ;
        RECT 142.900 183.210 143.200 187.890 ;
        RECT 143.680 187.750 144.760 188.050 ;
        RECT 147.640 187.750 148.720 188.050 ;
        RECT 144.070 187.170 144.370 187.750 ;
        RECT 148.030 187.170 148.330 187.750 ;
        RECT 143.680 186.870 144.760 187.170 ;
        RECT 147.640 186.870 148.720 187.170 ;
        RECT 143.680 186.290 144.600 186.330 ;
        RECT 147.640 186.290 148.560 186.330 ;
        RECT 143.680 185.990 144.760 186.290 ;
        RECT 147.640 185.990 148.720 186.290 ;
        RECT 147.640 185.410 148.560 185.450 ;
        RECT 143.680 185.110 148.720 185.410 ;
        RECT 143.680 184.530 144.600 184.570 ;
        RECT 147.640 184.530 148.560 184.570 ;
        RECT 143.680 184.230 144.760 184.530 ;
        RECT 147.640 184.230 148.720 184.530 ;
        RECT 143.680 183.650 144.600 183.690 ;
        RECT 143.680 183.350 148.720 183.650 ;
        RECT 141.520 182.910 143.200 183.210 ;
        RECT 141.520 181.150 142.600 181.450 ;
        RECT 141.520 179.690 142.440 179.730 ;
        RECT 141.520 179.390 142.600 179.690 ;
        RECT 141.520 177.630 142.600 177.930 ;
        RECT 142.900 176.610 143.200 182.910 ;
        RECT 143.680 182.470 144.760 182.770 ;
        RECT 144.070 181.890 144.370 182.470 ;
        RECT 143.680 181.590 144.760 181.890 ;
        RECT 143.680 181.010 144.600 181.050 ;
        RECT 143.680 180.710 144.760 181.010 ;
        RECT 145.060 180.130 145.360 183.350 ;
        RECT 147.640 182.470 148.720 182.770 ;
        RECT 148.030 181.890 148.330 182.470 ;
        RECT 147.640 181.590 148.720 181.890 ;
        RECT 147.640 181.010 148.560 181.050 ;
        RECT 147.640 180.710 148.720 181.010 ;
        RECT 143.680 179.830 148.720 180.130 ;
        RECT 149.020 179.690 149.320 193.470 ;
        RECT 149.800 192.010 150.720 192.050 ;
        RECT 149.800 191.710 150.880 192.010 ;
        RECT 149.800 189.950 150.880 190.250 ;
        RECT 149.800 188.490 150.720 188.530 ;
        RECT 149.800 188.190 150.880 188.490 ;
        RECT 149.800 186.730 150.720 186.770 ;
        RECT 149.800 186.430 150.880 186.730 ;
        RECT 149.800 184.670 150.880 184.970 ;
        RECT 149.800 183.210 150.720 183.250 ;
        RECT 149.800 182.910 150.880 183.210 ;
        RECT 149.800 181.450 150.720 181.490 ;
        RECT 149.800 181.150 150.880 181.450 ;
        RECT 149.020 179.390 150.880 179.690 ;
        RECT 143.680 178.950 144.760 179.250 ;
        RECT 147.640 178.950 148.720 179.250 ;
        RECT 144.070 178.370 144.370 178.950 ;
        RECT 148.030 178.370 148.330 178.950 ;
        RECT 143.680 178.070 144.760 178.370 ;
        RECT 147.640 178.070 148.720 178.370 ;
        RECT 143.680 177.490 144.600 177.530 ;
        RECT 147.640 177.490 148.560 177.530 ;
        RECT 143.680 177.190 144.760 177.490 ;
        RECT 147.640 177.190 148.720 177.490 ;
        RECT 149.020 176.610 149.320 179.390 ;
        RECT 149.800 177.630 150.880 177.930 ;
        RECT 142.900 176.310 149.320 176.610 ;
        RECT 141.520 175.870 142.600 176.170 ;
        RECT 149.800 175.870 150.880 176.170 ;
        RECT 143.680 175.730 144.600 175.770 ;
        RECT 147.640 175.730 148.560 175.770 ;
        RECT 143.680 175.430 144.760 175.730 ;
        RECT 147.640 175.430 148.720 175.730 ;
        RECT 149.020 175.570 150.100 175.870 ;
        RECT 143.680 174.850 144.600 174.890 ;
        RECT 147.640 174.850 148.560 174.890 ;
        RECT 143.680 174.550 145.360 174.850 ;
        RECT 147.640 174.550 148.720 174.850 ;
        RECT 141.520 174.410 142.440 174.450 ;
        RECT 141.520 174.110 142.600 174.410 ;
        RECT 145.060 173.970 145.360 174.550 ;
        RECT 143.680 173.670 144.760 173.970 ;
        RECT 145.060 173.670 148.720 173.970 ;
        RECT 144.070 173.090 144.370 173.670 ;
        RECT 145.060 173.090 145.360 173.670 ;
        RECT 147.640 173.090 148.560 173.130 ;
        RECT 149.020 173.090 149.320 175.570 ;
        RECT 149.800 174.110 150.880 174.410 ;
        RECT 143.680 172.790 144.760 173.090 ;
        RECT 145.060 172.790 149.320 173.090 ;
        RECT 141.520 172.350 142.600 172.650 ;
        RECT 149.800 172.350 150.880 172.650 ;
        RECT 143.680 172.210 144.600 172.250 ;
        RECT 147.640 172.210 148.560 172.250 ;
        RECT 143.680 171.910 144.760 172.210 ;
        RECT 147.640 171.910 148.720 172.210 ;
        RECT 147.640 171.330 148.560 171.370 ;
        RECT 143.680 171.030 148.720 171.330 ;
        RECT 141.520 170.590 143.200 170.890 ;
        RECT 149.800 170.590 150.880 170.890 ;
        RECT 142.900 169.570 143.200 170.590 ;
        RECT 143.680 170.450 144.600 170.490 ;
        RECT 147.640 170.450 148.560 170.490 ;
        RECT 143.680 170.150 144.760 170.450 ;
        RECT 147.640 170.150 148.720 170.450 ;
        RECT 143.680 169.570 144.600 169.610 ;
        RECT 142.900 169.270 148.720 169.570 ;
        RECT 141.520 169.130 142.440 169.170 ;
        RECT 141.520 168.830 142.600 169.130 ;
        RECT 149.020 168.830 150.880 169.130 ;
        RECT 143.680 168.390 144.760 168.690 ;
        RECT 147.640 168.390 148.720 168.690 ;
        RECT 144.070 167.810 144.370 168.390 ;
        RECT 148.030 167.810 148.330 168.390 ;
        RECT 143.680 167.510 148.720 167.810 ;
        RECT 141.520 167.070 142.600 167.370 ;
        RECT 143.680 166.630 144.760 166.930 ;
        RECT 144.070 166.050 144.370 166.630 ;
        RECT 143.680 165.750 144.760 166.050 ;
        RECT 141.520 165.610 142.440 165.650 ;
        RECT 141.520 165.310 142.600 165.610 ;
        RECT 143.680 165.170 144.600 165.210 ;
        RECT 147.040 165.170 147.340 167.510 ;
        RECT 147.640 166.930 148.560 166.970 ;
        RECT 147.640 166.630 148.720 166.930 ;
        RECT 147.640 166.050 148.560 166.090 ;
        RECT 147.640 165.750 148.720 166.050 ;
        RECT 143.680 164.870 144.760 165.170 ;
        RECT 147.040 164.870 148.720 165.170 ;
        RECT 143.680 164.290 144.600 164.330 ;
        RECT 143.680 163.990 148.720 164.290 ;
        RECT 141.520 163.550 142.600 163.850 ;
        RECT 142.300 163.250 143.200 163.550 ;
        RECT 141.520 161.790 142.600 162.090 ;
        RECT 141.520 160.330 142.440 160.370 ;
        RECT 141.520 160.030 142.600 160.330 ;
        RECT 142.900 158.570 143.200 163.250 ;
        RECT 143.680 163.110 144.760 163.410 ;
        RECT 147.640 163.110 148.720 163.410 ;
        RECT 144.070 162.530 144.370 163.110 ;
        RECT 148.030 162.530 148.330 163.110 ;
        RECT 143.680 162.230 144.760 162.530 ;
        RECT 147.640 162.230 148.720 162.530 ;
        RECT 143.680 161.650 144.600 161.690 ;
        RECT 147.640 161.650 148.560 161.690 ;
        RECT 143.680 161.350 144.760 161.650 ;
        RECT 147.640 161.350 148.720 161.650 ;
        RECT 147.640 160.770 148.560 160.810 ;
        RECT 143.680 160.470 148.720 160.770 ;
        RECT 143.680 159.890 144.600 159.930 ;
        RECT 147.640 159.890 148.560 159.930 ;
        RECT 143.680 159.590 144.760 159.890 ;
        RECT 147.640 159.590 148.720 159.890 ;
        RECT 143.680 159.010 144.600 159.050 ;
        RECT 143.680 158.710 148.720 159.010 ;
        RECT 141.520 158.270 143.200 158.570 ;
        RECT 141.520 156.510 142.600 156.810 ;
        RECT 141.520 155.050 142.440 155.090 ;
        RECT 141.520 154.750 142.600 155.050 ;
        RECT 141.520 152.990 142.600 153.290 ;
        RECT 142.900 151.970 143.200 158.270 ;
        RECT 143.680 157.830 144.760 158.130 ;
        RECT 144.070 157.250 144.370 157.830 ;
        RECT 143.680 156.950 144.760 157.250 ;
        RECT 143.680 156.370 144.600 156.410 ;
        RECT 143.680 156.070 144.760 156.370 ;
        RECT 145.060 155.490 145.360 158.710 ;
        RECT 147.640 157.830 148.720 158.130 ;
        RECT 148.030 157.250 148.330 157.830 ;
        RECT 147.640 156.950 148.720 157.250 ;
        RECT 147.640 156.370 148.560 156.410 ;
        RECT 147.640 156.070 148.720 156.370 ;
        RECT 143.680 155.190 148.720 155.490 ;
        RECT 149.020 155.050 149.320 168.830 ;
        RECT 149.800 167.370 150.720 167.410 ;
        RECT 149.800 167.070 150.880 167.370 ;
        RECT 149.800 165.310 150.880 165.610 ;
        RECT 149.800 163.850 150.720 163.890 ;
        RECT 149.800 163.550 150.880 163.850 ;
        RECT 149.800 162.090 150.720 162.130 ;
        RECT 149.800 161.790 150.880 162.090 ;
        RECT 149.800 160.030 150.880 160.330 ;
        RECT 149.800 158.570 150.720 158.610 ;
        RECT 149.800 158.270 150.880 158.570 ;
        RECT 149.800 156.810 150.720 156.850 ;
        RECT 149.800 156.510 150.880 156.810 ;
        RECT 149.020 154.750 150.880 155.050 ;
        RECT 143.680 154.310 144.760 154.610 ;
        RECT 147.640 154.310 148.720 154.610 ;
        RECT 144.070 153.730 144.370 154.310 ;
        RECT 148.030 153.730 148.330 154.310 ;
        RECT 143.680 153.430 144.760 153.730 ;
        RECT 147.640 153.430 148.720 153.730 ;
        RECT 143.680 152.850 144.600 152.890 ;
        RECT 147.640 152.850 148.560 152.890 ;
        RECT 143.680 152.550 144.760 152.850 ;
        RECT 147.640 152.550 148.720 152.850 ;
        RECT 149.020 151.970 149.320 154.750 ;
        RECT 149.800 152.990 150.880 153.290 ;
        RECT 142.900 151.670 149.320 151.970 ;
        RECT 141.520 151.230 142.600 151.530 ;
        RECT 149.800 151.230 150.880 151.530 ;
        RECT 143.680 151.090 144.600 151.130 ;
        RECT 147.640 151.090 148.560 151.130 ;
        RECT 143.680 150.790 144.760 151.090 ;
        RECT 147.640 150.790 148.720 151.090 ;
        RECT 149.020 150.930 150.100 151.230 ;
        RECT 143.680 150.210 144.600 150.250 ;
        RECT 147.640 150.210 148.560 150.250 ;
        RECT 143.680 149.910 145.360 150.210 ;
        RECT 147.640 149.910 148.720 150.210 ;
        RECT 141.520 149.770 142.440 149.810 ;
        RECT 141.520 149.470 142.600 149.770 ;
        RECT 145.060 149.330 145.360 149.910 ;
        RECT 143.680 149.030 144.760 149.330 ;
        RECT 145.060 149.030 148.720 149.330 ;
        RECT 144.070 148.450 144.370 149.030 ;
        RECT 145.060 148.450 145.360 149.030 ;
        RECT 147.640 148.450 148.560 148.490 ;
        RECT 149.020 148.450 149.320 150.930 ;
        RECT 149.800 149.470 150.880 149.770 ;
        RECT 143.680 148.150 144.760 148.450 ;
        RECT 145.060 148.150 149.320 148.450 ;
        RECT 141.520 147.710 142.600 148.010 ;
        RECT 149.800 147.710 150.880 148.010 ;
        RECT 143.680 147.570 144.600 147.610 ;
        RECT 147.640 147.570 148.560 147.610 ;
        RECT 143.680 147.270 144.760 147.570 ;
        RECT 147.640 147.270 148.720 147.570 ;
        RECT 147.640 146.690 148.560 146.730 ;
        RECT 143.680 146.390 148.720 146.690 ;
        RECT 141.520 145.950 143.200 146.250 ;
        RECT 149.800 145.950 150.880 146.250 ;
        RECT 142.900 144.930 143.200 145.950 ;
        RECT 143.680 145.810 144.600 145.850 ;
        RECT 147.640 145.810 148.560 145.850 ;
        RECT 143.680 145.510 144.760 145.810 ;
        RECT 147.640 145.510 148.720 145.810 ;
        RECT 143.680 144.930 144.600 144.970 ;
        RECT 142.900 144.630 148.720 144.930 ;
        RECT 141.520 144.490 142.440 144.530 ;
        RECT 141.520 144.190 142.600 144.490 ;
        RECT 149.020 144.190 150.880 144.490 ;
        RECT 143.680 143.750 144.760 144.050 ;
        RECT 147.640 143.750 148.720 144.050 ;
        RECT 144.070 143.170 144.370 143.750 ;
        RECT 148.030 143.170 148.330 143.750 ;
        RECT 143.680 142.870 148.720 143.170 ;
        RECT 141.520 142.430 142.600 142.730 ;
        RECT 143.680 141.990 144.760 142.290 ;
        RECT 144.070 141.410 144.370 141.990 ;
        RECT 143.680 141.110 144.760 141.410 ;
        RECT 141.520 140.970 142.440 141.010 ;
        RECT 141.520 140.670 142.600 140.970 ;
        RECT 143.680 140.530 144.600 140.570 ;
        RECT 147.040 140.530 147.340 142.870 ;
        RECT 147.640 142.290 148.560 142.330 ;
        RECT 147.640 141.990 148.720 142.290 ;
        RECT 147.640 141.410 148.560 141.450 ;
        RECT 147.640 141.110 148.720 141.410 ;
        RECT 143.680 140.230 144.760 140.530 ;
        RECT 147.040 140.230 148.720 140.530 ;
        RECT 143.680 139.650 144.600 139.690 ;
        RECT 143.680 139.350 148.720 139.650 ;
        RECT 141.520 138.910 142.600 139.210 ;
        RECT 142.300 138.610 143.200 138.910 ;
        RECT 141.520 137.150 142.600 137.450 ;
        RECT 141.520 135.690 142.440 135.730 ;
        RECT 141.520 135.390 142.600 135.690 ;
        RECT 142.900 133.930 143.200 138.610 ;
        RECT 143.680 138.470 144.760 138.770 ;
        RECT 147.640 138.470 148.720 138.770 ;
        RECT 144.070 137.890 144.370 138.470 ;
        RECT 148.030 137.890 148.330 138.470 ;
        RECT 143.680 137.590 144.760 137.890 ;
        RECT 147.640 137.590 148.720 137.890 ;
        RECT 143.680 137.010 144.600 137.050 ;
        RECT 147.640 137.010 148.560 137.050 ;
        RECT 143.680 136.710 144.760 137.010 ;
        RECT 147.640 136.710 148.720 137.010 ;
        RECT 147.640 136.130 148.560 136.170 ;
        RECT 143.680 135.830 148.720 136.130 ;
        RECT 143.680 135.250 144.600 135.290 ;
        RECT 147.640 135.250 148.560 135.290 ;
        RECT 143.680 134.950 144.760 135.250 ;
        RECT 147.640 134.950 148.720 135.250 ;
        RECT 143.680 134.370 144.600 134.410 ;
        RECT 143.680 134.070 148.720 134.370 ;
        RECT 141.520 133.630 143.200 133.930 ;
        RECT 141.520 131.870 142.600 132.170 ;
        RECT 141.520 130.410 142.440 130.450 ;
        RECT 141.520 130.110 142.600 130.410 ;
        RECT 141.520 128.350 142.600 128.650 ;
        RECT 142.900 127.330 143.200 133.630 ;
        RECT 143.680 133.190 144.760 133.490 ;
        RECT 144.070 132.610 144.370 133.190 ;
        RECT 143.680 132.310 144.760 132.610 ;
        RECT 143.680 131.730 144.600 131.770 ;
        RECT 143.680 131.430 144.760 131.730 ;
        RECT 145.060 130.850 145.360 134.070 ;
        RECT 147.640 133.190 148.720 133.490 ;
        RECT 148.030 132.610 148.330 133.190 ;
        RECT 147.640 132.310 148.720 132.610 ;
        RECT 147.640 131.730 148.560 131.770 ;
        RECT 147.640 131.430 148.720 131.730 ;
        RECT 143.680 130.550 148.720 130.850 ;
        RECT 149.020 130.410 149.320 144.190 ;
        RECT 149.800 142.730 150.720 142.770 ;
        RECT 149.800 142.430 150.880 142.730 ;
        RECT 149.800 140.670 150.880 140.970 ;
        RECT 149.800 139.210 150.720 139.250 ;
        RECT 149.800 138.910 150.880 139.210 ;
        RECT 149.800 137.450 150.720 137.490 ;
        RECT 149.800 137.150 150.880 137.450 ;
        RECT 149.800 135.390 150.880 135.690 ;
        RECT 149.800 133.930 150.720 133.970 ;
        RECT 149.800 133.630 150.880 133.930 ;
        RECT 149.800 132.170 150.720 132.210 ;
        RECT 149.800 131.870 150.880 132.170 ;
        RECT 149.020 130.110 150.880 130.410 ;
        RECT 143.680 129.670 144.760 129.970 ;
        RECT 147.640 129.670 148.720 129.970 ;
        RECT 144.070 129.090 144.370 129.670 ;
        RECT 148.030 129.090 148.330 129.670 ;
        RECT 143.680 128.790 144.760 129.090 ;
        RECT 147.640 128.790 148.720 129.090 ;
        RECT 143.680 128.210 144.600 128.250 ;
        RECT 147.640 128.210 148.560 128.250 ;
        RECT 143.680 127.910 144.760 128.210 ;
        RECT 147.640 127.910 148.720 128.210 ;
        RECT 149.020 127.330 149.320 130.110 ;
        RECT 149.800 128.350 150.880 128.650 ;
        RECT 142.900 127.030 149.320 127.330 ;
        RECT 141.520 126.590 142.600 126.890 ;
        RECT 149.800 126.590 150.880 126.890 ;
        RECT 143.680 126.450 144.600 126.490 ;
        RECT 147.640 126.450 148.560 126.490 ;
        RECT 143.680 126.150 144.760 126.450 ;
        RECT 147.640 126.150 148.720 126.450 ;
        RECT 149.020 126.290 150.100 126.590 ;
        RECT 143.680 125.570 144.600 125.610 ;
        RECT 147.640 125.570 148.560 125.610 ;
        RECT 143.680 125.270 145.360 125.570 ;
        RECT 147.640 125.270 148.720 125.570 ;
        RECT 141.520 125.130 142.440 125.170 ;
        RECT 141.520 124.830 142.600 125.130 ;
        RECT 145.060 124.690 145.360 125.270 ;
        RECT 143.680 124.390 144.760 124.690 ;
        RECT 145.060 124.390 148.720 124.690 ;
        RECT 144.070 123.810 144.370 124.390 ;
        RECT 145.060 123.810 145.360 124.390 ;
        RECT 147.640 123.810 148.560 123.850 ;
        RECT 149.020 123.810 149.320 126.290 ;
        RECT 149.800 124.830 150.880 125.130 ;
        RECT 143.680 123.510 144.760 123.810 ;
        RECT 145.060 123.510 149.320 123.810 ;
        RECT 141.520 123.070 142.600 123.370 ;
        RECT 149.800 123.070 150.880 123.370 ;
        RECT 143.680 122.930 144.600 122.970 ;
        RECT 147.640 122.930 148.560 122.970 ;
        RECT 143.680 122.630 144.760 122.930 ;
        RECT 147.640 122.630 148.720 122.930 ;
        RECT 147.640 122.050 148.560 122.090 ;
        RECT 143.680 121.750 148.720 122.050 ;
        RECT 141.520 121.310 143.200 121.610 ;
        RECT 149.800 121.310 150.880 121.610 ;
        RECT 142.900 120.290 143.200 121.310 ;
        RECT 143.680 121.170 144.600 121.210 ;
        RECT 147.640 121.170 148.560 121.210 ;
        RECT 143.680 120.870 144.760 121.170 ;
        RECT 147.640 120.870 148.720 121.170 ;
        RECT 143.680 120.290 144.600 120.330 ;
        RECT 142.900 119.990 148.720 120.290 ;
        RECT 141.520 119.850 142.440 119.890 ;
        RECT 141.520 119.550 142.600 119.850 ;
        RECT 149.020 119.550 150.880 119.850 ;
        RECT 143.680 119.110 144.760 119.410 ;
        RECT 147.640 119.110 148.720 119.410 ;
        RECT 144.070 118.530 144.370 119.110 ;
        RECT 148.030 118.530 148.330 119.110 ;
        RECT 143.680 118.230 148.720 118.530 ;
        RECT 141.520 117.790 142.600 118.090 ;
        RECT 143.680 117.350 144.760 117.650 ;
        RECT 144.070 116.770 144.370 117.350 ;
        RECT 143.680 116.470 144.760 116.770 ;
        RECT 141.520 116.330 142.440 116.370 ;
        RECT 141.520 116.030 142.600 116.330 ;
        RECT 143.680 115.890 144.600 115.930 ;
        RECT 147.040 115.890 147.340 118.230 ;
        RECT 147.640 117.650 148.560 117.690 ;
        RECT 147.640 117.350 148.720 117.650 ;
        RECT 147.640 116.770 148.560 116.810 ;
        RECT 147.640 116.470 148.720 116.770 ;
        RECT 143.680 115.590 144.760 115.890 ;
        RECT 147.040 115.590 148.720 115.890 ;
        RECT 143.680 115.010 144.600 115.050 ;
        RECT 143.680 114.710 148.720 115.010 ;
        RECT 141.520 114.270 142.600 114.570 ;
        RECT 142.300 113.970 143.200 114.270 ;
        RECT 141.520 112.510 142.600 112.810 ;
        RECT 141.520 111.050 142.440 111.090 ;
        RECT 141.520 110.750 142.600 111.050 ;
        RECT 142.900 109.290 143.200 113.970 ;
        RECT 143.680 113.830 144.760 114.130 ;
        RECT 147.640 113.830 148.720 114.130 ;
        RECT 144.070 113.250 144.370 113.830 ;
        RECT 148.030 113.250 148.330 113.830 ;
        RECT 143.680 112.950 144.760 113.250 ;
        RECT 147.640 112.950 148.720 113.250 ;
        RECT 143.680 112.370 144.600 112.410 ;
        RECT 147.640 112.370 148.560 112.410 ;
        RECT 143.680 112.070 144.760 112.370 ;
        RECT 147.640 112.070 148.720 112.370 ;
        RECT 147.640 111.490 148.560 111.530 ;
        RECT 143.680 111.190 148.720 111.490 ;
        RECT 143.680 110.610 144.600 110.650 ;
        RECT 147.640 110.610 148.560 110.650 ;
        RECT 143.680 110.310 144.760 110.610 ;
        RECT 147.640 110.310 148.720 110.610 ;
        RECT 143.680 109.730 144.600 109.770 ;
        RECT 143.680 109.430 148.720 109.730 ;
        RECT 141.520 108.990 143.200 109.290 ;
        RECT 141.520 107.230 142.600 107.530 ;
        RECT 141.520 105.770 142.440 105.810 ;
        RECT 141.520 105.470 142.600 105.770 ;
        RECT 141.520 103.710 142.600 104.010 ;
        RECT 142.900 102.690 143.200 108.990 ;
        RECT 143.680 108.550 144.760 108.850 ;
        RECT 144.070 107.970 144.370 108.550 ;
        RECT 143.680 107.670 144.760 107.970 ;
        RECT 143.680 107.090 144.600 107.130 ;
        RECT 143.680 106.790 144.760 107.090 ;
        RECT 145.060 106.210 145.360 109.430 ;
        RECT 147.640 108.550 148.720 108.850 ;
        RECT 148.030 107.970 148.330 108.550 ;
        RECT 147.640 107.670 148.720 107.970 ;
        RECT 147.640 107.090 148.560 107.130 ;
        RECT 147.640 106.790 148.720 107.090 ;
        RECT 143.680 105.910 148.720 106.210 ;
        RECT 149.020 105.770 149.320 119.550 ;
        RECT 149.800 118.090 150.720 118.130 ;
        RECT 149.800 117.790 150.880 118.090 ;
        RECT 149.800 116.030 150.880 116.330 ;
        RECT 149.800 114.570 150.720 114.610 ;
        RECT 149.800 114.270 150.880 114.570 ;
        RECT 149.800 112.810 150.720 112.850 ;
        RECT 149.800 112.510 150.880 112.810 ;
        RECT 149.800 110.750 150.880 111.050 ;
        RECT 149.800 109.290 150.720 109.330 ;
        RECT 149.800 108.990 150.880 109.290 ;
        RECT 149.800 107.530 150.720 107.570 ;
        RECT 149.800 107.230 150.880 107.530 ;
        RECT 149.020 105.470 150.880 105.770 ;
        RECT 143.680 105.030 144.760 105.330 ;
        RECT 147.640 105.030 148.720 105.330 ;
        RECT 144.070 104.450 144.370 105.030 ;
        RECT 148.030 104.450 148.330 105.030 ;
        RECT 143.680 104.150 144.760 104.450 ;
        RECT 147.640 104.150 148.720 104.450 ;
        RECT 143.680 103.570 144.600 103.610 ;
        RECT 147.640 103.570 148.560 103.610 ;
        RECT 143.680 103.270 144.760 103.570 ;
        RECT 147.640 103.270 148.720 103.570 ;
        RECT 149.020 102.690 149.320 105.470 ;
        RECT 149.800 103.710 150.880 104.010 ;
        RECT 142.900 102.390 149.320 102.690 ;
        RECT 141.520 101.950 142.600 102.250 ;
        RECT 149.800 101.950 150.880 102.250 ;
        RECT 143.680 101.810 144.600 101.850 ;
        RECT 147.640 101.810 148.560 101.850 ;
        RECT 143.680 101.510 144.760 101.810 ;
        RECT 147.640 101.510 148.720 101.810 ;
        RECT 149.020 101.650 150.100 101.950 ;
        RECT 143.680 100.930 144.600 100.970 ;
        RECT 147.640 100.930 148.560 100.970 ;
        RECT 143.680 100.630 145.360 100.930 ;
        RECT 147.640 100.630 148.720 100.930 ;
        RECT 141.520 100.490 142.440 100.530 ;
        RECT 141.520 100.190 142.600 100.490 ;
        RECT 145.060 100.050 145.360 100.630 ;
        RECT 143.680 99.750 144.760 100.050 ;
        RECT 145.060 99.750 148.720 100.050 ;
        RECT 144.070 99.170 144.370 99.750 ;
        RECT 145.060 99.170 145.360 99.750 ;
        RECT 147.640 99.170 148.560 99.210 ;
        RECT 149.020 99.170 149.320 101.650 ;
        RECT 149.800 100.190 150.880 100.490 ;
        RECT 143.680 98.870 144.760 99.170 ;
        RECT 145.060 98.870 149.320 99.170 ;
        RECT 141.520 98.430 142.600 98.730 ;
        RECT 149.800 98.430 150.880 98.730 ;
        RECT 143.680 98.290 144.600 98.330 ;
        RECT 147.640 98.290 148.560 98.330 ;
        RECT 143.680 97.990 144.760 98.290 ;
        RECT 147.640 97.990 148.720 98.290 ;
        RECT 147.640 97.410 148.560 97.450 ;
        RECT 143.680 97.110 148.720 97.410 ;
        RECT 141.520 96.670 143.200 96.970 ;
        RECT 149.800 96.670 150.880 96.970 ;
        RECT 142.900 95.650 143.200 96.670 ;
        RECT 143.680 96.530 144.600 96.570 ;
        RECT 147.640 96.530 148.560 96.570 ;
        RECT 143.680 96.230 144.760 96.530 ;
        RECT 147.640 96.230 148.720 96.530 ;
        RECT 143.680 95.650 144.600 95.690 ;
        RECT 142.900 95.350 148.720 95.650 ;
        RECT 141.520 95.210 142.440 95.250 ;
        RECT 141.520 94.910 142.600 95.210 ;
        RECT 149.020 94.910 150.880 95.210 ;
        RECT 143.680 94.470 144.760 94.770 ;
        RECT 147.640 94.470 148.720 94.770 ;
        RECT 144.070 93.890 144.370 94.470 ;
        RECT 148.030 93.890 148.330 94.470 ;
        RECT 143.680 93.590 148.720 93.890 ;
        RECT 141.520 93.150 142.600 93.450 ;
        RECT 143.680 92.710 144.760 93.010 ;
        RECT 144.070 92.130 144.370 92.710 ;
        RECT 143.680 91.830 144.760 92.130 ;
        RECT 141.520 91.690 142.440 91.730 ;
        RECT 141.520 91.390 142.600 91.690 ;
        RECT 143.680 91.250 144.600 91.290 ;
        RECT 147.040 91.250 147.340 93.590 ;
        RECT 147.640 93.010 148.560 93.050 ;
        RECT 147.640 92.710 148.720 93.010 ;
        RECT 147.640 92.130 148.560 92.170 ;
        RECT 147.640 91.830 148.720 92.130 ;
        RECT 143.680 90.950 144.760 91.250 ;
        RECT 147.040 90.950 148.720 91.250 ;
        RECT 143.680 90.370 144.600 90.410 ;
        RECT 143.680 90.070 148.720 90.370 ;
        RECT 141.520 89.630 142.600 89.930 ;
        RECT 142.300 89.330 143.200 89.630 ;
        RECT 141.520 87.870 142.600 88.170 ;
        RECT 141.520 86.410 142.440 86.450 ;
        RECT 141.520 86.110 142.600 86.410 ;
        RECT 142.900 84.650 143.200 89.330 ;
        RECT 143.680 89.190 144.760 89.490 ;
        RECT 147.640 89.190 148.720 89.490 ;
        RECT 144.070 88.610 144.370 89.190 ;
        RECT 148.030 88.610 148.330 89.190 ;
        RECT 143.680 88.310 144.760 88.610 ;
        RECT 147.640 88.310 148.720 88.610 ;
        RECT 143.680 87.730 144.600 87.770 ;
        RECT 147.640 87.730 148.560 87.770 ;
        RECT 143.680 87.430 144.760 87.730 ;
        RECT 147.640 87.430 148.720 87.730 ;
        RECT 147.640 86.850 148.560 86.890 ;
        RECT 143.680 86.550 148.720 86.850 ;
        RECT 143.680 85.970 144.600 86.010 ;
        RECT 147.640 85.970 148.560 86.010 ;
        RECT 143.680 85.670 144.760 85.970 ;
        RECT 147.640 85.670 148.720 85.970 ;
        RECT 143.680 85.090 144.600 85.130 ;
        RECT 143.680 84.790 148.720 85.090 ;
        RECT 141.520 84.350 143.200 84.650 ;
        RECT 141.520 82.590 142.600 82.890 ;
        RECT 141.520 81.130 142.440 81.170 ;
        RECT 141.520 80.830 142.600 81.130 ;
        RECT 141.520 79.070 142.600 79.370 ;
        RECT 142.900 78.050 143.200 84.350 ;
        RECT 143.680 83.910 144.760 84.210 ;
        RECT 144.070 83.330 144.370 83.910 ;
        RECT 143.680 83.030 144.760 83.330 ;
        RECT 143.680 82.450 144.600 82.490 ;
        RECT 143.680 82.150 144.760 82.450 ;
        RECT 145.060 81.570 145.360 84.790 ;
        RECT 147.640 83.910 148.720 84.210 ;
        RECT 148.030 83.330 148.330 83.910 ;
        RECT 147.640 83.030 148.720 83.330 ;
        RECT 147.640 82.450 148.560 82.490 ;
        RECT 147.640 82.150 148.720 82.450 ;
        RECT 143.680 81.270 148.720 81.570 ;
        RECT 149.020 81.130 149.320 94.910 ;
        RECT 149.800 93.450 150.720 93.490 ;
        RECT 149.800 93.150 150.880 93.450 ;
        RECT 149.800 91.390 150.880 91.690 ;
        RECT 149.800 89.930 150.720 89.970 ;
        RECT 149.800 89.630 150.880 89.930 ;
        RECT 149.800 88.170 150.720 88.210 ;
        RECT 149.800 87.870 150.880 88.170 ;
        RECT 149.800 86.110 150.880 86.410 ;
        RECT 149.800 84.650 150.720 84.690 ;
        RECT 149.800 84.350 150.880 84.650 ;
        RECT 149.800 82.890 150.720 82.930 ;
        RECT 149.800 82.590 150.880 82.890 ;
        RECT 149.020 80.830 150.880 81.130 ;
        RECT 143.680 80.390 144.760 80.690 ;
        RECT 147.640 80.390 148.720 80.690 ;
        RECT 144.070 79.810 144.370 80.390 ;
        RECT 148.030 79.810 148.330 80.390 ;
        RECT 143.680 79.510 144.760 79.810 ;
        RECT 147.640 79.510 148.720 79.810 ;
        RECT 143.680 78.930 144.600 78.970 ;
        RECT 147.640 78.930 148.560 78.970 ;
        RECT 143.680 78.630 144.760 78.930 ;
        RECT 147.640 78.630 148.720 78.930 ;
        RECT 149.020 78.050 149.320 80.830 ;
        RECT 149.800 79.070 150.880 79.370 ;
        RECT 142.900 77.750 149.320 78.050 ;
        RECT 141.520 77.310 142.600 77.610 ;
        RECT 149.800 77.310 150.880 77.610 ;
        RECT 143.680 77.170 144.600 77.210 ;
        RECT 147.640 77.170 148.560 77.210 ;
        RECT 143.680 76.870 144.760 77.170 ;
        RECT 147.640 76.870 148.720 77.170 ;
        RECT 149.020 77.010 150.100 77.310 ;
        RECT 143.680 76.290 144.600 76.330 ;
        RECT 147.640 76.290 148.560 76.330 ;
        RECT 143.680 75.990 145.360 76.290 ;
        RECT 147.640 75.990 148.720 76.290 ;
        RECT 141.520 75.850 142.440 75.890 ;
        RECT 141.520 75.550 142.600 75.850 ;
        RECT 145.060 75.410 145.360 75.990 ;
        RECT 143.680 75.110 144.760 75.410 ;
        RECT 145.060 75.110 148.720 75.410 ;
        RECT 144.070 74.530 144.370 75.110 ;
        RECT 145.060 74.530 145.360 75.110 ;
        RECT 147.640 74.530 148.560 74.570 ;
        RECT 149.020 74.530 149.320 77.010 ;
        RECT 149.800 75.550 150.880 75.850 ;
        RECT 143.680 74.230 144.760 74.530 ;
        RECT 145.060 74.230 149.320 74.530 ;
        RECT 141.520 73.790 142.600 74.090 ;
        RECT 149.800 73.790 150.880 74.090 ;
        RECT 143.680 73.650 144.600 73.690 ;
        RECT 147.640 73.650 148.560 73.690 ;
        RECT 143.680 73.350 144.760 73.650 ;
        RECT 147.640 73.350 148.720 73.650 ;
        RECT 147.640 72.770 148.560 72.810 ;
        RECT 143.680 72.470 148.720 72.770 ;
        RECT 141.520 72.030 143.200 72.330 ;
        RECT 149.800 72.030 150.880 72.330 ;
        RECT 142.900 71.010 143.200 72.030 ;
        RECT 143.680 71.890 144.600 71.930 ;
        RECT 147.640 71.890 148.560 71.930 ;
        RECT 143.680 71.590 144.760 71.890 ;
        RECT 147.640 71.590 148.720 71.890 ;
        RECT 143.680 71.010 144.600 71.050 ;
        RECT 142.900 70.710 148.720 71.010 ;
        RECT 141.520 70.570 142.440 70.610 ;
        RECT 141.520 70.270 142.600 70.570 ;
        RECT 149.020 70.270 150.880 70.570 ;
        RECT 143.680 69.830 144.760 70.130 ;
        RECT 147.640 69.830 148.720 70.130 ;
        RECT 144.070 69.250 144.370 69.830 ;
        RECT 148.030 69.250 148.330 69.830 ;
        RECT 143.680 68.950 148.720 69.250 ;
        RECT 141.520 68.510 142.600 68.810 ;
        RECT 143.680 68.070 144.760 68.370 ;
        RECT 144.070 67.490 144.370 68.070 ;
        RECT 143.680 67.190 144.760 67.490 ;
        RECT 141.520 67.050 142.440 67.090 ;
        RECT 141.520 66.750 142.600 67.050 ;
        RECT 143.680 66.610 144.600 66.650 ;
        RECT 147.040 66.610 147.340 68.950 ;
        RECT 147.640 68.370 148.560 68.410 ;
        RECT 147.640 68.070 148.720 68.370 ;
        RECT 147.640 67.490 148.560 67.530 ;
        RECT 147.640 67.190 148.720 67.490 ;
        RECT 143.680 66.310 144.760 66.610 ;
        RECT 147.040 66.310 148.720 66.610 ;
        RECT 143.680 65.730 144.600 65.770 ;
        RECT 143.680 65.430 148.720 65.730 ;
        RECT 141.520 64.990 142.600 65.290 ;
        RECT 142.300 64.690 143.200 64.990 ;
        RECT 141.520 63.230 142.600 63.530 ;
        RECT 141.520 61.770 142.440 61.810 ;
        RECT 141.520 61.470 142.600 61.770 ;
        RECT 142.900 60.010 143.200 64.690 ;
        RECT 143.680 64.550 144.760 64.850 ;
        RECT 147.640 64.550 148.720 64.850 ;
        RECT 144.070 63.970 144.370 64.550 ;
        RECT 148.030 63.970 148.330 64.550 ;
        RECT 143.680 63.670 144.760 63.970 ;
        RECT 147.640 63.670 148.720 63.970 ;
        RECT 143.680 63.090 144.600 63.130 ;
        RECT 147.640 63.090 148.560 63.130 ;
        RECT 143.680 62.790 144.760 63.090 ;
        RECT 147.640 62.790 148.720 63.090 ;
        RECT 147.640 62.210 148.560 62.250 ;
        RECT 143.680 61.910 148.720 62.210 ;
        RECT 143.680 61.330 144.600 61.370 ;
        RECT 147.640 61.330 148.560 61.370 ;
        RECT 143.680 61.030 144.760 61.330 ;
        RECT 147.640 61.030 148.720 61.330 ;
        RECT 143.680 60.450 144.600 60.490 ;
        RECT 143.680 60.150 148.720 60.450 ;
        RECT 141.520 59.710 143.200 60.010 ;
        RECT 141.520 57.950 142.600 58.250 ;
        RECT 141.520 56.490 142.440 56.530 ;
        RECT 141.520 56.190 142.600 56.490 ;
        RECT 141.520 54.430 142.600 54.730 ;
        RECT 142.900 53.410 143.200 59.710 ;
        RECT 143.680 59.270 144.760 59.570 ;
        RECT 144.070 58.690 144.370 59.270 ;
        RECT 143.680 58.390 144.760 58.690 ;
        RECT 143.680 57.810 144.600 57.850 ;
        RECT 143.680 57.510 144.760 57.810 ;
        RECT 145.060 56.930 145.360 60.150 ;
        RECT 147.640 59.270 148.720 59.570 ;
        RECT 148.030 58.690 148.330 59.270 ;
        RECT 147.640 58.390 148.720 58.690 ;
        RECT 147.640 57.810 148.560 57.850 ;
        RECT 147.640 57.510 148.720 57.810 ;
        RECT 143.680 56.630 148.720 56.930 ;
        RECT 149.020 56.490 149.320 70.270 ;
        RECT 149.800 68.810 150.720 68.850 ;
        RECT 149.800 68.510 150.880 68.810 ;
        RECT 149.800 66.750 150.880 67.050 ;
        RECT 149.800 65.290 150.720 65.330 ;
        RECT 149.800 64.990 150.880 65.290 ;
        RECT 149.800 63.530 150.720 63.570 ;
        RECT 149.800 63.230 150.880 63.530 ;
        RECT 149.800 61.470 150.880 61.770 ;
        RECT 149.800 60.010 150.720 60.050 ;
        RECT 149.800 59.710 150.880 60.010 ;
        RECT 149.800 58.250 150.720 58.290 ;
        RECT 149.800 57.950 150.880 58.250 ;
        RECT 149.020 56.190 150.880 56.490 ;
        RECT 143.680 55.750 144.760 56.050 ;
        RECT 147.640 55.750 148.720 56.050 ;
        RECT 144.070 55.170 144.370 55.750 ;
        RECT 148.030 55.170 148.330 55.750 ;
        RECT 143.680 54.870 144.760 55.170 ;
        RECT 147.640 54.870 148.720 55.170 ;
        RECT 143.680 54.290 144.600 54.330 ;
        RECT 147.640 54.290 148.560 54.330 ;
        RECT 143.680 53.990 144.760 54.290 ;
        RECT 147.640 53.990 148.720 54.290 ;
        RECT 149.020 53.410 149.320 56.190 ;
        RECT 149.800 54.430 150.880 54.730 ;
        RECT 142.900 53.110 149.320 53.410 ;
        RECT 141.520 52.670 142.600 52.970 ;
        RECT 149.800 52.670 150.880 52.970 ;
        RECT 143.680 52.530 144.600 52.570 ;
        RECT 147.640 52.530 148.560 52.570 ;
        RECT 143.680 52.230 144.760 52.530 ;
        RECT 147.640 52.230 148.720 52.530 ;
        RECT 149.020 52.370 150.100 52.670 ;
        RECT 143.680 51.650 144.600 51.690 ;
        RECT 147.640 51.650 148.560 51.690 ;
        RECT 143.680 51.350 145.360 51.650 ;
        RECT 147.640 51.350 148.720 51.650 ;
        RECT 141.520 51.210 142.440 51.250 ;
        RECT 141.520 50.910 142.600 51.210 ;
        RECT 145.060 50.770 145.360 51.350 ;
        RECT 143.680 50.470 144.760 50.770 ;
        RECT 145.060 50.470 148.720 50.770 ;
        RECT 144.070 49.890 144.370 50.470 ;
        RECT 145.060 49.890 145.360 50.470 ;
        RECT 147.640 49.890 148.560 49.930 ;
        RECT 149.020 49.890 149.320 52.370 ;
        RECT 149.800 50.910 150.880 51.210 ;
        RECT 143.680 49.590 144.760 49.890 ;
        RECT 145.060 49.590 149.320 49.890 ;
        RECT 141.520 49.150 142.600 49.450 ;
        RECT 149.800 49.150 150.880 49.450 ;
        RECT 143.680 49.010 144.600 49.050 ;
        RECT 147.640 49.010 148.560 49.050 ;
        RECT 143.680 48.710 144.760 49.010 ;
        RECT 147.640 48.710 148.720 49.010 ;
        RECT 147.640 48.130 148.560 48.170 ;
        RECT 143.680 47.830 148.720 48.130 ;
        RECT 141.520 47.390 143.200 47.690 ;
        RECT 149.800 47.390 150.880 47.690 ;
        RECT 142.900 46.370 143.200 47.390 ;
        RECT 143.680 47.250 144.600 47.290 ;
        RECT 147.640 47.250 148.560 47.290 ;
        RECT 143.680 46.950 144.760 47.250 ;
        RECT 147.640 46.950 148.720 47.250 ;
        RECT 143.680 46.370 144.600 46.410 ;
        RECT 142.900 46.070 148.720 46.370 ;
        RECT 141.520 45.930 142.440 45.970 ;
        RECT 141.520 45.630 142.600 45.930 ;
        RECT 149.020 45.630 150.880 45.930 ;
        RECT 143.680 45.190 144.760 45.490 ;
        RECT 147.640 45.190 148.720 45.490 ;
        RECT 144.070 44.610 144.370 45.190 ;
        RECT 148.030 44.610 148.330 45.190 ;
        RECT 143.680 44.310 148.720 44.610 ;
        RECT 141.520 43.870 142.600 44.170 ;
        RECT 143.680 43.430 144.760 43.730 ;
        RECT 144.070 42.850 144.370 43.430 ;
        RECT 143.680 42.550 144.760 42.850 ;
        RECT 141.520 42.410 142.440 42.450 ;
        RECT 141.520 42.110 142.600 42.410 ;
        RECT 143.680 41.970 144.600 42.010 ;
        RECT 147.040 41.970 147.340 44.310 ;
        RECT 147.640 43.730 148.560 43.770 ;
        RECT 147.640 43.430 148.720 43.730 ;
        RECT 147.640 42.850 148.560 42.890 ;
        RECT 147.640 42.550 148.720 42.850 ;
        RECT 143.680 41.670 144.760 41.970 ;
        RECT 147.040 41.670 148.720 41.970 ;
        RECT 143.680 41.090 144.600 41.130 ;
        RECT 143.680 40.790 148.720 41.090 ;
        RECT 141.520 40.350 142.600 40.650 ;
        RECT 142.300 40.050 143.200 40.350 ;
        RECT 141.520 38.590 142.600 38.890 ;
        RECT 141.520 37.130 142.440 37.170 ;
        RECT 141.520 36.830 142.600 37.130 ;
        RECT 142.900 35.370 143.200 40.050 ;
        RECT 143.680 39.910 144.760 40.210 ;
        RECT 147.640 39.910 148.720 40.210 ;
        RECT 144.070 39.330 144.370 39.910 ;
        RECT 148.030 39.330 148.330 39.910 ;
        RECT 143.680 39.030 144.760 39.330 ;
        RECT 147.640 39.030 148.720 39.330 ;
        RECT 143.680 38.450 144.600 38.490 ;
        RECT 147.640 38.450 148.560 38.490 ;
        RECT 143.680 38.150 144.760 38.450 ;
        RECT 147.640 38.150 148.720 38.450 ;
        RECT 147.640 37.570 148.560 37.610 ;
        RECT 143.680 37.270 148.720 37.570 ;
        RECT 143.680 36.690 144.600 36.730 ;
        RECT 147.640 36.690 148.560 36.730 ;
        RECT 143.680 36.390 144.760 36.690 ;
        RECT 147.640 36.390 148.720 36.690 ;
        RECT 143.680 35.810 144.600 35.850 ;
        RECT 143.680 35.510 148.720 35.810 ;
        RECT 141.520 35.070 143.200 35.370 ;
        RECT 141.520 33.310 142.600 33.610 ;
        RECT 141.520 31.850 142.440 31.890 ;
        RECT 141.520 31.550 142.600 31.850 ;
        RECT 141.520 29.790 142.600 30.090 ;
        RECT 142.900 28.770 143.200 35.070 ;
        RECT 143.680 34.630 144.760 34.930 ;
        RECT 144.070 34.050 144.370 34.630 ;
        RECT 143.680 33.750 144.760 34.050 ;
        RECT 143.680 33.170 144.600 33.210 ;
        RECT 143.680 32.870 144.760 33.170 ;
        RECT 145.060 32.290 145.360 35.510 ;
        RECT 147.640 34.630 148.720 34.930 ;
        RECT 148.030 34.050 148.330 34.630 ;
        RECT 147.640 33.750 148.720 34.050 ;
        RECT 147.640 33.170 148.560 33.210 ;
        RECT 147.640 32.870 148.720 33.170 ;
        RECT 143.680 31.990 148.720 32.290 ;
        RECT 149.020 31.850 149.320 45.630 ;
        RECT 149.800 44.170 150.720 44.210 ;
        RECT 149.800 43.870 150.880 44.170 ;
        RECT 149.800 42.110 150.880 42.410 ;
        RECT 149.800 40.650 150.720 40.690 ;
        RECT 149.800 40.350 150.880 40.650 ;
        RECT 149.800 38.890 150.720 38.930 ;
        RECT 149.800 38.590 150.880 38.890 ;
        RECT 149.800 36.830 150.880 37.130 ;
        RECT 149.800 35.370 150.720 35.410 ;
        RECT 149.800 35.070 150.880 35.370 ;
        RECT 149.800 33.610 150.720 33.650 ;
        RECT 149.800 33.310 150.880 33.610 ;
        RECT 149.020 31.550 150.880 31.850 ;
        RECT 143.680 31.110 144.760 31.410 ;
        RECT 147.640 31.110 148.720 31.410 ;
        RECT 144.070 30.530 144.370 31.110 ;
        RECT 148.030 30.530 148.330 31.110 ;
        RECT 143.680 30.230 144.760 30.530 ;
        RECT 147.640 30.230 148.720 30.530 ;
        RECT 143.680 29.650 144.600 29.690 ;
        RECT 147.640 29.650 148.560 29.690 ;
        RECT 143.680 29.350 144.760 29.650 ;
        RECT 147.640 29.350 148.720 29.650 ;
        RECT 149.020 28.770 149.320 31.550 ;
        RECT 149.800 29.790 150.880 30.090 ;
        RECT 142.900 28.470 149.320 28.770 ;
        RECT 141.520 28.030 142.600 28.330 ;
        RECT 149.800 28.030 150.880 28.330 ;
        RECT 143.680 27.890 144.600 27.930 ;
        RECT 147.640 27.890 148.560 27.930 ;
        RECT 143.680 27.590 144.760 27.890 ;
        RECT 147.640 27.590 148.720 27.890 ;
        RECT 149.020 27.730 150.100 28.030 ;
        RECT 143.680 27.010 144.600 27.050 ;
        RECT 147.640 27.010 148.560 27.050 ;
        RECT 143.680 26.710 145.360 27.010 ;
        RECT 147.640 26.710 148.720 27.010 ;
        RECT 141.520 26.570 142.440 26.610 ;
        RECT 141.520 26.270 142.600 26.570 ;
        RECT 145.060 26.130 145.360 26.710 ;
        RECT 143.680 25.830 144.760 26.130 ;
        RECT 145.060 25.830 148.720 26.130 ;
        RECT 144.070 25.250 144.370 25.830 ;
        RECT 145.060 25.250 145.360 25.830 ;
        RECT 147.640 25.250 148.560 25.290 ;
        RECT 149.020 25.250 149.320 27.730 ;
        RECT 149.800 26.270 150.880 26.570 ;
        RECT 143.680 24.950 144.760 25.250 ;
        RECT 145.060 24.950 149.320 25.250 ;
        RECT 141.520 24.510 142.600 24.810 ;
        RECT 149.800 24.510 150.880 24.810 ;
        RECT 143.680 24.370 144.600 24.410 ;
        RECT 147.640 24.370 148.560 24.410 ;
        RECT 143.680 24.070 144.760 24.370 ;
        RECT 147.640 24.070 148.720 24.370 ;
        RECT 143.680 23.190 148.720 23.490 ;
        RECT 141.520 22.750 143.200 23.050 ;
        RECT 149.800 22.750 150.880 23.050 ;
        RECT 142.900 21.730 143.200 22.750 ;
        RECT 143.680 22.610 144.600 22.650 ;
        RECT 147.640 22.610 148.560 22.650 ;
        RECT 143.680 22.310 144.760 22.610 ;
        RECT 147.640 22.310 148.720 22.610 ;
        RECT 147.640 21.730 148.560 21.770 ;
        RECT 142.900 21.430 145.360 21.730 ;
        RECT 147.640 21.430 148.720 21.730 ;
        RECT 141.520 20.990 142.600 21.290 ;
        RECT 145.060 20.850 145.360 21.430 ;
        RECT 149.800 20.990 150.880 21.290 ;
        RECT 143.680 20.550 144.760 20.850 ;
        RECT 145.060 20.550 148.720 20.850 ;
        RECT 144.070 19.970 144.370 20.550 ;
        RECT 145.060 19.970 145.360 20.550 ;
        RECT 143.680 19.670 144.760 19.970 ;
        RECT 145.060 19.670 148.720 19.970 ;
        RECT 141.520 19.230 142.600 19.530 ;
        RECT 149.800 19.230 150.880 19.530 ;
        RECT 143.680 19.090 144.600 19.130 ;
        RECT 147.640 19.090 148.560 19.130 ;
        RECT 143.680 18.790 144.760 19.090 ;
        RECT 147.640 18.790 148.720 19.090 ;
        RECT 143.680 17.910 148.720 18.210 ;
        RECT 141.520 17.470 142.600 17.770 ;
        RECT 149.800 17.470 150.880 17.770 ;
        RECT 143.680 17.330 144.600 17.370 ;
        RECT 147.640 17.330 148.560 17.370 ;
        RECT 143.680 17.030 144.760 17.330 ;
        RECT 147.640 17.030 148.720 17.330 ;
        RECT 143.680 16.150 148.720 16.450 ;
        RECT 141.520 15.710 143.200 16.010 ;
        RECT 149.800 15.710 150.880 16.010 ;
        RECT 141.520 13.950 142.600 14.250 ;
        RECT 142.900 13.810 143.200 15.710 ;
        RECT 143.680 15.570 144.600 15.610 ;
        RECT 147.640 15.570 148.560 15.610 ;
        RECT 143.680 15.270 144.760 15.570 ;
        RECT 147.640 15.270 148.720 15.570 ;
        RECT 143.680 14.690 144.600 14.730 ;
        RECT 143.680 14.390 144.760 14.690 ;
        RECT 145.060 14.390 148.720 14.690 ;
        RECT 145.060 13.810 145.360 14.390 ;
        RECT 149.800 13.950 150.880 14.250 ;
        RECT 142.900 13.510 145.360 13.810 ;
        RECT 147.640 13.510 148.720 13.810 ;
        RECT 145.060 12.930 145.360 13.510 ;
        RECT 148.030 12.930 148.330 13.510 ;
        RECT 143.680 12.630 145.360 12.930 ;
        RECT 147.640 12.630 148.720 12.930 ;
        RECT 141.520 12.190 142.600 12.490 ;
        RECT 149.800 12.190 150.880 12.490 ;
        RECT 143.680 12.050 144.600 12.090 ;
        RECT 147.640 12.050 148.560 12.090 ;
        RECT 143.680 11.750 144.760 12.050 ;
        RECT 147.640 11.750 148.720 12.050 ;
        RECT 143.680 10.870 148.720 11.170 ;
        RECT 141.520 10.430 143.200 10.730 ;
        RECT 149.800 10.430 150.880 10.730 ;
        RECT 141.520 8.670 142.600 8.970 ;
        RECT 142.900 8.530 143.200 10.430 ;
        RECT 143.680 10.290 144.600 10.330 ;
        RECT 147.640 10.290 148.560 10.330 ;
        RECT 143.680 9.990 144.760 10.290 ;
        RECT 147.640 9.990 148.720 10.290 ;
        RECT 143.680 9.410 144.600 9.450 ;
        RECT 147.640 9.410 148.560 9.450 ;
        RECT 143.680 9.110 144.760 9.410 ;
        RECT 147.640 9.110 148.720 9.410 ;
        RECT 149.800 8.670 150.880 8.970 ;
        RECT 142.900 8.230 148.720 8.530 ;
        RECT 143.680 7.350 148.720 7.650 ;
        RECT 141.520 6.910 142.600 7.210 ;
        RECT 149.800 6.910 150.880 7.210 ;
        RECT 143.680 6.770 144.600 6.810 ;
        RECT 147.640 6.770 148.560 6.810 ;
        RECT 143.680 6.470 144.760 6.770 ;
        RECT 147.640 6.470 148.720 6.770 ;
        RECT 143.680 5.590 148.720 5.890 ;
        RECT 141.520 5.150 142.600 5.450 ;
        RECT 149.800 5.150 150.880 5.450 ;
        RECT 143.680 5.010 144.600 5.050 ;
        RECT 147.640 5.010 148.560 5.050 ;
        RECT 143.680 4.710 144.760 5.010 ;
        RECT 147.640 4.710 148.720 5.010 ;
        RECT 143.680 4.130 144.600 4.170 ;
        RECT 147.640 4.130 148.560 4.170 ;
        RECT 142.900 3.830 144.760 4.130 ;
        RECT 147.640 3.830 149.320 4.130 ;
        RECT 142.900 3.690 143.200 3.830 ;
        RECT 139.360 3.390 143.200 3.690 ;
        RECT 139.360 2.440 140.440 3.390 ;
        RECT 142.900 3.250 143.200 3.390 ;
        RECT 149.020 3.690 149.320 3.830 ;
        RECT 151.960 3.690 153.040 221.630 ;
        RECT 149.020 3.390 153.040 3.690 ;
        RECT 143.680 3.250 144.600 3.290 ;
        RECT 147.640 3.250 148.560 3.290 ;
        RECT 149.020 3.250 149.320 3.390 ;
        RECT 142.900 2.950 144.760 3.250 ;
        RECT 147.640 2.950 149.320 3.250 ;
        RECT 151.960 2.440 153.040 3.390 ;
      LAYER mcon ;
        RECT 24.640 221.770 24.920 222.050 ;
        RECT 25.160 221.770 25.440 222.050 ;
        RECT 27.600 221.770 27.880 222.050 ;
        RECT 28.120 221.770 28.400 222.050 ;
        RECT 49.840 221.770 50.120 222.050 ;
        RECT 50.360 221.770 50.640 222.050 ;
        RECT 52.800 221.770 53.080 222.050 ;
        RECT 53.320 221.770 53.600 222.050 ;
        RECT 75.040 221.770 75.320 222.050 ;
        RECT 75.560 221.770 75.840 222.050 ;
        RECT 78.000 221.770 78.280 222.050 ;
        RECT 78.520 221.770 78.800 222.050 ;
        RECT 100.240 221.770 100.520 222.050 ;
        RECT 100.760 221.770 101.040 222.050 ;
        RECT 103.200 221.770 103.480 222.050 ;
        RECT 103.720 221.770 104.000 222.050 ;
        RECT 24.640 221.250 24.920 221.530 ;
        RECT 25.160 221.250 25.440 221.530 ;
        RECT 27.600 221.250 27.880 221.530 ;
        RECT 28.120 221.250 28.400 221.530 ;
        RECT 49.840 221.250 50.120 221.530 ;
        RECT 50.360 221.250 50.640 221.530 ;
        RECT 52.800 221.250 53.080 221.530 ;
        RECT 53.320 221.250 53.600 221.530 ;
        RECT 75.040 221.250 75.320 221.530 ;
        RECT 75.560 221.250 75.840 221.530 ;
        RECT 78.000 221.250 78.280 221.530 ;
        RECT 78.520 221.250 78.800 221.530 ;
        RECT 100.240 221.250 100.520 221.530 ;
        RECT 100.760 221.250 101.040 221.530 ;
        RECT 103.200 221.250 103.480 221.530 ;
        RECT 103.720 221.250 104.000 221.530 ;
        RECT 21.760 218.170 22.040 218.450 ;
        RECT 22.280 218.170 22.560 218.450 ;
        RECT 30.480 218.170 30.760 218.450 ;
        RECT 31.000 218.170 31.280 218.450 ;
        RECT 46.960 218.170 47.240 218.450 ;
        RECT 47.480 218.170 47.760 218.450 ;
        RECT 55.680 218.170 55.960 218.450 ;
        RECT 56.200 218.170 56.480 218.450 ;
        RECT 72.160 218.170 72.440 218.450 ;
        RECT 72.680 218.170 72.960 218.450 ;
        RECT 80.880 218.170 81.160 218.450 ;
        RECT 81.400 218.170 81.680 218.450 ;
        RECT 97.360 218.170 97.640 218.450 ;
        RECT 97.880 218.170 98.160 218.450 ;
        RECT 106.080 218.170 106.360 218.450 ;
        RECT 106.600 218.170 106.880 218.450 ;
        RECT 122.560 218.170 122.840 218.450 ;
        RECT 123.080 218.170 123.360 218.450 ;
        RECT 21.760 217.650 22.040 217.930 ;
        RECT 22.280 217.650 22.560 217.930 ;
        RECT 30.480 217.650 30.760 217.930 ;
        RECT 31.000 217.650 31.280 217.930 ;
        RECT 46.960 217.650 47.240 217.930 ;
        RECT 47.480 217.650 47.760 217.930 ;
        RECT 55.680 217.650 55.960 217.930 ;
        RECT 56.200 217.650 56.480 217.930 ;
        RECT 72.160 217.650 72.440 217.930 ;
        RECT 72.680 217.650 72.960 217.930 ;
        RECT 80.880 217.650 81.160 217.930 ;
        RECT 81.400 217.650 81.680 217.930 ;
        RECT 97.360 217.650 97.640 217.930 ;
        RECT 97.880 217.650 98.160 217.930 ;
        RECT 106.080 217.650 106.360 217.930 ;
        RECT 106.600 217.650 106.880 217.930 ;
        RECT 122.560 217.650 122.840 217.930 ;
        RECT 123.080 217.650 123.360 217.930 ;
        RECT 4.030 207.110 4.310 207.390 ;
        RECT 4.030 206.590 4.310 206.870 ;
        RECT 17.800 214.570 18.080 214.850 ;
        RECT 18.320 214.570 18.600 214.850 ;
        RECT 34.440 214.570 34.720 214.850 ;
        RECT 34.960 214.570 35.240 214.850 ;
        RECT 43.000 214.570 43.280 214.850 ;
        RECT 43.520 214.570 43.800 214.850 ;
        RECT 59.640 214.570 59.920 214.850 ;
        RECT 60.160 214.570 60.440 214.850 ;
        RECT 68.200 214.570 68.480 214.850 ;
        RECT 68.720 214.570 69.000 214.850 ;
        RECT 84.840 214.570 85.120 214.850 ;
        RECT 85.360 214.570 85.640 214.850 ;
        RECT 93.400 214.570 93.680 214.850 ;
        RECT 93.920 214.570 94.200 214.850 ;
        RECT 110.040 214.570 110.320 214.850 ;
        RECT 110.560 214.570 110.840 214.850 ;
        RECT 118.600 214.570 118.880 214.850 ;
        RECT 119.120 214.570 119.400 214.850 ;
        RECT 17.800 214.050 18.080 214.330 ;
        RECT 18.320 214.050 18.600 214.330 ;
        RECT 34.440 214.050 34.720 214.330 ;
        RECT 34.960 214.050 35.240 214.330 ;
        RECT 43.000 214.050 43.280 214.330 ;
        RECT 43.520 214.050 43.800 214.330 ;
        RECT 59.640 214.050 59.920 214.330 ;
        RECT 60.160 214.050 60.440 214.330 ;
        RECT 68.200 214.050 68.480 214.330 ;
        RECT 68.720 214.050 69.000 214.330 ;
        RECT 84.840 214.050 85.120 214.330 ;
        RECT 85.360 214.050 85.640 214.330 ;
        RECT 93.400 214.050 93.680 214.330 ;
        RECT 93.920 214.050 94.200 214.330 ;
        RECT 110.040 214.050 110.320 214.330 ;
        RECT 110.560 214.050 110.840 214.330 ;
        RECT 118.600 214.050 118.880 214.330 ;
        RECT 119.120 214.050 119.400 214.330 ;
        RECT 17.800 210.830 18.080 211.110 ;
        RECT 18.320 210.830 18.600 211.110 ;
        RECT 21.760 210.830 22.040 211.110 ;
        RECT 22.280 210.830 22.560 211.110 ;
        RECT 30.560 210.830 30.840 211.110 ;
        RECT 31.080 210.830 31.360 211.110 ;
        RECT 34.520 210.830 34.800 211.110 ;
        RECT 35.040 210.830 35.320 211.110 ;
        RECT 17.800 209.950 18.080 210.230 ;
        RECT 18.320 209.950 18.600 210.230 ;
        RECT 21.760 209.950 22.040 210.230 ;
        RECT 22.280 209.950 22.560 210.230 ;
        RECT 21.760 209.260 22.040 209.540 ;
        RECT 22.280 209.260 22.560 209.540 ;
        RECT 15.640 206.870 15.920 207.150 ;
        RECT 16.160 206.870 16.440 207.150 ;
        RECT 17.800 208.190 18.080 208.470 ;
        RECT 18.320 208.190 18.600 208.470 ;
        RECT 21.760 208.190 22.040 208.470 ;
        RECT 22.280 208.190 22.560 208.470 ;
        RECT 17.800 207.310 18.080 207.590 ;
        RECT 18.320 207.310 18.600 207.590 ;
        RECT 17.800 204.670 18.080 204.950 ;
        RECT 18.320 204.670 18.600 204.950 ;
        RECT 21.760 204.670 22.040 204.950 ;
        RECT 22.280 204.670 22.560 204.950 ;
        RECT 17.800 202.910 18.080 203.190 ;
        RECT 18.320 202.910 18.600 203.190 ;
        RECT 21.760 202.910 22.040 203.190 ;
        RECT 22.280 202.910 22.560 203.190 ;
        RECT 21.760 202.030 22.040 202.310 ;
        RECT 22.280 202.030 22.560 202.310 ;
        RECT 15.640 201.590 15.920 201.870 ;
        RECT 16.160 201.590 16.440 201.870 ;
        RECT 17.800 199.390 18.080 199.670 ;
        RECT 18.320 199.390 18.600 199.670 ;
        RECT 21.760 199.390 22.040 199.670 ;
        RECT 22.280 199.390 22.560 199.670 ;
        RECT 17.800 197.630 18.080 197.910 ;
        RECT 18.320 197.630 18.600 197.910 ;
        RECT 21.760 197.630 22.040 197.910 ;
        RECT 22.280 197.630 22.560 197.910 ;
        RECT 23.920 196.310 24.200 196.590 ;
        RECT 24.440 196.310 24.720 196.590 ;
        RECT 17.800 195.870 18.080 196.150 ;
        RECT 18.320 195.870 18.600 196.150 ;
        RECT 21.760 195.870 22.040 196.150 ;
        RECT 22.280 195.870 22.560 196.150 ;
        RECT 17.800 194.990 18.080 195.270 ;
        RECT 18.320 194.990 18.600 195.270 ;
        RECT 17.800 192.350 18.080 192.630 ;
        RECT 18.320 192.350 18.600 192.630 ;
        RECT 17.800 191.470 18.080 191.750 ;
        RECT 18.320 191.470 18.600 191.750 ;
        RECT 15.640 191.030 15.920 191.310 ;
        RECT 16.160 191.030 16.440 191.310 ;
        RECT 17.800 188.830 18.080 189.110 ;
        RECT 18.320 188.830 18.600 189.110 ;
        RECT 23.920 192.790 24.200 193.070 ;
        RECT 24.440 192.790 24.720 193.070 ;
        RECT 21.760 192.350 22.040 192.630 ;
        RECT 22.280 192.350 22.560 192.630 ;
        RECT 21.760 191.470 22.040 191.750 ;
        RECT 22.280 191.470 22.560 191.750 ;
        RECT 17.800 187.950 18.080 188.230 ;
        RECT 18.320 187.950 18.600 188.230 ;
        RECT 21.760 187.950 22.040 188.230 ;
        RECT 22.280 187.950 22.560 188.230 ;
        RECT 17.800 185.310 18.080 185.590 ;
        RECT 18.320 185.310 18.600 185.590 ;
        RECT 17.800 184.430 18.080 184.710 ;
        RECT 18.320 184.430 18.600 184.710 ;
        RECT 21.760 184.430 22.040 184.710 ;
        RECT 22.280 184.430 22.560 184.710 ;
        RECT 20.940 182.870 21.220 183.150 ;
        RECT 20.940 182.350 21.220 182.630 ;
        RECT 17.800 181.790 18.080 182.070 ;
        RECT 18.320 181.790 18.600 182.070 ;
        RECT 21.760 181.790 22.040 182.070 ;
        RECT 22.280 181.790 22.560 182.070 ;
        RECT 17.800 180.910 18.080 181.190 ;
        RECT 18.320 180.910 18.600 181.190 ;
        RECT 21.760 180.910 22.040 181.190 ;
        RECT 22.280 180.910 22.560 181.190 ;
        RECT 17.800 178.270 18.080 178.550 ;
        RECT 18.320 178.270 18.600 178.550 ;
        RECT 17.800 177.390 18.080 177.670 ;
        RECT 18.320 177.390 18.600 177.670 ;
        RECT 21.760 177.390 22.040 177.670 ;
        RECT 22.280 177.390 22.560 177.670 ;
        RECT 20.065 175.830 20.345 176.110 ;
        RECT 15.640 175.190 15.920 175.470 ;
        RECT 16.160 175.190 16.440 175.470 ;
        RECT 20.065 175.310 20.345 175.590 ;
        RECT 17.800 174.750 18.080 175.030 ;
        RECT 18.320 174.750 18.600 175.030 ;
        RECT 21.760 174.750 22.040 175.030 ;
        RECT 22.280 174.750 22.560 175.030 ;
        RECT 17.800 173.870 18.080 174.150 ;
        RECT 18.320 173.870 18.600 174.150 ;
        RECT 21.760 173.870 22.040 174.150 ;
        RECT 22.280 173.870 22.560 174.150 ;
        RECT 17.800 171.230 18.080 171.510 ;
        RECT 18.320 171.230 18.600 171.510 ;
        RECT 17.800 170.350 18.080 170.630 ;
        RECT 18.320 170.350 18.600 170.630 ;
        RECT 21.760 170.350 22.040 170.630 ;
        RECT 22.280 170.350 22.560 170.630 ;
        RECT 19.265 168.790 19.545 169.070 ;
        RECT 21.760 168.590 22.040 168.870 ;
        RECT 22.280 168.590 22.560 168.870 ;
        RECT 15.720 168.110 16.000 168.390 ;
        RECT 16.240 168.110 16.520 168.390 ;
        RECT 19.265 168.270 19.545 168.550 ;
        RECT 17.800 167.710 18.080 167.990 ;
        RECT 18.320 167.710 18.600 167.990 ;
        RECT 21.760 167.710 22.040 167.990 ;
        RECT 22.280 167.710 22.560 167.990 ;
        RECT 17.800 166.830 18.080 167.110 ;
        RECT 18.320 166.830 18.600 167.110 ;
        RECT 21.760 166.830 22.040 167.110 ;
        RECT 22.280 166.830 22.560 167.110 ;
        RECT 17.800 164.190 18.080 164.470 ;
        RECT 18.320 164.190 18.600 164.470 ;
        RECT 17.800 163.310 18.080 163.590 ;
        RECT 18.320 163.310 18.600 163.590 ;
        RECT 21.760 163.310 22.040 163.590 ;
        RECT 22.280 163.310 22.560 163.590 ;
        RECT 17.800 160.670 18.080 160.950 ;
        RECT 18.320 160.670 18.600 160.950 ;
        RECT 21.760 160.670 22.040 160.950 ;
        RECT 22.280 160.670 22.560 160.950 ;
        RECT 15.640 159.350 15.920 159.630 ;
        RECT 16.160 159.350 16.440 159.630 ;
        RECT 23.920 159.350 24.200 159.630 ;
        RECT 24.440 159.350 24.720 159.630 ;
        RECT 15.640 155.830 15.920 156.110 ;
        RECT 16.160 155.830 16.440 156.110 ;
        RECT 15.640 154.070 15.920 154.350 ;
        RECT 16.160 154.070 16.440 154.350 ;
        RECT 17.800 155.390 18.080 155.670 ;
        RECT 18.320 155.390 18.600 155.670 ;
        RECT 21.760 155.390 22.040 155.670 ;
        RECT 22.280 155.390 22.560 155.670 ;
        RECT 17.800 154.510 18.080 154.790 ;
        RECT 18.320 154.510 18.600 154.790 ;
        RECT 15.800 150.550 16.080 150.830 ;
        RECT 16.320 150.550 16.600 150.830 ;
        RECT 17.800 150.110 18.080 150.390 ;
        RECT 18.320 150.110 18.600 150.390 ;
        RECT 21.760 150.110 22.040 150.390 ;
        RECT 22.280 150.110 22.560 150.390 ;
        RECT 17.800 148.350 18.080 148.630 ;
        RECT 18.320 148.350 18.600 148.630 ;
        RECT 21.760 148.350 22.040 148.630 ;
        RECT 22.280 148.350 22.560 148.630 ;
        RECT 21.760 147.470 22.040 147.750 ;
        RECT 22.280 147.470 22.560 147.750 ;
        RECT 17.800 146.590 18.080 146.870 ;
        RECT 18.320 146.590 18.600 146.870 ;
        RECT 17.800 145.710 18.080 145.990 ;
        RECT 18.320 145.710 18.600 145.990 ;
        RECT 15.800 145.270 16.080 145.550 ;
        RECT 16.320 145.270 16.600 145.550 ;
        RECT 17.800 143.070 18.080 143.350 ;
        RECT 18.320 143.070 18.600 143.350 ;
        RECT 21.760 143.070 22.040 143.350 ;
        RECT 22.280 143.070 22.560 143.350 ;
        RECT 21.760 142.190 22.040 142.470 ;
        RECT 22.280 142.190 22.560 142.470 ;
        RECT 15.640 141.750 15.920 142.030 ;
        RECT 16.160 141.750 16.440 142.030 ;
        RECT 17.800 140.430 18.080 140.710 ;
        RECT 18.320 140.430 18.600 140.710 ;
        RECT 21.760 140.430 22.040 140.710 ;
        RECT 22.280 140.430 22.560 140.710 ;
        RECT 43.000 210.830 43.280 211.110 ;
        RECT 43.520 210.830 43.800 211.110 ;
        RECT 46.960 210.830 47.240 211.110 ;
        RECT 47.480 210.830 47.760 211.110 ;
        RECT 30.560 209.950 30.840 210.230 ;
        RECT 31.080 209.950 31.360 210.230 ;
        RECT 34.520 209.950 34.800 210.230 ;
        RECT 35.040 209.950 35.320 210.230 ;
        RECT 30.400 209.070 30.680 209.350 ;
        RECT 30.920 209.070 31.200 209.350 ;
        RECT 30.560 208.190 30.840 208.470 ;
        RECT 31.080 208.190 31.360 208.470 ;
        RECT 34.520 208.190 34.800 208.470 ;
        RECT 35.040 208.190 35.320 208.470 ;
        RECT 34.520 207.310 34.800 207.590 ;
        RECT 35.040 207.310 35.320 207.590 ;
        RECT 36.520 206.870 36.800 207.150 ;
        RECT 37.040 206.870 37.320 207.150 ;
        RECT 30.560 204.670 30.840 204.950 ;
        RECT 31.080 204.670 31.360 204.950 ;
        RECT 34.520 204.670 34.800 204.950 ;
        RECT 35.040 204.670 35.320 204.950 ;
        RECT 30.560 202.910 30.840 203.190 ;
        RECT 31.080 202.910 31.360 203.190 ;
        RECT 34.520 202.910 34.800 203.190 ;
        RECT 35.040 202.910 35.320 203.190 ;
        RECT 30.560 202.030 30.840 202.310 ;
        RECT 31.080 202.030 31.360 202.310 ;
        RECT 36.680 201.590 36.960 201.870 ;
        RECT 37.200 201.590 37.480 201.870 ;
        RECT 30.560 199.390 30.840 199.670 ;
        RECT 31.080 199.390 31.360 199.670 ;
        RECT 34.520 199.390 34.800 199.670 ;
        RECT 35.040 199.390 35.320 199.670 ;
        RECT 30.560 197.630 30.840 197.910 ;
        RECT 31.080 197.630 31.360 197.910 ;
        RECT 34.520 197.630 34.800 197.910 ;
        RECT 35.040 197.630 35.320 197.910 ;
        RECT 28.400 196.310 28.680 196.590 ;
        RECT 28.920 196.310 29.200 196.590 ;
        RECT 30.560 195.870 30.840 196.150 ;
        RECT 31.080 195.870 31.360 196.150 ;
        RECT 34.520 195.870 34.800 196.150 ;
        RECT 35.040 195.870 35.320 196.150 ;
        RECT 34.520 194.990 34.800 195.270 ;
        RECT 35.040 194.990 35.320 195.270 ;
        RECT 28.400 192.790 28.680 193.070 ;
        RECT 28.920 192.790 29.200 193.070 ;
        RECT 30.560 192.350 30.840 192.630 ;
        RECT 31.080 192.350 31.360 192.630 ;
        RECT 30.560 191.470 30.840 191.750 ;
        RECT 31.080 191.470 31.360 191.750 ;
        RECT 34.520 192.350 34.800 192.630 ;
        RECT 35.040 192.350 35.320 192.630 ;
        RECT 34.520 191.470 34.800 191.750 ;
        RECT 35.040 191.470 35.320 191.750 ;
        RECT 36.520 191.030 36.800 191.310 ;
        RECT 37.040 191.030 37.320 191.310 ;
        RECT 34.520 188.830 34.800 189.110 ;
        RECT 35.040 188.830 35.320 189.110 ;
        RECT 30.560 187.950 30.840 188.230 ;
        RECT 31.080 187.950 31.360 188.230 ;
        RECT 34.520 187.950 34.800 188.230 ;
        RECT 35.040 187.950 35.320 188.230 ;
        RECT 30.560 184.430 30.840 184.710 ;
        RECT 31.080 184.430 31.360 184.710 ;
        RECT 31.900 182.870 32.180 183.150 ;
        RECT 34.520 185.310 34.800 185.590 ;
        RECT 35.040 185.310 35.320 185.590 ;
        RECT 34.520 184.430 34.800 184.710 ;
        RECT 35.040 184.430 35.320 184.710 ;
        RECT 31.900 182.350 32.180 182.630 ;
        RECT 30.560 181.790 30.840 182.070 ;
        RECT 31.080 181.790 31.360 182.070 ;
        RECT 34.520 181.790 34.800 182.070 ;
        RECT 35.040 181.790 35.320 182.070 ;
        RECT 30.560 180.910 30.840 181.190 ;
        RECT 31.080 180.910 31.360 181.190 ;
        RECT 34.520 180.910 34.800 181.190 ;
        RECT 35.040 180.910 35.320 181.190 ;
        RECT 30.560 177.390 30.840 177.670 ;
        RECT 31.080 177.390 31.360 177.670 ;
        RECT 32.775 175.830 33.055 176.110 ;
        RECT 34.520 178.270 34.800 178.550 ;
        RECT 35.040 178.270 35.320 178.550 ;
        RECT 34.520 177.390 34.800 177.670 ;
        RECT 35.040 177.390 35.320 177.670 ;
        RECT 32.775 175.310 33.055 175.590 ;
        RECT 36.680 175.190 36.960 175.470 ;
        RECT 37.200 175.190 37.480 175.470 ;
        RECT 30.560 174.750 30.840 175.030 ;
        RECT 31.080 174.750 31.360 175.030 ;
        RECT 34.520 174.750 34.800 175.030 ;
        RECT 35.040 174.750 35.320 175.030 ;
        RECT 30.560 173.870 30.840 174.150 ;
        RECT 31.080 173.870 31.360 174.150 ;
        RECT 34.520 173.870 34.800 174.150 ;
        RECT 35.040 173.870 35.320 174.150 ;
        RECT 30.560 170.350 30.840 170.630 ;
        RECT 31.080 170.350 31.360 170.630 ;
        RECT 34.520 171.230 34.800 171.510 ;
        RECT 35.040 171.230 35.320 171.510 ;
        RECT 34.520 170.350 34.800 170.630 ;
        RECT 35.040 170.350 35.320 170.630 ;
        RECT 30.560 168.590 30.840 168.870 ;
        RECT 31.080 168.590 31.360 168.870 ;
        RECT 33.575 168.790 33.855 169.070 ;
        RECT 33.575 168.270 33.855 168.550 ;
        RECT 30.560 167.710 30.840 167.990 ;
        RECT 31.080 167.710 31.360 167.990 ;
        RECT 34.520 167.710 34.800 167.990 ;
        RECT 35.040 167.710 35.320 167.990 ;
        RECT 30.560 166.830 30.840 167.110 ;
        RECT 31.080 166.830 31.360 167.110 ;
        RECT 34.520 166.830 34.800 167.110 ;
        RECT 35.040 166.830 35.320 167.110 ;
        RECT 30.560 163.310 30.840 163.590 ;
        RECT 31.080 163.310 31.360 163.590 ;
        RECT 34.520 164.190 34.800 164.470 ;
        RECT 35.040 164.190 35.320 164.470 ;
        RECT 34.520 163.310 34.800 163.590 ;
        RECT 35.040 163.310 35.320 163.590 ;
        RECT 36.600 168.110 36.880 168.390 ;
        RECT 37.120 168.110 37.400 168.390 ;
        RECT 30.560 160.670 30.840 160.950 ;
        RECT 31.080 160.670 31.360 160.950 ;
        RECT 34.520 160.670 34.800 160.950 ;
        RECT 35.040 160.670 35.320 160.950 ;
        RECT 28.240 159.350 28.520 159.630 ;
        RECT 28.760 159.350 29.040 159.630 ;
        RECT 36.680 159.350 36.960 159.630 ;
        RECT 37.200 159.350 37.480 159.630 ;
        RECT 30.560 155.390 30.840 155.670 ;
        RECT 31.080 155.390 31.360 155.670 ;
        RECT 34.520 155.390 34.800 155.670 ;
        RECT 35.040 155.390 35.320 155.670 ;
        RECT 34.520 154.510 34.800 154.790 ;
        RECT 35.040 154.510 35.320 154.790 ;
        RECT 36.520 155.830 36.800 156.110 ;
        RECT 37.040 155.830 37.320 156.110 ;
        RECT 36.680 154.070 36.960 154.350 ;
        RECT 37.200 154.070 37.480 154.350 ;
        RECT 30.560 150.110 30.840 150.390 ;
        RECT 31.080 150.110 31.360 150.390 ;
        RECT 34.520 150.110 34.800 150.390 ;
        RECT 35.040 150.110 35.320 150.390 ;
        RECT 36.520 150.550 36.800 150.830 ;
        RECT 37.040 150.550 37.320 150.830 ;
        RECT 30.560 148.350 30.840 148.630 ;
        RECT 31.080 148.350 31.360 148.630 ;
        RECT 34.520 148.350 34.800 148.630 ;
        RECT 35.040 148.350 35.320 148.630 ;
        RECT 30.560 147.470 30.840 147.750 ;
        RECT 31.080 147.470 31.360 147.750 ;
        RECT 30.560 143.070 30.840 143.350 ;
        RECT 31.080 143.070 31.360 143.350 ;
        RECT 34.520 146.590 34.800 146.870 ;
        RECT 35.040 146.590 35.320 146.870 ;
        RECT 34.520 145.710 34.800 145.990 ;
        RECT 35.040 145.710 35.320 145.990 ;
        RECT 36.520 145.270 36.800 145.550 ;
        RECT 37.040 145.270 37.320 145.550 ;
        RECT 30.560 142.190 30.840 142.470 ;
        RECT 31.080 142.190 31.360 142.470 ;
        RECT 34.520 143.070 34.800 143.350 ;
        RECT 35.040 143.070 35.320 143.350 ;
        RECT 36.680 141.750 36.960 142.030 ;
        RECT 37.200 141.750 37.480 142.030 ;
        RECT 30.560 140.430 30.840 140.710 ;
        RECT 31.080 140.430 31.360 140.710 ;
        RECT 34.520 140.430 34.800 140.710 ;
        RECT 35.040 140.430 35.320 140.710 ;
        RECT 17.800 139.550 18.080 139.830 ;
        RECT 18.320 139.550 18.600 139.830 ;
        RECT 21.760 139.550 22.040 139.830 ;
        RECT 22.280 139.550 22.560 139.830 ;
        RECT 55.760 210.830 56.040 211.110 ;
        RECT 56.280 210.830 56.560 211.110 ;
        RECT 59.720 210.830 60.000 211.110 ;
        RECT 60.240 210.830 60.520 211.110 ;
        RECT 43.000 209.950 43.280 210.230 ;
        RECT 43.520 209.950 43.800 210.230 ;
        RECT 46.960 209.950 47.240 210.230 ;
        RECT 47.480 209.950 47.760 210.230 ;
        RECT 46.960 209.260 47.240 209.540 ;
        RECT 47.480 209.260 47.760 209.540 ;
        RECT 40.840 206.870 41.120 207.150 ;
        RECT 41.360 206.870 41.640 207.150 ;
        RECT 43.000 208.190 43.280 208.470 ;
        RECT 43.520 208.190 43.800 208.470 ;
        RECT 46.960 208.190 47.240 208.470 ;
        RECT 47.480 208.190 47.760 208.470 ;
        RECT 43.000 207.310 43.280 207.590 ;
        RECT 43.520 207.310 43.800 207.590 ;
        RECT 43.000 204.670 43.280 204.950 ;
        RECT 43.520 204.670 43.800 204.950 ;
        RECT 46.960 204.670 47.240 204.950 ;
        RECT 47.480 204.670 47.760 204.950 ;
        RECT 43.000 202.910 43.280 203.190 ;
        RECT 43.520 202.910 43.800 203.190 ;
        RECT 46.960 202.910 47.240 203.190 ;
        RECT 47.480 202.910 47.760 203.190 ;
        RECT 46.960 202.030 47.240 202.310 ;
        RECT 47.480 202.030 47.760 202.310 ;
        RECT 40.840 201.590 41.120 201.870 ;
        RECT 41.360 201.590 41.640 201.870 ;
        RECT 43.000 199.390 43.280 199.670 ;
        RECT 43.520 199.390 43.800 199.670 ;
        RECT 46.960 199.390 47.240 199.670 ;
        RECT 47.480 199.390 47.760 199.670 ;
        RECT 43.000 197.630 43.280 197.910 ;
        RECT 43.520 197.630 43.800 197.910 ;
        RECT 46.960 197.630 47.240 197.910 ;
        RECT 47.480 197.630 47.760 197.910 ;
        RECT 49.120 196.310 49.400 196.590 ;
        RECT 49.640 196.310 49.920 196.590 ;
        RECT 43.000 195.870 43.280 196.150 ;
        RECT 43.520 195.870 43.800 196.150 ;
        RECT 46.960 195.870 47.240 196.150 ;
        RECT 47.480 195.870 47.760 196.150 ;
        RECT 43.000 194.990 43.280 195.270 ;
        RECT 43.520 194.990 43.800 195.270 ;
        RECT 43.000 192.350 43.280 192.630 ;
        RECT 43.520 192.350 43.800 192.630 ;
        RECT 43.000 191.470 43.280 191.750 ;
        RECT 43.520 191.470 43.800 191.750 ;
        RECT 40.840 191.030 41.120 191.310 ;
        RECT 41.360 191.030 41.640 191.310 ;
        RECT 43.000 188.830 43.280 189.110 ;
        RECT 43.520 188.830 43.800 189.110 ;
        RECT 49.120 192.790 49.400 193.070 ;
        RECT 49.640 192.790 49.920 193.070 ;
        RECT 46.960 192.350 47.240 192.630 ;
        RECT 47.480 192.350 47.760 192.630 ;
        RECT 46.960 191.470 47.240 191.750 ;
        RECT 47.480 191.470 47.760 191.750 ;
        RECT 43.000 187.950 43.280 188.230 ;
        RECT 43.520 187.950 43.800 188.230 ;
        RECT 46.960 187.950 47.240 188.230 ;
        RECT 47.480 187.950 47.760 188.230 ;
        RECT 43.000 185.310 43.280 185.590 ;
        RECT 43.520 185.310 43.800 185.590 ;
        RECT 43.000 184.430 43.280 184.710 ;
        RECT 43.520 184.430 43.800 184.710 ;
        RECT 46.960 184.430 47.240 184.710 ;
        RECT 47.480 184.430 47.760 184.710 ;
        RECT 46.140 182.870 46.420 183.150 ;
        RECT 46.140 182.350 46.420 182.630 ;
        RECT 43.000 181.790 43.280 182.070 ;
        RECT 43.520 181.790 43.800 182.070 ;
        RECT 46.960 181.790 47.240 182.070 ;
        RECT 47.480 181.790 47.760 182.070 ;
        RECT 43.000 180.910 43.280 181.190 ;
        RECT 43.520 180.910 43.800 181.190 ;
        RECT 46.960 180.910 47.240 181.190 ;
        RECT 47.480 180.910 47.760 181.190 ;
        RECT 43.000 178.270 43.280 178.550 ;
        RECT 43.520 178.270 43.800 178.550 ;
        RECT 43.000 177.390 43.280 177.670 ;
        RECT 43.520 177.390 43.800 177.670 ;
        RECT 46.960 177.390 47.240 177.670 ;
        RECT 47.480 177.390 47.760 177.670 ;
        RECT 45.265 175.830 45.545 176.110 ;
        RECT 40.840 175.190 41.120 175.470 ;
        RECT 41.360 175.190 41.640 175.470 ;
        RECT 45.265 175.310 45.545 175.590 ;
        RECT 43.000 174.750 43.280 175.030 ;
        RECT 43.520 174.750 43.800 175.030 ;
        RECT 46.960 174.750 47.240 175.030 ;
        RECT 47.480 174.750 47.760 175.030 ;
        RECT 43.000 173.870 43.280 174.150 ;
        RECT 43.520 173.870 43.800 174.150 ;
        RECT 46.960 173.870 47.240 174.150 ;
        RECT 47.480 173.870 47.760 174.150 ;
        RECT 43.000 171.230 43.280 171.510 ;
        RECT 43.520 171.230 43.800 171.510 ;
        RECT 43.000 170.350 43.280 170.630 ;
        RECT 43.520 170.350 43.800 170.630 ;
        RECT 46.960 170.350 47.240 170.630 ;
        RECT 47.480 170.350 47.760 170.630 ;
        RECT 44.465 168.790 44.745 169.070 ;
        RECT 46.960 168.590 47.240 168.870 ;
        RECT 47.480 168.590 47.760 168.870 ;
        RECT 40.920 168.110 41.200 168.390 ;
        RECT 41.440 168.110 41.720 168.390 ;
        RECT 44.465 168.270 44.745 168.550 ;
        RECT 43.000 167.710 43.280 167.990 ;
        RECT 43.520 167.710 43.800 167.990 ;
        RECT 46.960 167.710 47.240 167.990 ;
        RECT 47.480 167.710 47.760 167.990 ;
        RECT 43.000 166.830 43.280 167.110 ;
        RECT 43.520 166.830 43.800 167.110 ;
        RECT 46.960 166.830 47.240 167.110 ;
        RECT 47.480 166.830 47.760 167.110 ;
        RECT 43.000 164.190 43.280 164.470 ;
        RECT 43.520 164.190 43.800 164.470 ;
        RECT 43.000 163.310 43.280 163.590 ;
        RECT 43.520 163.310 43.800 163.590 ;
        RECT 46.960 163.310 47.240 163.590 ;
        RECT 47.480 163.310 47.760 163.590 ;
        RECT 43.000 160.670 43.280 160.950 ;
        RECT 43.520 160.670 43.800 160.950 ;
        RECT 46.960 160.670 47.240 160.950 ;
        RECT 47.480 160.670 47.760 160.950 ;
        RECT 40.840 159.350 41.120 159.630 ;
        RECT 41.360 159.350 41.640 159.630 ;
        RECT 49.120 159.350 49.400 159.630 ;
        RECT 49.640 159.350 49.920 159.630 ;
        RECT 40.840 155.830 41.120 156.110 ;
        RECT 41.360 155.830 41.640 156.110 ;
        RECT 40.840 154.070 41.120 154.350 ;
        RECT 41.360 154.070 41.640 154.350 ;
        RECT 43.000 155.390 43.280 155.670 ;
        RECT 43.520 155.390 43.800 155.670 ;
        RECT 46.960 155.390 47.240 155.670 ;
        RECT 47.480 155.390 47.760 155.670 ;
        RECT 43.000 154.510 43.280 154.790 ;
        RECT 43.520 154.510 43.800 154.790 ;
        RECT 41.000 150.550 41.280 150.830 ;
        RECT 41.520 150.550 41.800 150.830 ;
        RECT 43.000 150.110 43.280 150.390 ;
        RECT 43.520 150.110 43.800 150.390 ;
        RECT 46.960 150.110 47.240 150.390 ;
        RECT 47.480 150.110 47.760 150.390 ;
        RECT 43.000 148.350 43.280 148.630 ;
        RECT 43.520 148.350 43.800 148.630 ;
        RECT 46.960 148.350 47.240 148.630 ;
        RECT 47.480 148.350 47.760 148.630 ;
        RECT 46.960 147.470 47.240 147.750 ;
        RECT 47.480 147.470 47.760 147.750 ;
        RECT 43.000 146.590 43.280 146.870 ;
        RECT 43.520 146.590 43.800 146.870 ;
        RECT 43.000 145.710 43.280 145.990 ;
        RECT 43.520 145.710 43.800 145.990 ;
        RECT 41.000 145.270 41.280 145.550 ;
        RECT 41.520 145.270 41.800 145.550 ;
        RECT 43.000 143.070 43.280 143.350 ;
        RECT 43.520 143.070 43.800 143.350 ;
        RECT 46.960 143.070 47.240 143.350 ;
        RECT 47.480 143.070 47.760 143.350 ;
        RECT 46.960 142.190 47.240 142.470 ;
        RECT 47.480 142.190 47.760 142.470 ;
        RECT 40.840 141.750 41.120 142.030 ;
        RECT 41.360 141.750 41.640 142.030 ;
        RECT 43.000 140.430 43.280 140.710 ;
        RECT 43.520 140.430 43.800 140.710 ;
        RECT 46.960 140.430 47.240 140.710 ;
        RECT 47.480 140.430 47.760 140.710 ;
        RECT 30.560 139.550 30.840 139.830 ;
        RECT 31.080 139.550 31.360 139.830 ;
        RECT 34.520 139.550 34.800 139.830 ;
        RECT 35.040 139.550 35.320 139.830 ;
        RECT 68.200 210.830 68.480 211.110 ;
        RECT 68.720 210.830 69.000 211.110 ;
        RECT 72.160 210.830 72.440 211.110 ;
        RECT 72.680 210.830 72.960 211.110 ;
        RECT 55.760 209.950 56.040 210.230 ;
        RECT 56.280 209.950 56.560 210.230 ;
        RECT 59.720 209.950 60.000 210.230 ;
        RECT 60.240 209.950 60.520 210.230 ;
        RECT 55.600 209.070 55.880 209.350 ;
        RECT 56.120 209.070 56.400 209.350 ;
        RECT 55.760 208.190 56.040 208.470 ;
        RECT 56.280 208.190 56.560 208.470 ;
        RECT 59.720 208.190 60.000 208.470 ;
        RECT 60.240 208.190 60.520 208.470 ;
        RECT 59.720 207.310 60.000 207.590 ;
        RECT 60.240 207.310 60.520 207.590 ;
        RECT 61.720 206.870 62.000 207.150 ;
        RECT 62.240 206.870 62.520 207.150 ;
        RECT 55.760 204.670 56.040 204.950 ;
        RECT 56.280 204.670 56.560 204.950 ;
        RECT 59.720 204.670 60.000 204.950 ;
        RECT 60.240 204.670 60.520 204.950 ;
        RECT 55.760 202.910 56.040 203.190 ;
        RECT 56.280 202.910 56.560 203.190 ;
        RECT 59.720 202.910 60.000 203.190 ;
        RECT 60.240 202.910 60.520 203.190 ;
        RECT 55.760 202.030 56.040 202.310 ;
        RECT 56.280 202.030 56.560 202.310 ;
        RECT 61.880 201.590 62.160 201.870 ;
        RECT 62.400 201.590 62.680 201.870 ;
        RECT 55.760 199.390 56.040 199.670 ;
        RECT 56.280 199.390 56.560 199.670 ;
        RECT 59.720 199.390 60.000 199.670 ;
        RECT 60.240 199.390 60.520 199.670 ;
        RECT 55.760 197.630 56.040 197.910 ;
        RECT 56.280 197.630 56.560 197.910 ;
        RECT 59.720 197.630 60.000 197.910 ;
        RECT 60.240 197.630 60.520 197.910 ;
        RECT 53.600 196.310 53.880 196.590 ;
        RECT 54.120 196.310 54.400 196.590 ;
        RECT 55.760 195.870 56.040 196.150 ;
        RECT 56.280 195.870 56.560 196.150 ;
        RECT 59.720 195.870 60.000 196.150 ;
        RECT 60.240 195.870 60.520 196.150 ;
        RECT 59.720 194.990 60.000 195.270 ;
        RECT 60.240 194.990 60.520 195.270 ;
        RECT 53.600 192.790 53.880 193.070 ;
        RECT 54.120 192.790 54.400 193.070 ;
        RECT 55.760 192.350 56.040 192.630 ;
        RECT 56.280 192.350 56.560 192.630 ;
        RECT 55.760 191.470 56.040 191.750 ;
        RECT 56.280 191.470 56.560 191.750 ;
        RECT 59.720 192.350 60.000 192.630 ;
        RECT 60.240 192.350 60.520 192.630 ;
        RECT 59.720 191.470 60.000 191.750 ;
        RECT 60.240 191.470 60.520 191.750 ;
        RECT 61.720 191.030 62.000 191.310 ;
        RECT 62.240 191.030 62.520 191.310 ;
        RECT 59.720 188.830 60.000 189.110 ;
        RECT 60.240 188.830 60.520 189.110 ;
        RECT 55.760 187.950 56.040 188.230 ;
        RECT 56.280 187.950 56.560 188.230 ;
        RECT 59.720 187.950 60.000 188.230 ;
        RECT 60.240 187.950 60.520 188.230 ;
        RECT 55.760 184.430 56.040 184.710 ;
        RECT 56.280 184.430 56.560 184.710 ;
        RECT 57.100 182.870 57.380 183.150 ;
        RECT 59.720 185.310 60.000 185.590 ;
        RECT 60.240 185.310 60.520 185.590 ;
        RECT 59.720 184.430 60.000 184.710 ;
        RECT 60.240 184.430 60.520 184.710 ;
        RECT 57.100 182.350 57.380 182.630 ;
        RECT 55.760 181.790 56.040 182.070 ;
        RECT 56.280 181.790 56.560 182.070 ;
        RECT 59.720 181.790 60.000 182.070 ;
        RECT 60.240 181.790 60.520 182.070 ;
        RECT 55.760 180.910 56.040 181.190 ;
        RECT 56.280 180.910 56.560 181.190 ;
        RECT 59.720 180.910 60.000 181.190 ;
        RECT 60.240 180.910 60.520 181.190 ;
        RECT 55.760 177.390 56.040 177.670 ;
        RECT 56.280 177.390 56.560 177.670 ;
        RECT 57.975 175.830 58.255 176.110 ;
        RECT 59.720 178.270 60.000 178.550 ;
        RECT 60.240 178.270 60.520 178.550 ;
        RECT 59.720 177.390 60.000 177.670 ;
        RECT 60.240 177.390 60.520 177.670 ;
        RECT 57.975 175.310 58.255 175.590 ;
        RECT 61.880 175.190 62.160 175.470 ;
        RECT 62.400 175.190 62.680 175.470 ;
        RECT 55.760 174.750 56.040 175.030 ;
        RECT 56.280 174.750 56.560 175.030 ;
        RECT 59.720 174.750 60.000 175.030 ;
        RECT 60.240 174.750 60.520 175.030 ;
        RECT 55.760 173.870 56.040 174.150 ;
        RECT 56.280 173.870 56.560 174.150 ;
        RECT 59.720 173.870 60.000 174.150 ;
        RECT 60.240 173.870 60.520 174.150 ;
        RECT 55.760 170.350 56.040 170.630 ;
        RECT 56.280 170.350 56.560 170.630 ;
        RECT 59.720 171.230 60.000 171.510 ;
        RECT 60.240 171.230 60.520 171.510 ;
        RECT 59.720 170.350 60.000 170.630 ;
        RECT 60.240 170.350 60.520 170.630 ;
        RECT 55.760 168.590 56.040 168.870 ;
        RECT 56.280 168.590 56.560 168.870 ;
        RECT 58.775 168.790 59.055 169.070 ;
        RECT 58.775 168.270 59.055 168.550 ;
        RECT 55.760 167.710 56.040 167.990 ;
        RECT 56.280 167.710 56.560 167.990 ;
        RECT 59.720 167.710 60.000 167.990 ;
        RECT 60.240 167.710 60.520 167.990 ;
        RECT 55.760 166.830 56.040 167.110 ;
        RECT 56.280 166.830 56.560 167.110 ;
        RECT 59.720 166.830 60.000 167.110 ;
        RECT 60.240 166.830 60.520 167.110 ;
        RECT 55.760 163.310 56.040 163.590 ;
        RECT 56.280 163.310 56.560 163.590 ;
        RECT 59.720 164.190 60.000 164.470 ;
        RECT 60.240 164.190 60.520 164.470 ;
        RECT 59.720 163.310 60.000 163.590 ;
        RECT 60.240 163.310 60.520 163.590 ;
        RECT 61.800 168.110 62.080 168.390 ;
        RECT 62.320 168.110 62.600 168.390 ;
        RECT 55.760 160.670 56.040 160.950 ;
        RECT 56.280 160.670 56.560 160.950 ;
        RECT 59.720 160.670 60.000 160.950 ;
        RECT 60.240 160.670 60.520 160.950 ;
        RECT 53.440 159.350 53.720 159.630 ;
        RECT 53.960 159.350 54.240 159.630 ;
        RECT 61.880 159.350 62.160 159.630 ;
        RECT 62.400 159.350 62.680 159.630 ;
        RECT 55.760 155.390 56.040 155.670 ;
        RECT 56.280 155.390 56.560 155.670 ;
        RECT 59.720 155.390 60.000 155.670 ;
        RECT 60.240 155.390 60.520 155.670 ;
        RECT 59.720 154.510 60.000 154.790 ;
        RECT 60.240 154.510 60.520 154.790 ;
        RECT 61.720 155.830 62.000 156.110 ;
        RECT 62.240 155.830 62.520 156.110 ;
        RECT 61.880 154.070 62.160 154.350 ;
        RECT 62.400 154.070 62.680 154.350 ;
        RECT 55.760 150.110 56.040 150.390 ;
        RECT 56.280 150.110 56.560 150.390 ;
        RECT 59.720 150.110 60.000 150.390 ;
        RECT 60.240 150.110 60.520 150.390 ;
        RECT 61.720 150.550 62.000 150.830 ;
        RECT 62.240 150.550 62.520 150.830 ;
        RECT 55.760 148.350 56.040 148.630 ;
        RECT 56.280 148.350 56.560 148.630 ;
        RECT 59.720 148.350 60.000 148.630 ;
        RECT 60.240 148.350 60.520 148.630 ;
        RECT 55.760 147.470 56.040 147.750 ;
        RECT 56.280 147.470 56.560 147.750 ;
        RECT 55.760 143.070 56.040 143.350 ;
        RECT 56.280 143.070 56.560 143.350 ;
        RECT 59.720 146.590 60.000 146.870 ;
        RECT 60.240 146.590 60.520 146.870 ;
        RECT 59.720 145.710 60.000 145.990 ;
        RECT 60.240 145.710 60.520 145.990 ;
        RECT 61.720 145.270 62.000 145.550 ;
        RECT 62.240 145.270 62.520 145.550 ;
        RECT 55.760 142.190 56.040 142.470 ;
        RECT 56.280 142.190 56.560 142.470 ;
        RECT 59.720 143.070 60.000 143.350 ;
        RECT 60.240 143.070 60.520 143.350 ;
        RECT 61.880 141.750 62.160 142.030 ;
        RECT 62.400 141.750 62.680 142.030 ;
        RECT 55.760 140.430 56.040 140.710 ;
        RECT 56.280 140.430 56.560 140.710 ;
        RECT 59.720 140.430 60.000 140.710 ;
        RECT 60.240 140.430 60.520 140.710 ;
        RECT 43.000 139.550 43.280 139.830 ;
        RECT 43.520 139.550 43.800 139.830 ;
        RECT 46.960 139.550 47.240 139.830 ;
        RECT 47.480 139.550 47.760 139.830 ;
        RECT 80.960 210.830 81.240 211.110 ;
        RECT 81.480 210.830 81.760 211.110 ;
        RECT 84.920 210.830 85.200 211.110 ;
        RECT 85.440 210.830 85.720 211.110 ;
        RECT 68.200 209.950 68.480 210.230 ;
        RECT 68.720 209.950 69.000 210.230 ;
        RECT 72.160 209.950 72.440 210.230 ;
        RECT 72.680 209.950 72.960 210.230 ;
        RECT 72.160 209.260 72.440 209.540 ;
        RECT 72.680 209.260 72.960 209.540 ;
        RECT 66.040 206.870 66.320 207.150 ;
        RECT 66.560 206.870 66.840 207.150 ;
        RECT 68.200 208.190 68.480 208.470 ;
        RECT 68.720 208.190 69.000 208.470 ;
        RECT 72.160 208.190 72.440 208.470 ;
        RECT 72.680 208.190 72.960 208.470 ;
        RECT 68.200 207.310 68.480 207.590 ;
        RECT 68.720 207.310 69.000 207.590 ;
        RECT 68.200 204.670 68.480 204.950 ;
        RECT 68.720 204.670 69.000 204.950 ;
        RECT 72.160 204.670 72.440 204.950 ;
        RECT 72.680 204.670 72.960 204.950 ;
        RECT 68.200 202.910 68.480 203.190 ;
        RECT 68.720 202.910 69.000 203.190 ;
        RECT 72.160 202.910 72.440 203.190 ;
        RECT 72.680 202.910 72.960 203.190 ;
        RECT 72.160 202.030 72.440 202.310 ;
        RECT 72.680 202.030 72.960 202.310 ;
        RECT 66.040 201.590 66.320 201.870 ;
        RECT 66.560 201.590 66.840 201.870 ;
        RECT 68.200 199.390 68.480 199.670 ;
        RECT 68.720 199.390 69.000 199.670 ;
        RECT 72.160 199.390 72.440 199.670 ;
        RECT 72.680 199.390 72.960 199.670 ;
        RECT 68.200 197.630 68.480 197.910 ;
        RECT 68.720 197.630 69.000 197.910 ;
        RECT 72.160 197.630 72.440 197.910 ;
        RECT 72.680 197.630 72.960 197.910 ;
        RECT 74.320 196.310 74.600 196.590 ;
        RECT 74.840 196.310 75.120 196.590 ;
        RECT 68.200 195.870 68.480 196.150 ;
        RECT 68.720 195.870 69.000 196.150 ;
        RECT 72.160 195.870 72.440 196.150 ;
        RECT 72.680 195.870 72.960 196.150 ;
        RECT 68.200 194.990 68.480 195.270 ;
        RECT 68.720 194.990 69.000 195.270 ;
        RECT 68.200 192.350 68.480 192.630 ;
        RECT 68.720 192.350 69.000 192.630 ;
        RECT 68.200 191.470 68.480 191.750 ;
        RECT 68.720 191.470 69.000 191.750 ;
        RECT 66.040 191.030 66.320 191.310 ;
        RECT 66.560 191.030 66.840 191.310 ;
        RECT 68.200 188.830 68.480 189.110 ;
        RECT 68.720 188.830 69.000 189.110 ;
        RECT 74.320 192.790 74.600 193.070 ;
        RECT 74.840 192.790 75.120 193.070 ;
        RECT 72.160 192.350 72.440 192.630 ;
        RECT 72.680 192.350 72.960 192.630 ;
        RECT 72.160 191.470 72.440 191.750 ;
        RECT 72.680 191.470 72.960 191.750 ;
        RECT 68.200 187.950 68.480 188.230 ;
        RECT 68.720 187.950 69.000 188.230 ;
        RECT 72.160 187.950 72.440 188.230 ;
        RECT 72.680 187.950 72.960 188.230 ;
        RECT 68.200 185.310 68.480 185.590 ;
        RECT 68.720 185.310 69.000 185.590 ;
        RECT 68.200 184.430 68.480 184.710 ;
        RECT 68.720 184.430 69.000 184.710 ;
        RECT 72.160 184.430 72.440 184.710 ;
        RECT 72.680 184.430 72.960 184.710 ;
        RECT 71.340 182.870 71.620 183.150 ;
        RECT 71.340 182.350 71.620 182.630 ;
        RECT 68.200 181.790 68.480 182.070 ;
        RECT 68.720 181.790 69.000 182.070 ;
        RECT 72.160 181.790 72.440 182.070 ;
        RECT 72.680 181.790 72.960 182.070 ;
        RECT 68.200 180.910 68.480 181.190 ;
        RECT 68.720 180.910 69.000 181.190 ;
        RECT 72.160 180.910 72.440 181.190 ;
        RECT 72.680 180.910 72.960 181.190 ;
        RECT 68.200 178.270 68.480 178.550 ;
        RECT 68.720 178.270 69.000 178.550 ;
        RECT 68.200 177.390 68.480 177.670 ;
        RECT 68.720 177.390 69.000 177.670 ;
        RECT 72.160 177.390 72.440 177.670 ;
        RECT 72.680 177.390 72.960 177.670 ;
        RECT 70.465 175.830 70.745 176.110 ;
        RECT 66.040 175.190 66.320 175.470 ;
        RECT 66.560 175.190 66.840 175.470 ;
        RECT 70.465 175.310 70.745 175.590 ;
        RECT 68.200 174.750 68.480 175.030 ;
        RECT 68.720 174.750 69.000 175.030 ;
        RECT 72.160 174.750 72.440 175.030 ;
        RECT 72.680 174.750 72.960 175.030 ;
        RECT 68.200 173.870 68.480 174.150 ;
        RECT 68.720 173.870 69.000 174.150 ;
        RECT 72.160 173.870 72.440 174.150 ;
        RECT 72.680 173.870 72.960 174.150 ;
        RECT 68.200 171.230 68.480 171.510 ;
        RECT 68.720 171.230 69.000 171.510 ;
        RECT 68.200 170.350 68.480 170.630 ;
        RECT 68.720 170.350 69.000 170.630 ;
        RECT 72.160 170.350 72.440 170.630 ;
        RECT 72.680 170.350 72.960 170.630 ;
        RECT 69.665 168.790 69.945 169.070 ;
        RECT 72.160 168.590 72.440 168.870 ;
        RECT 72.680 168.590 72.960 168.870 ;
        RECT 66.120 168.110 66.400 168.390 ;
        RECT 66.640 168.110 66.920 168.390 ;
        RECT 69.665 168.270 69.945 168.550 ;
        RECT 68.200 167.710 68.480 167.990 ;
        RECT 68.720 167.710 69.000 167.990 ;
        RECT 72.160 167.710 72.440 167.990 ;
        RECT 72.680 167.710 72.960 167.990 ;
        RECT 68.200 166.830 68.480 167.110 ;
        RECT 68.720 166.830 69.000 167.110 ;
        RECT 72.160 166.830 72.440 167.110 ;
        RECT 72.680 166.830 72.960 167.110 ;
        RECT 68.200 164.190 68.480 164.470 ;
        RECT 68.720 164.190 69.000 164.470 ;
        RECT 68.200 163.310 68.480 163.590 ;
        RECT 68.720 163.310 69.000 163.590 ;
        RECT 72.160 163.310 72.440 163.590 ;
        RECT 72.680 163.310 72.960 163.590 ;
        RECT 68.200 160.670 68.480 160.950 ;
        RECT 68.720 160.670 69.000 160.950 ;
        RECT 72.160 160.670 72.440 160.950 ;
        RECT 72.680 160.670 72.960 160.950 ;
        RECT 66.040 159.350 66.320 159.630 ;
        RECT 66.560 159.350 66.840 159.630 ;
        RECT 74.320 159.350 74.600 159.630 ;
        RECT 74.840 159.350 75.120 159.630 ;
        RECT 66.040 155.830 66.320 156.110 ;
        RECT 66.560 155.830 66.840 156.110 ;
        RECT 66.040 154.070 66.320 154.350 ;
        RECT 66.560 154.070 66.840 154.350 ;
        RECT 68.200 155.390 68.480 155.670 ;
        RECT 68.720 155.390 69.000 155.670 ;
        RECT 72.160 155.390 72.440 155.670 ;
        RECT 72.680 155.390 72.960 155.670 ;
        RECT 68.200 154.510 68.480 154.790 ;
        RECT 68.720 154.510 69.000 154.790 ;
        RECT 66.200 150.550 66.480 150.830 ;
        RECT 66.720 150.550 67.000 150.830 ;
        RECT 68.200 150.110 68.480 150.390 ;
        RECT 68.720 150.110 69.000 150.390 ;
        RECT 72.160 150.110 72.440 150.390 ;
        RECT 72.680 150.110 72.960 150.390 ;
        RECT 68.200 148.350 68.480 148.630 ;
        RECT 68.720 148.350 69.000 148.630 ;
        RECT 72.160 148.350 72.440 148.630 ;
        RECT 72.680 148.350 72.960 148.630 ;
        RECT 72.160 147.470 72.440 147.750 ;
        RECT 72.680 147.470 72.960 147.750 ;
        RECT 68.200 146.590 68.480 146.870 ;
        RECT 68.720 146.590 69.000 146.870 ;
        RECT 68.200 145.710 68.480 145.990 ;
        RECT 68.720 145.710 69.000 145.990 ;
        RECT 66.200 145.270 66.480 145.550 ;
        RECT 66.720 145.270 67.000 145.550 ;
        RECT 68.200 143.070 68.480 143.350 ;
        RECT 68.720 143.070 69.000 143.350 ;
        RECT 72.160 143.070 72.440 143.350 ;
        RECT 72.680 143.070 72.960 143.350 ;
        RECT 72.160 142.190 72.440 142.470 ;
        RECT 72.680 142.190 72.960 142.470 ;
        RECT 66.040 141.750 66.320 142.030 ;
        RECT 66.560 141.750 66.840 142.030 ;
        RECT 68.200 140.430 68.480 140.710 ;
        RECT 68.720 140.430 69.000 140.710 ;
        RECT 72.160 140.430 72.440 140.710 ;
        RECT 72.680 140.430 72.960 140.710 ;
        RECT 55.760 139.550 56.040 139.830 ;
        RECT 56.280 139.550 56.560 139.830 ;
        RECT 59.720 139.550 60.000 139.830 ;
        RECT 60.240 139.550 60.520 139.830 ;
        RECT 93.400 210.830 93.680 211.110 ;
        RECT 93.920 210.830 94.200 211.110 ;
        RECT 97.360 210.830 97.640 211.110 ;
        RECT 97.880 210.830 98.160 211.110 ;
        RECT 80.960 209.950 81.240 210.230 ;
        RECT 81.480 209.950 81.760 210.230 ;
        RECT 84.920 209.950 85.200 210.230 ;
        RECT 85.440 209.950 85.720 210.230 ;
        RECT 80.800 209.070 81.080 209.350 ;
        RECT 81.320 209.070 81.600 209.350 ;
        RECT 80.960 208.190 81.240 208.470 ;
        RECT 81.480 208.190 81.760 208.470 ;
        RECT 84.920 208.190 85.200 208.470 ;
        RECT 85.440 208.190 85.720 208.470 ;
        RECT 84.920 207.310 85.200 207.590 ;
        RECT 85.440 207.310 85.720 207.590 ;
        RECT 86.920 206.870 87.200 207.150 ;
        RECT 87.440 206.870 87.720 207.150 ;
        RECT 80.960 204.670 81.240 204.950 ;
        RECT 81.480 204.670 81.760 204.950 ;
        RECT 84.920 204.670 85.200 204.950 ;
        RECT 85.440 204.670 85.720 204.950 ;
        RECT 80.960 202.910 81.240 203.190 ;
        RECT 81.480 202.910 81.760 203.190 ;
        RECT 84.920 202.910 85.200 203.190 ;
        RECT 85.440 202.910 85.720 203.190 ;
        RECT 80.960 202.030 81.240 202.310 ;
        RECT 81.480 202.030 81.760 202.310 ;
        RECT 87.080 201.590 87.360 201.870 ;
        RECT 87.600 201.590 87.880 201.870 ;
        RECT 80.960 199.390 81.240 199.670 ;
        RECT 81.480 199.390 81.760 199.670 ;
        RECT 84.920 199.390 85.200 199.670 ;
        RECT 85.440 199.390 85.720 199.670 ;
        RECT 80.960 197.630 81.240 197.910 ;
        RECT 81.480 197.630 81.760 197.910 ;
        RECT 84.920 197.630 85.200 197.910 ;
        RECT 85.440 197.630 85.720 197.910 ;
        RECT 78.800 196.310 79.080 196.590 ;
        RECT 79.320 196.310 79.600 196.590 ;
        RECT 80.960 195.870 81.240 196.150 ;
        RECT 81.480 195.870 81.760 196.150 ;
        RECT 84.920 195.870 85.200 196.150 ;
        RECT 85.440 195.870 85.720 196.150 ;
        RECT 84.920 194.990 85.200 195.270 ;
        RECT 85.440 194.990 85.720 195.270 ;
        RECT 78.800 192.790 79.080 193.070 ;
        RECT 79.320 192.790 79.600 193.070 ;
        RECT 80.960 192.350 81.240 192.630 ;
        RECT 81.480 192.350 81.760 192.630 ;
        RECT 80.960 191.470 81.240 191.750 ;
        RECT 81.480 191.470 81.760 191.750 ;
        RECT 84.920 192.350 85.200 192.630 ;
        RECT 85.440 192.350 85.720 192.630 ;
        RECT 84.920 191.470 85.200 191.750 ;
        RECT 85.440 191.470 85.720 191.750 ;
        RECT 86.920 191.030 87.200 191.310 ;
        RECT 87.440 191.030 87.720 191.310 ;
        RECT 84.920 188.830 85.200 189.110 ;
        RECT 85.440 188.830 85.720 189.110 ;
        RECT 80.960 187.950 81.240 188.230 ;
        RECT 81.480 187.950 81.760 188.230 ;
        RECT 84.920 187.950 85.200 188.230 ;
        RECT 85.440 187.950 85.720 188.230 ;
        RECT 80.960 184.430 81.240 184.710 ;
        RECT 81.480 184.430 81.760 184.710 ;
        RECT 82.300 182.870 82.580 183.150 ;
        RECT 84.920 185.310 85.200 185.590 ;
        RECT 85.440 185.310 85.720 185.590 ;
        RECT 84.920 184.430 85.200 184.710 ;
        RECT 85.440 184.430 85.720 184.710 ;
        RECT 82.300 182.350 82.580 182.630 ;
        RECT 80.960 181.790 81.240 182.070 ;
        RECT 81.480 181.790 81.760 182.070 ;
        RECT 84.920 181.790 85.200 182.070 ;
        RECT 85.440 181.790 85.720 182.070 ;
        RECT 80.960 180.910 81.240 181.190 ;
        RECT 81.480 180.910 81.760 181.190 ;
        RECT 84.920 180.910 85.200 181.190 ;
        RECT 85.440 180.910 85.720 181.190 ;
        RECT 80.960 177.390 81.240 177.670 ;
        RECT 81.480 177.390 81.760 177.670 ;
        RECT 83.175 175.830 83.455 176.110 ;
        RECT 84.920 178.270 85.200 178.550 ;
        RECT 85.440 178.270 85.720 178.550 ;
        RECT 84.920 177.390 85.200 177.670 ;
        RECT 85.440 177.390 85.720 177.670 ;
        RECT 83.175 175.310 83.455 175.590 ;
        RECT 87.080 175.190 87.360 175.470 ;
        RECT 87.600 175.190 87.880 175.470 ;
        RECT 80.960 174.750 81.240 175.030 ;
        RECT 81.480 174.750 81.760 175.030 ;
        RECT 84.920 174.750 85.200 175.030 ;
        RECT 85.440 174.750 85.720 175.030 ;
        RECT 80.960 173.870 81.240 174.150 ;
        RECT 81.480 173.870 81.760 174.150 ;
        RECT 84.920 173.870 85.200 174.150 ;
        RECT 85.440 173.870 85.720 174.150 ;
        RECT 80.960 170.350 81.240 170.630 ;
        RECT 81.480 170.350 81.760 170.630 ;
        RECT 84.920 171.230 85.200 171.510 ;
        RECT 85.440 171.230 85.720 171.510 ;
        RECT 84.920 170.350 85.200 170.630 ;
        RECT 85.440 170.350 85.720 170.630 ;
        RECT 80.960 168.590 81.240 168.870 ;
        RECT 81.480 168.590 81.760 168.870 ;
        RECT 83.975 168.790 84.255 169.070 ;
        RECT 83.975 168.270 84.255 168.550 ;
        RECT 80.960 167.710 81.240 167.990 ;
        RECT 81.480 167.710 81.760 167.990 ;
        RECT 84.920 167.710 85.200 167.990 ;
        RECT 85.440 167.710 85.720 167.990 ;
        RECT 80.960 166.830 81.240 167.110 ;
        RECT 81.480 166.830 81.760 167.110 ;
        RECT 84.920 166.830 85.200 167.110 ;
        RECT 85.440 166.830 85.720 167.110 ;
        RECT 80.960 163.310 81.240 163.590 ;
        RECT 81.480 163.310 81.760 163.590 ;
        RECT 84.920 164.190 85.200 164.470 ;
        RECT 85.440 164.190 85.720 164.470 ;
        RECT 84.920 163.310 85.200 163.590 ;
        RECT 85.440 163.310 85.720 163.590 ;
        RECT 87.000 168.110 87.280 168.390 ;
        RECT 87.520 168.110 87.800 168.390 ;
        RECT 80.960 160.670 81.240 160.950 ;
        RECT 81.480 160.670 81.760 160.950 ;
        RECT 84.920 160.670 85.200 160.950 ;
        RECT 85.440 160.670 85.720 160.950 ;
        RECT 78.640 159.350 78.920 159.630 ;
        RECT 79.160 159.350 79.440 159.630 ;
        RECT 87.080 159.350 87.360 159.630 ;
        RECT 87.600 159.350 87.880 159.630 ;
        RECT 80.960 155.390 81.240 155.670 ;
        RECT 81.480 155.390 81.760 155.670 ;
        RECT 84.920 155.390 85.200 155.670 ;
        RECT 85.440 155.390 85.720 155.670 ;
        RECT 84.920 154.510 85.200 154.790 ;
        RECT 85.440 154.510 85.720 154.790 ;
        RECT 86.920 155.830 87.200 156.110 ;
        RECT 87.440 155.830 87.720 156.110 ;
        RECT 87.080 154.070 87.360 154.350 ;
        RECT 87.600 154.070 87.880 154.350 ;
        RECT 80.960 150.110 81.240 150.390 ;
        RECT 81.480 150.110 81.760 150.390 ;
        RECT 84.920 150.110 85.200 150.390 ;
        RECT 85.440 150.110 85.720 150.390 ;
        RECT 86.920 150.550 87.200 150.830 ;
        RECT 87.440 150.550 87.720 150.830 ;
        RECT 80.960 148.350 81.240 148.630 ;
        RECT 81.480 148.350 81.760 148.630 ;
        RECT 84.920 148.350 85.200 148.630 ;
        RECT 85.440 148.350 85.720 148.630 ;
        RECT 80.960 147.470 81.240 147.750 ;
        RECT 81.480 147.470 81.760 147.750 ;
        RECT 80.960 143.070 81.240 143.350 ;
        RECT 81.480 143.070 81.760 143.350 ;
        RECT 84.920 146.590 85.200 146.870 ;
        RECT 85.440 146.590 85.720 146.870 ;
        RECT 84.920 145.710 85.200 145.990 ;
        RECT 85.440 145.710 85.720 145.990 ;
        RECT 86.920 145.270 87.200 145.550 ;
        RECT 87.440 145.270 87.720 145.550 ;
        RECT 80.960 142.190 81.240 142.470 ;
        RECT 81.480 142.190 81.760 142.470 ;
        RECT 84.920 143.070 85.200 143.350 ;
        RECT 85.440 143.070 85.720 143.350 ;
        RECT 87.080 141.750 87.360 142.030 ;
        RECT 87.600 141.750 87.880 142.030 ;
        RECT 80.960 140.430 81.240 140.710 ;
        RECT 81.480 140.430 81.760 140.710 ;
        RECT 84.920 140.430 85.200 140.710 ;
        RECT 85.440 140.430 85.720 140.710 ;
        RECT 68.200 139.550 68.480 139.830 ;
        RECT 68.720 139.550 69.000 139.830 ;
        RECT 72.160 139.550 72.440 139.830 ;
        RECT 72.680 139.550 72.960 139.830 ;
        RECT 106.160 210.830 106.440 211.110 ;
        RECT 106.680 210.830 106.960 211.110 ;
        RECT 110.120 210.830 110.400 211.110 ;
        RECT 110.640 210.830 110.920 211.110 ;
        RECT 93.400 209.950 93.680 210.230 ;
        RECT 93.920 209.950 94.200 210.230 ;
        RECT 97.360 209.950 97.640 210.230 ;
        RECT 97.880 209.950 98.160 210.230 ;
        RECT 97.360 209.260 97.640 209.540 ;
        RECT 97.880 209.260 98.160 209.540 ;
        RECT 91.240 206.870 91.520 207.150 ;
        RECT 91.760 206.870 92.040 207.150 ;
        RECT 93.400 208.190 93.680 208.470 ;
        RECT 93.920 208.190 94.200 208.470 ;
        RECT 97.360 208.190 97.640 208.470 ;
        RECT 97.880 208.190 98.160 208.470 ;
        RECT 93.400 207.310 93.680 207.590 ;
        RECT 93.920 207.310 94.200 207.590 ;
        RECT 93.400 204.670 93.680 204.950 ;
        RECT 93.920 204.670 94.200 204.950 ;
        RECT 97.360 204.670 97.640 204.950 ;
        RECT 97.880 204.670 98.160 204.950 ;
        RECT 93.400 202.910 93.680 203.190 ;
        RECT 93.920 202.910 94.200 203.190 ;
        RECT 97.360 202.910 97.640 203.190 ;
        RECT 97.880 202.910 98.160 203.190 ;
        RECT 97.360 202.030 97.640 202.310 ;
        RECT 97.880 202.030 98.160 202.310 ;
        RECT 91.240 201.590 91.520 201.870 ;
        RECT 91.760 201.590 92.040 201.870 ;
        RECT 93.400 199.390 93.680 199.670 ;
        RECT 93.920 199.390 94.200 199.670 ;
        RECT 97.360 199.390 97.640 199.670 ;
        RECT 97.880 199.390 98.160 199.670 ;
        RECT 93.400 197.630 93.680 197.910 ;
        RECT 93.920 197.630 94.200 197.910 ;
        RECT 97.360 197.630 97.640 197.910 ;
        RECT 97.880 197.630 98.160 197.910 ;
        RECT 99.520 196.310 99.800 196.590 ;
        RECT 100.040 196.310 100.320 196.590 ;
        RECT 93.400 195.870 93.680 196.150 ;
        RECT 93.920 195.870 94.200 196.150 ;
        RECT 97.360 195.870 97.640 196.150 ;
        RECT 97.880 195.870 98.160 196.150 ;
        RECT 93.400 194.990 93.680 195.270 ;
        RECT 93.920 194.990 94.200 195.270 ;
        RECT 93.400 192.350 93.680 192.630 ;
        RECT 93.920 192.350 94.200 192.630 ;
        RECT 93.400 191.470 93.680 191.750 ;
        RECT 93.920 191.470 94.200 191.750 ;
        RECT 91.240 191.030 91.520 191.310 ;
        RECT 91.760 191.030 92.040 191.310 ;
        RECT 93.400 188.830 93.680 189.110 ;
        RECT 93.920 188.830 94.200 189.110 ;
        RECT 99.520 192.790 99.800 193.070 ;
        RECT 100.040 192.790 100.320 193.070 ;
        RECT 97.360 192.350 97.640 192.630 ;
        RECT 97.880 192.350 98.160 192.630 ;
        RECT 97.360 191.470 97.640 191.750 ;
        RECT 97.880 191.470 98.160 191.750 ;
        RECT 93.400 187.950 93.680 188.230 ;
        RECT 93.920 187.950 94.200 188.230 ;
        RECT 97.360 187.950 97.640 188.230 ;
        RECT 97.880 187.950 98.160 188.230 ;
        RECT 93.400 185.310 93.680 185.590 ;
        RECT 93.920 185.310 94.200 185.590 ;
        RECT 93.400 184.430 93.680 184.710 ;
        RECT 93.920 184.430 94.200 184.710 ;
        RECT 97.360 184.430 97.640 184.710 ;
        RECT 97.880 184.430 98.160 184.710 ;
        RECT 96.540 182.870 96.820 183.150 ;
        RECT 96.540 182.350 96.820 182.630 ;
        RECT 93.400 181.790 93.680 182.070 ;
        RECT 93.920 181.790 94.200 182.070 ;
        RECT 97.360 181.790 97.640 182.070 ;
        RECT 97.880 181.790 98.160 182.070 ;
        RECT 93.400 180.910 93.680 181.190 ;
        RECT 93.920 180.910 94.200 181.190 ;
        RECT 97.360 180.910 97.640 181.190 ;
        RECT 97.880 180.910 98.160 181.190 ;
        RECT 93.400 178.270 93.680 178.550 ;
        RECT 93.920 178.270 94.200 178.550 ;
        RECT 93.400 177.390 93.680 177.670 ;
        RECT 93.920 177.390 94.200 177.670 ;
        RECT 97.360 177.390 97.640 177.670 ;
        RECT 97.880 177.390 98.160 177.670 ;
        RECT 95.665 175.830 95.945 176.110 ;
        RECT 91.240 175.190 91.520 175.470 ;
        RECT 91.760 175.190 92.040 175.470 ;
        RECT 95.665 175.310 95.945 175.590 ;
        RECT 93.400 174.750 93.680 175.030 ;
        RECT 93.920 174.750 94.200 175.030 ;
        RECT 97.360 174.750 97.640 175.030 ;
        RECT 97.880 174.750 98.160 175.030 ;
        RECT 93.400 173.870 93.680 174.150 ;
        RECT 93.920 173.870 94.200 174.150 ;
        RECT 97.360 173.870 97.640 174.150 ;
        RECT 97.880 173.870 98.160 174.150 ;
        RECT 93.400 171.230 93.680 171.510 ;
        RECT 93.920 171.230 94.200 171.510 ;
        RECT 93.400 170.350 93.680 170.630 ;
        RECT 93.920 170.350 94.200 170.630 ;
        RECT 97.360 170.350 97.640 170.630 ;
        RECT 97.880 170.350 98.160 170.630 ;
        RECT 94.865 168.790 95.145 169.070 ;
        RECT 97.360 168.590 97.640 168.870 ;
        RECT 97.880 168.590 98.160 168.870 ;
        RECT 91.320 168.110 91.600 168.390 ;
        RECT 91.840 168.110 92.120 168.390 ;
        RECT 94.865 168.270 95.145 168.550 ;
        RECT 93.400 167.710 93.680 167.990 ;
        RECT 93.920 167.710 94.200 167.990 ;
        RECT 97.360 167.710 97.640 167.990 ;
        RECT 97.880 167.710 98.160 167.990 ;
        RECT 93.400 166.830 93.680 167.110 ;
        RECT 93.920 166.830 94.200 167.110 ;
        RECT 97.360 166.830 97.640 167.110 ;
        RECT 97.880 166.830 98.160 167.110 ;
        RECT 93.400 164.190 93.680 164.470 ;
        RECT 93.920 164.190 94.200 164.470 ;
        RECT 93.400 163.310 93.680 163.590 ;
        RECT 93.920 163.310 94.200 163.590 ;
        RECT 97.360 163.310 97.640 163.590 ;
        RECT 97.880 163.310 98.160 163.590 ;
        RECT 93.400 160.670 93.680 160.950 ;
        RECT 93.920 160.670 94.200 160.950 ;
        RECT 97.360 160.670 97.640 160.950 ;
        RECT 97.880 160.670 98.160 160.950 ;
        RECT 91.240 159.350 91.520 159.630 ;
        RECT 91.760 159.350 92.040 159.630 ;
        RECT 99.520 159.350 99.800 159.630 ;
        RECT 100.040 159.350 100.320 159.630 ;
        RECT 91.240 155.830 91.520 156.110 ;
        RECT 91.760 155.830 92.040 156.110 ;
        RECT 91.240 154.070 91.520 154.350 ;
        RECT 91.760 154.070 92.040 154.350 ;
        RECT 93.400 155.390 93.680 155.670 ;
        RECT 93.920 155.390 94.200 155.670 ;
        RECT 97.360 155.390 97.640 155.670 ;
        RECT 97.880 155.390 98.160 155.670 ;
        RECT 93.400 154.510 93.680 154.790 ;
        RECT 93.920 154.510 94.200 154.790 ;
        RECT 91.400 150.550 91.680 150.830 ;
        RECT 91.920 150.550 92.200 150.830 ;
        RECT 93.400 150.110 93.680 150.390 ;
        RECT 93.920 150.110 94.200 150.390 ;
        RECT 97.360 150.110 97.640 150.390 ;
        RECT 97.880 150.110 98.160 150.390 ;
        RECT 93.400 148.350 93.680 148.630 ;
        RECT 93.920 148.350 94.200 148.630 ;
        RECT 97.360 148.350 97.640 148.630 ;
        RECT 97.880 148.350 98.160 148.630 ;
        RECT 97.360 147.470 97.640 147.750 ;
        RECT 97.880 147.470 98.160 147.750 ;
        RECT 93.400 146.590 93.680 146.870 ;
        RECT 93.920 146.590 94.200 146.870 ;
        RECT 93.400 145.710 93.680 145.990 ;
        RECT 93.920 145.710 94.200 145.990 ;
        RECT 91.400 145.270 91.680 145.550 ;
        RECT 91.920 145.270 92.200 145.550 ;
        RECT 93.400 143.070 93.680 143.350 ;
        RECT 93.920 143.070 94.200 143.350 ;
        RECT 97.360 143.070 97.640 143.350 ;
        RECT 97.880 143.070 98.160 143.350 ;
        RECT 97.360 142.190 97.640 142.470 ;
        RECT 97.880 142.190 98.160 142.470 ;
        RECT 91.240 141.750 91.520 142.030 ;
        RECT 91.760 141.750 92.040 142.030 ;
        RECT 93.400 140.430 93.680 140.710 ;
        RECT 93.920 140.430 94.200 140.710 ;
        RECT 97.360 140.430 97.640 140.710 ;
        RECT 97.880 140.430 98.160 140.710 ;
        RECT 80.960 139.550 81.240 139.830 ;
        RECT 81.480 139.550 81.760 139.830 ;
        RECT 84.920 139.550 85.200 139.830 ;
        RECT 85.440 139.550 85.720 139.830 ;
        RECT 106.160 209.950 106.440 210.230 ;
        RECT 106.680 209.950 106.960 210.230 ;
        RECT 110.120 209.950 110.400 210.230 ;
        RECT 110.640 209.950 110.920 210.230 ;
        RECT 106.000 209.070 106.280 209.350 ;
        RECT 106.520 209.070 106.800 209.350 ;
        RECT 118.600 209.070 118.880 209.350 ;
        RECT 119.120 209.070 119.400 209.350 ;
        RECT 122.560 209.070 122.840 209.350 ;
        RECT 123.080 209.070 123.360 209.350 ;
        RECT 106.160 208.190 106.440 208.470 ;
        RECT 106.680 208.190 106.960 208.470 ;
        RECT 110.120 208.190 110.400 208.470 ;
        RECT 110.640 208.190 110.920 208.470 ;
        RECT 110.120 207.310 110.400 207.590 ;
        RECT 110.640 207.310 110.920 207.590 ;
        RECT 112.120 206.870 112.400 207.150 ;
        RECT 112.640 206.870 112.920 207.150 ;
        RECT 106.160 204.670 106.440 204.950 ;
        RECT 106.680 204.670 106.960 204.950 ;
        RECT 110.120 204.670 110.400 204.950 ;
        RECT 110.640 204.670 110.920 204.950 ;
        RECT 106.160 202.910 106.440 203.190 ;
        RECT 106.680 202.910 106.960 203.190 ;
        RECT 110.120 202.910 110.400 203.190 ;
        RECT 110.640 202.910 110.920 203.190 ;
        RECT 106.160 202.030 106.440 202.310 ;
        RECT 106.680 202.030 106.960 202.310 ;
        RECT 112.280 201.590 112.560 201.870 ;
        RECT 112.800 201.590 113.080 201.870 ;
        RECT 106.160 199.390 106.440 199.670 ;
        RECT 106.680 199.390 106.960 199.670 ;
        RECT 110.120 199.390 110.400 199.670 ;
        RECT 110.640 199.390 110.920 199.670 ;
        RECT 110.040 198.510 110.320 198.790 ;
        RECT 110.560 198.510 110.840 198.790 ;
        RECT 106.160 197.630 106.440 197.910 ;
        RECT 106.680 197.630 106.960 197.910 ;
        RECT 110.120 197.630 110.400 197.910 ;
        RECT 110.640 197.630 110.920 197.910 ;
        RECT 104.000 196.310 104.280 196.590 ;
        RECT 104.520 196.310 104.800 196.590 ;
        RECT 106.160 195.870 106.440 196.150 ;
        RECT 106.680 195.870 106.960 196.150 ;
        RECT 110.120 195.870 110.400 196.150 ;
        RECT 110.640 195.870 110.920 196.150 ;
        RECT 110.120 194.990 110.400 195.270 ;
        RECT 110.640 194.990 110.920 195.270 ;
        RECT 104.000 192.790 104.280 193.070 ;
        RECT 104.520 192.790 104.800 193.070 ;
        RECT 106.160 192.350 106.440 192.630 ;
        RECT 106.680 192.350 106.960 192.630 ;
        RECT 106.160 191.470 106.440 191.750 ;
        RECT 106.680 191.470 106.960 191.750 ;
        RECT 112.120 194.550 112.400 194.830 ;
        RECT 112.640 194.550 112.920 194.830 ;
        RECT 110.120 192.350 110.400 192.630 ;
        RECT 110.640 192.350 110.920 192.630 ;
        RECT 110.120 191.470 110.400 191.750 ;
        RECT 110.640 191.470 110.920 191.750 ;
        RECT 112.120 191.030 112.400 191.310 ;
        RECT 112.640 191.030 112.920 191.310 ;
        RECT 110.120 188.830 110.400 189.110 ;
        RECT 110.640 188.830 110.920 189.110 ;
        RECT 106.160 187.950 106.440 188.230 ;
        RECT 106.680 187.950 106.960 188.230 ;
        RECT 110.120 187.950 110.400 188.230 ;
        RECT 110.640 187.950 110.920 188.230 ;
        RECT 106.160 184.430 106.440 184.710 ;
        RECT 106.680 184.430 106.960 184.710 ;
        RECT 107.500 182.870 107.780 183.150 ;
        RECT 110.120 185.310 110.400 185.590 ;
        RECT 110.640 185.310 110.920 185.590 ;
        RECT 110.120 184.430 110.400 184.710 ;
        RECT 110.640 184.430 110.920 184.710 ;
        RECT 107.500 182.350 107.780 182.630 ;
        RECT 106.160 181.790 106.440 182.070 ;
        RECT 106.680 181.790 106.960 182.070 ;
        RECT 110.120 181.790 110.400 182.070 ;
        RECT 110.640 181.790 110.920 182.070 ;
        RECT 106.160 180.910 106.440 181.190 ;
        RECT 106.680 180.910 106.960 181.190 ;
        RECT 110.120 180.910 110.400 181.190 ;
        RECT 110.640 180.910 110.920 181.190 ;
        RECT 106.160 177.390 106.440 177.670 ;
        RECT 106.680 177.390 106.960 177.670 ;
        RECT 108.375 175.830 108.655 176.110 ;
        RECT 110.120 178.270 110.400 178.550 ;
        RECT 110.640 178.270 110.920 178.550 ;
        RECT 110.120 177.390 110.400 177.670 ;
        RECT 110.640 177.390 110.920 177.670 ;
        RECT 108.375 175.310 108.655 175.590 ;
        RECT 112.280 175.190 112.560 175.470 ;
        RECT 112.800 175.190 113.080 175.470 ;
        RECT 106.160 174.750 106.440 175.030 ;
        RECT 106.680 174.750 106.960 175.030 ;
        RECT 110.120 174.750 110.400 175.030 ;
        RECT 110.640 174.750 110.920 175.030 ;
        RECT 106.160 173.870 106.440 174.150 ;
        RECT 106.680 173.870 106.960 174.150 ;
        RECT 110.120 173.870 110.400 174.150 ;
        RECT 110.640 173.870 110.920 174.150 ;
        RECT 106.160 170.350 106.440 170.630 ;
        RECT 106.680 170.350 106.960 170.630 ;
        RECT 110.120 171.230 110.400 171.510 ;
        RECT 110.640 171.230 110.920 171.510 ;
        RECT 110.120 170.350 110.400 170.630 ;
        RECT 110.640 170.350 110.920 170.630 ;
        RECT 106.160 168.590 106.440 168.870 ;
        RECT 106.680 168.590 106.960 168.870 ;
        RECT 109.175 168.790 109.455 169.070 ;
        RECT 109.175 168.270 109.455 168.550 ;
        RECT 106.160 167.710 106.440 167.990 ;
        RECT 106.680 167.710 106.960 167.990 ;
        RECT 110.120 167.710 110.400 167.990 ;
        RECT 110.640 167.710 110.920 167.990 ;
        RECT 106.160 166.830 106.440 167.110 ;
        RECT 106.680 166.830 106.960 167.110 ;
        RECT 110.120 166.830 110.400 167.110 ;
        RECT 110.640 166.830 110.920 167.110 ;
        RECT 106.160 163.310 106.440 163.590 ;
        RECT 106.680 163.310 106.960 163.590 ;
        RECT 110.120 164.190 110.400 164.470 ;
        RECT 110.640 164.190 110.920 164.470 ;
        RECT 110.120 163.310 110.400 163.590 ;
        RECT 110.640 163.310 110.920 163.590 ;
        RECT 112.200 168.110 112.480 168.390 ;
        RECT 112.720 168.110 113.000 168.390 ;
        RECT 106.160 160.670 106.440 160.950 ;
        RECT 106.680 160.670 106.960 160.950 ;
        RECT 110.120 160.670 110.400 160.950 ;
        RECT 110.640 160.670 110.920 160.950 ;
        RECT 103.840 159.350 104.120 159.630 ;
        RECT 104.360 159.350 104.640 159.630 ;
        RECT 112.280 159.350 112.560 159.630 ;
        RECT 112.800 159.350 113.080 159.630 ;
        RECT 106.160 155.390 106.440 155.670 ;
        RECT 106.680 155.390 106.960 155.670 ;
        RECT 110.120 155.390 110.400 155.670 ;
        RECT 110.640 155.390 110.920 155.670 ;
        RECT 110.120 154.510 110.400 154.790 ;
        RECT 110.640 154.510 110.920 154.790 ;
        RECT 112.120 155.830 112.400 156.110 ;
        RECT 112.640 155.830 112.920 156.110 ;
        RECT 112.280 154.070 112.560 154.350 ;
        RECT 112.800 154.070 113.080 154.350 ;
        RECT 106.160 150.110 106.440 150.390 ;
        RECT 106.680 150.110 106.960 150.390 ;
        RECT 110.120 150.110 110.400 150.390 ;
        RECT 110.640 150.110 110.920 150.390 ;
        RECT 112.120 150.550 112.400 150.830 ;
        RECT 112.640 150.550 112.920 150.830 ;
        RECT 106.160 148.350 106.440 148.630 ;
        RECT 106.680 148.350 106.960 148.630 ;
        RECT 110.120 148.350 110.400 148.630 ;
        RECT 110.640 148.350 110.920 148.630 ;
        RECT 106.160 147.470 106.440 147.750 ;
        RECT 106.680 147.470 106.960 147.750 ;
        RECT 106.160 143.070 106.440 143.350 ;
        RECT 106.680 143.070 106.960 143.350 ;
        RECT 110.120 146.590 110.400 146.870 ;
        RECT 110.640 146.590 110.920 146.870 ;
        RECT 110.120 145.710 110.400 145.990 ;
        RECT 110.640 145.710 110.920 145.990 ;
        RECT 112.120 145.270 112.400 145.550 ;
        RECT 112.640 145.270 112.920 145.550 ;
        RECT 106.160 142.190 106.440 142.470 ;
        RECT 106.680 142.190 106.960 142.470 ;
        RECT 110.120 143.070 110.400 143.350 ;
        RECT 110.640 143.070 110.920 143.350 ;
        RECT 112.280 141.750 112.560 142.030 ;
        RECT 112.800 141.750 113.080 142.030 ;
        RECT 106.160 140.430 106.440 140.710 ;
        RECT 106.680 140.430 106.960 140.710 ;
        RECT 110.120 140.430 110.400 140.710 ;
        RECT 110.640 140.430 110.920 140.710 ;
        RECT 93.400 139.550 93.680 139.830 ;
        RECT 93.920 139.550 94.200 139.830 ;
        RECT 97.360 139.550 97.640 139.830 ;
        RECT 97.880 139.550 98.160 139.830 ;
        RECT 118.600 208.190 118.880 208.470 ;
        RECT 119.120 208.190 119.400 208.470 ;
        RECT 122.560 208.190 122.840 208.470 ;
        RECT 123.080 208.190 123.360 208.470 ;
        RECT 116.440 207.060 116.720 207.340 ;
        RECT 116.960 207.060 117.240 207.340 ;
        RECT 118.600 206.430 118.880 206.710 ;
        RECT 119.120 206.430 119.400 206.710 ;
        RECT 122.560 206.430 122.840 206.710 ;
        RECT 123.080 206.430 123.360 206.710 ;
        RECT 118.600 205.550 118.880 205.830 ;
        RECT 119.120 205.550 119.400 205.830 ;
        RECT 118.600 202.910 118.880 203.190 ;
        RECT 119.120 202.910 119.400 203.190 ;
        RECT 122.560 202.910 122.840 203.190 ;
        RECT 123.080 202.910 123.360 203.190 ;
        RECT 118.600 202.030 118.880 202.310 ;
        RECT 119.120 202.030 119.400 202.310 ;
        RECT 122.560 202.030 122.840 202.310 ;
        RECT 123.080 202.030 123.360 202.310 ;
        RECT 124.800 205.110 125.080 205.390 ;
        RECT 125.320 205.110 125.600 205.390 ;
        RECT 124.720 203.350 125.000 203.630 ;
        RECT 125.240 203.350 125.520 203.630 ;
        RECT 118.600 199.390 118.880 199.670 ;
        RECT 119.120 199.390 119.400 199.670 ;
        RECT 122.560 199.390 122.840 199.670 ;
        RECT 123.080 199.390 123.360 199.670 ;
        RECT 116.440 198.070 116.720 198.350 ;
        RECT 116.960 198.070 117.240 198.350 ;
        RECT 118.600 197.630 118.880 197.910 ;
        RECT 119.120 197.630 119.400 197.910 ;
        RECT 122.560 197.630 122.840 197.910 ;
        RECT 123.080 197.630 123.360 197.910 ;
        RECT 116.600 187.510 116.880 187.790 ;
        RECT 117.120 187.510 117.400 187.790 ;
        RECT 122.560 186.190 122.840 186.470 ;
        RECT 123.080 186.190 123.360 186.470 ;
        RECT 116.440 185.750 116.720 186.030 ;
        RECT 116.960 185.750 117.240 186.030 ;
        RECT 118.600 185.310 118.880 185.590 ;
        RECT 119.120 185.310 119.400 185.590 ;
        RECT 122.560 184.430 122.840 184.710 ;
        RECT 123.080 184.430 123.360 184.710 ;
        RECT 116.600 182.230 116.880 182.510 ;
        RECT 117.120 182.230 117.400 182.510 ;
        RECT 122.560 181.790 122.840 182.070 ;
        RECT 123.080 181.790 123.360 182.070 ;
        RECT 122.560 180.910 122.840 181.190 ;
        RECT 123.080 180.910 123.360 181.190 ;
        RECT 122.560 180.030 122.840 180.310 ;
        RECT 123.080 180.030 123.360 180.310 ;
        RECT 122.560 178.270 122.840 178.550 ;
        RECT 123.080 178.270 123.360 178.550 ;
        RECT 122.560 177.390 122.840 177.670 ;
        RECT 123.080 177.390 123.360 177.670 ;
        RECT 122.560 174.750 122.840 175.030 ;
        RECT 123.080 174.750 123.360 175.030 ;
        RECT 122.560 173.870 122.840 174.150 ;
        RECT 123.080 173.870 123.360 174.150 ;
        RECT 118.600 172.990 118.880 173.270 ;
        RECT 119.120 172.990 119.400 173.270 ;
        RECT 118.600 172.110 118.880 172.390 ;
        RECT 119.120 172.110 119.400 172.390 ;
        RECT 122.560 172.110 122.840 172.390 ;
        RECT 123.080 172.110 123.360 172.390 ;
        RECT 122.560 170.350 122.840 170.630 ;
        RECT 123.080 170.350 123.360 170.630 ;
        RECT 124.720 176.950 125.000 177.230 ;
        RECT 125.240 176.950 125.520 177.230 ;
        RECT 118.600 169.470 118.880 169.750 ;
        RECT 119.120 169.470 119.400 169.750 ;
        RECT 122.560 169.470 122.840 169.750 ;
        RECT 123.080 169.470 123.360 169.750 ;
        RECT 118.600 168.590 118.880 168.870 ;
        RECT 119.120 168.590 119.400 168.870 ;
        RECT 122.560 168.590 122.840 168.870 ;
        RECT 123.080 168.590 123.360 168.870 ;
        RECT 118.680 167.020 118.960 167.300 ;
        RECT 119.200 167.020 119.480 167.300 ;
        RECT 118.600 165.950 118.880 166.230 ;
        RECT 119.120 165.950 119.400 166.230 ;
        RECT 122.560 165.950 122.840 166.230 ;
        RECT 123.080 165.950 123.360 166.230 ;
        RECT 122.560 165.070 122.840 165.350 ;
        RECT 123.080 165.070 123.360 165.350 ;
        RECT 124.720 166.390 125.000 166.670 ;
        RECT 125.240 166.390 125.520 166.670 ;
        RECT 124.720 162.870 125.000 163.150 ;
        RECT 125.240 162.870 125.520 163.150 ;
        RECT 122.560 162.430 122.840 162.710 ;
        RECT 123.080 162.430 123.360 162.710 ;
        RECT 122.560 161.550 122.840 161.830 ;
        RECT 123.080 161.550 123.360 161.830 ;
        RECT 116.600 155.830 116.880 156.110 ;
        RECT 117.120 155.830 117.400 156.110 ;
        RECT 122.560 158.910 122.840 159.190 ;
        RECT 123.080 158.910 123.360 159.190 ;
        RECT 122.560 158.030 122.840 158.310 ;
        RECT 123.080 158.030 123.360 158.310 ;
        RECT 124.720 157.590 125.000 157.870 ;
        RECT 125.240 157.590 125.520 157.870 ;
        RECT 122.560 155.390 122.840 155.670 ;
        RECT 123.080 155.390 123.360 155.670 ;
        RECT 122.560 154.510 122.840 154.790 ;
        RECT 123.080 154.510 123.360 154.790 ;
        RECT 118.600 153.630 118.880 153.910 ;
        RECT 119.120 153.630 119.400 153.910 ;
        RECT 116.600 150.550 116.880 150.830 ;
        RECT 117.120 150.550 117.400 150.830 ;
        RECT 122.560 142.190 122.840 142.470 ;
        RECT 123.080 142.190 123.360 142.470 ;
        RECT 116.440 141.750 116.720 142.030 ;
        RECT 116.960 141.750 117.240 142.030 ;
        RECT 118.600 141.310 118.880 141.590 ;
        RECT 119.120 141.310 119.400 141.590 ;
        RECT 118.600 140.430 118.880 140.710 ;
        RECT 119.120 140.430 119.400 140.710 ;
        RECT 122.560 140.430 122.840 140.710 ;
        RECT 123.080 140.430 123.360 140.710 ;
        RECT 106.160 139.550 106.440 139.830 ;
        RECT 106.680 139.550 106.960 139.830 ;
        RECT 110.120 139.550 110.400 139.830 ;
        RECT 110.640 139.550 110.920 139.830 ;
        RECT 118.600 139.550 118.880 139.830 ;
        RECT 119.120 139.550 119.400 139.830 ;
        RECT 122.560 139.550 122.840 139.830 ;
        RECT 123.080 139.550 123.360 139.830 ;
        RECT 23.510 109.390 23.790 109.670 ;
        RECT 23.510 108.870 23.790 109.150 ;
        RECT 58.900 109.150 59.180 109.430 ;
        RECT 59.420 109.150 59.700 109.430 ;
        RECT 81.420 109.150 81.700 109.430 ;
        RECT 81.940 109.150 82.220 109.430 ;
        RECT 117.330 109.390 117.610 109.670 ;
        RECT 117.330 108.870 117.610 109.150 ;
        RECT 22.110 106.330 22.390 106.610 ;
        RECT 26.310 106.330 26.590 106.610 ;
        RECT 44.510 106.330 44.790 106.610 ;
        RECT 48.710 106.330 48.990 106.610 ;
        RECT 22.110 105.810 22.390 106.090 ;
        RECT 26.310 105.810 26.590 106.090 ;
        RECT 44.510 105.810 44.790 106.090 ;
        RECT 48.710 105.810 48.990 106.090 ;
        RECT 58.900 106.090 59.180 106.370 ;
        RECT 59.420 106.090 59.700 106.370 ;
        RECT 81.420 106.090 81.700 106.370 ;
        RECT 81.940 106.090 82.220 106.370 ;
        RECT 92.130 106.330 92.410 106.610 ;
        RECT 96.330 106.330 96.610 106.610 ;
        RECT 114.530 106.330 114.810 106.610 ;
        RECT 118.730 106.330 119.010 106.610 ;
        RECT 92.130 105.810 92.410 106.090 ;
        RECT 96.330 105.810 96.610 106.090 ;
        RECT 114.530 105.810 114.810 106.090 ;
        RECT 118.730 105.810 119.010 106.090 ;
        RECT 19.310 103.270 19.590 103.550 ;
        RECT 20.710 103.270 20.990 103.550 ;
        RECT 27.710 103.270 27.990 103.550 ;
        RECT 29.110 103.270 29.390 103.550 ;
        RECT 41.710 103.270 41.990 103.550 ;
        RECT 43.110 103.270 43.390 103.550 ;
        RECT 50.110 103.270 50.390 103.550 ;
        RECT 51.510 103.270 51.790 103.550 ;
        RECT 19.310 102.750 19.590 103.030 ;
        RECT 20.710 102.750 20.990 103.030 ;
        RECT 27.710 102.750 27.990 103.030 ;
        RECT 29.110 102.750 29.390 103.030 ;
        RECT 41.710 102.750 41.990 103.030 ;
        RECT 43.110 102.750 43.390 103.030 ;
        RECT 50.110 102.750 50.390 103.030 ;
        RECT 51.510 102.750 51.790 103.030 ;
        RECT 58.900 103.030 59.180 103.310 ;
        RECT 59.420 103.030 59.700 103.310 ;
        RECT 81.420 103.030 81.700 103.310 ;
        RECT 81.940 103.030 82.220 103.310 ;
        RECT 89.330 103.270 89.610 103.550 ;
        RECT 90.730 103.270 91.010 103.550 ;
        RECT 97.730 103.270 98.010 103.550 ;
        RECT 99.130 103.270 99.410 103.550 ;
        RECT 111.730 103.270 112.010 103.550 ;
        RECT 113.130 103.270 113.410 103.550 ;
        RECT 120.130 103.270 120.410 103.550 ;
        RECT 121.530 103.270 121.810 103.550 ;
        RECT 89.330 102.750 89.610 103.030 ;
        RECT 90.730 102.750 91.010 103.030 ;
        RECT 97.730 102.750 98.010 103.030 ;
        RECT 99.130 102.750 99.410 103.030 ;
        RECT 111.730 102.750 112.010 103.030 ;
        RECT 113.130 102.750 113.410 103.030 ;
        RECT 120.130 102.750 120.410 103.030 ;
        RECT 121.530 102.750 121.810 103.030 ;
        RECT 24.910 100.210 25.190 100.490 ;
        RECT 45.910 100.210 46.190 100.490 ;
        RECT 24.910 99.690 25.190 99.970 ;
        RECT 45.910 99.690 46.190 99.970 ;
        RECT 58.900 99.970 59.180 100.250 ;
        RECT 59.420 99.970 59.700 100.250 ;
        RECT 81.420 99.970 81.700 100.250 ;
        RECT 81.940 99.970 82.220 100.250 ;
        RECT 94.930 100.210 95.210 100.490 ;
        RECT 115.930 100.210 116.210 100.490 ;
        RECT 94.930 99.690 95.210 99.970 ;
        RECT 115.930 99.690 116.210 99.970 ;
        RECT 13.710 97.150 13.990 97.430 ;
        RECT 15.110 97.150 15.390 97.430 ;
        RECT 16.510 97.150 16.790 97.430 ;
        RECT 17.910 97.150 18.190 97.430 ;
        RECT 30.510 97.150 30.790 97.430 ;
        RECT 31.910 97.150 32.190 97.430 ;
        RECT 33.310 97.150 33.590 97.430 ;
        RECT 34.710 97.150 34.990 97.430 ;
        RECT 36.110 97.150 36.390 97.430 ;
        RECT 37.510 97.150 37.790 97.430 ;
        RECT 38.910 97.150 39.190 97.430 ;
        RECT 40.310 97.150 40.590 97.430 ;
        RECT 52.910 97.150 53.190 97.430 ;
        RECT 54.310 97.150 54.590 97.430 ;
        RECT 55.710 97.150 55.990 97.430 ;
        RECT 57.110 97.150 57.390 97.430 ;
        RECT 13.710 96.630 13.990 96.910 ;
        RECT 15.110 96.630 15.390 96.910 ;
        RECT 16.510 96.630 16.790 96.910 ;
        RECT 17.910 96.630 18.190 96.910 ;
        RECT 30.510 96.630 30.790 96.910 ;
        RECT 31.910 96.630 32.190 96.910 ;
        RECT 33.310 96.630 33.590 96.910 ;
        RECT 34.710 96.630 34.990 96.910 ;
        RECT 36.110 96.630 36.390 96.910 ;
        RECT 37.510 96.630 37.790 96.910 ;
        RECT 38.910 96.630 39.190 96.910 ;
        RECT 40.310 96.630 40.590 96.910 ;
        RECT 52.910 96.630 53.190 96.910 ;
        RECT 54.310 96.630 54.590 96.910 ;
        RECT 55.710 96.630 55.990 96.910 ;
        RECT 57.110 96.630 57.390 96.910 ;
        RECT 58.900 96.910 59.180 97.190 ;
        RECT 59.420 96.910 59.700 97.190 ;
        RECT 81.420 96.910 81.700 97.190 ;
        RECT 81.940 96.910 82.220 97.190 ;
        RECT 83.730 97.150 84.010 97.430 ;
        RECT 85.130 97.150 85.410 97.430 ;
        RECT 86.530 97.150 86.810 97.430 ;
        RECT 87.930 97.150 88.210 97.430 ;
        RECT 100.530 97.150 100.810 97.430 ;
        RECT 101.930 97.150 102.210 97.430 ;
        RECT 103.330 97.150 103.610 97.430 ;
        RECT 104.730 97.150 105.010 97.430 ;
        RECT 106.130 97.150 106.410 97.430 ;
        RECT 107.530 97.150 107.810 97.430 ;
        RECT 108.930 97.150 109.210 97.430 ;
        RECT 110.330 97.150 110.610 97.430 ;
        RECT 122.930 97.150 123.210 97.430 ;
        RECT 124.330 97.150 124.610 97.430 ;
        RECT 125.730 97.150 126.010 97.430 ;
        RECT 127.130 97.150 127.410 97.430 ;
        RECT 83.730 96.630 84.010 96.910 ;
        RECT 85.130 96.630 85.410 96.910 ;
        RECT 86.530 96.630 86.810 96.910 ;
        RECT 87.930 96.630 88.210 96.910 ;
        RECT 100.530 96.630 100.810 96.910 ;
        RECT 101.930 96.630 102.210 96.910 ;
        RECT 103.330 96.630 103.610 96.910 ;
        RECT 104.730 96.630 105.010 96.910 ;
        RECT 106.130 96.630 106.410 96.910 ;
        RECT 107.530 96.630 107.810 96.910 ;
        RECT 108.930 96.630 109.210 96.910 ;
        RECT 110.330 96.630 110.610 96.910 ;
        RECT 122.930 96.630 123.210 96.910 ;
        RECT 124.330 96.630 124.610 96.910 ;
        RECT 125.730 96.630 126.010 96.910 ;
        RECT 127.130 96.630 127.410 96.910 ;
        RECT 8.700 93.690 8.980 93.970 ;
        RECT 9.220 93.690 9.500 93.970 ;
        RECT 47.310 94.090 47.590 94.370 ;
        RECT 47.310 93.570 47.590 93.850 ;
        RECT 58.900 93.850 59.180 94.130 ;
        RECT 59.420 93.850 59.700 94.130 ;
        RECT 81.420 93.850 81.700 94.130 ;
        RECT 81.940 93.850 82.220 94.130 ;
        RECT 93.530 94.090 93.810 94.370 ;
        RECT 93.530 93.570 93.810 93.850 ;
        RECT 8.700 93.170 8.980 93.450 ;
        RECT 9.220 93.170 9.500 93.450 ;
        RECT 131.610 93.390 131.890 93.670 ;
        RECT 131.610 92.870 131.890 93.150 ;
        RECT 23.510 91.990 23.790 92.270 ;
        RECT 23.510 91.470 23.790 91.750 ;
        RECT 58.900 91.750 59.180 92.030 ;
        RECT 59.420 91.750 59.700 92.030 ;
        RECT 81.420 91.750 81.700 92.030 ;
        RECT 81.940 91.750 82.220 92.030 ;
        RECT 117.330 91.990 117.610 92.270 ;
        RECT 117.330 91.470 117.610 91.750 ;
        RECT 22.110 88.930 22.390 89.210 ;
        RECT 26.310 88.930 26.590 89.210 ;
        RECT 44.510 88.930 44.790 89.210 ;
        RECT 48.710 88.930 48.990 89.210 ;
        RECT 22.110 88.410 22.390 88.690 ;
        RECT 26.310 88.410 26.590 88.690 ;
        RECT 44.510 88.410 44.790 88.690 ;
        RECT 48.710 88.410 48.990 88.690 ;
        RECT 58.900 88.690 59.180 88.970 ;
        RECT 59.420 88.690 59.700 88.970 ;
        RECT 81.420 88.690 81.700 88.970 ;
        RECT 81.940 88.690 82.220 88.970 ;
        RECT 92.130 88.930 92.410 89.210 ;
        RECT 96.330 88.930 96.610 89.210 ;
        RECT 114.530 88.930 114.810 89.210 ;
        RECT 118.730 88.930 119.010 89.210 ;
        RECT 92.130 88.410 92.410 88.690 ;
        RECT 96.330 88.410 96.610 88.690 ;
        RECT 114.530 88.410 114.810 88.690 ;
        RECT 118.730 88.410 119.010 88.690 ;
        RECT 19.310 85.870 19.590 86.150 ;
        RECT 20.710 85.870 20.990 86.150 ;
        RECT 27.710 85.870 27.990 86.150 ;
        RECT 29.110 85.870 29.390 86.150 ;
        RECT 41.710 85.870 41.990 86.150 ;
        RECT 43.110 85.870 43.390 86.150 ;
        RECT 50.110 85.870 50.390 86.150 ;
        RECT 51.510 85.870 51.790 86.150 ;
        RECT 19.310 85.350 19.590 85.630 ;
        RECT 20.710 85.350 20.990 85.630 ;
        RECT 27.710 85.350 27.990 85.630 ;
        RECT 29.110 85.350 29.390 85.630 ;
        RECT 41.710 85.350 41.990 85.630 ;
        RECT 43.110 85.350 43.390 85.630 ;
        RECT 50.110 85.350 50.390 85.630 ;
        RECT 51.510 85.350 51.790 85.630 ;
        RECT 58.900 85.630 59.180 85.910 ;
        RECT 59.420 85.630 59.700 85.910 ;
        RECT 81.420 85.630 81.700 85.910 ;
        RECT 81.940 85.630 82.220 85.910 ;
        RECT 89.330 85.870 89.610 86.150 ;
        RECT 90.730 85.870 91.010 86.150 ;
        RECT 97.730 85.870 98.010 86.150 ;
        RECT 99.130 85.870 99.410 86.150 ;
        RECT 111.730 85.870 112.010 86.150 ;
        RECT 113.130 85.870 113.410 86.150 ;
        RECT 120.130 85.870 120.410 86.150 ;
        RECT 121.530 85.870 121.810 86.150 ;
        RECT 89.330 85.350 89.610 85.630 ;
        RECT 90.730 85.350 91.010 85.630 ;
        RECT 97.730 85.350 98.010 85.630 ;
        RECT 99.130 85.350 99.410 85.630 ;
        RECT 111.730 85.350 112.010 85.630 ;
        RECT 113.130 85.350 113.410 85.630 ;
        RECT 120.130 85.350 120.410 85.630 ;
        RECT 121.530 85.350 121.810 85.630 ;
        RECT 24.910 82.810 25.190 83.090 ;
        RECT 45.910 82.810 46.190 83.090 ;
        RECT 24.910 82.290 25.190 82.570 ;
        RECT 45.910 82.290 46.190 82.570 ;
        RECT 58.900 82.570 59.180 82.850 ;
        RECT 59.420 82.570 59.700 82.850 ;
        RECT 81.420 82.570 81.700 82.850 ;
        RECT 81.940 82.570 82.220 82.850 ;
        RECT 94.930 82.810 95.210 83.090 ;
        RECT 115.930 82.810 116.210 83.090 ;
        RECT 94.930 82.290 95.210 82.570 ;
        RECT 115.930 82.290 116.210 82.570 ;
        RECT 13.710 79.750 13.990 80.030 ;
        RECT 15.110 79.750 15.390 80.030 ;
        RECT 16.510 79.750 16.790 80.030 ;
        RECT 17.910 79.750 18.190 80.030 ;
        RECT 30.510 79.750 30.790 80.030 ;
        RECT 31.910 79.750 32.190 80.030 ;
        RECT 33.310 79.750 33.590 80.030 ;
        RECT 34.710 79.750 34.990 80.030 ;
        RECT 36.110 79.750 36.390 80.030 ;
        RECT 37.510 79.750 37.790 80.030 ;
        RECT 38.910 79.750 39.190 80.030 ;
        RECT 40.310 79.750 40.590 80.030 ;
        RECT 52.910 79.750 53.190 80.030 ;
        RECT 54.310 79.750 54.590 80.030 ;
        RECT 55.710 79.750 55.990 80.030 ;
        RECT 57.110 79.750 57.390 80.030 ;
        RECT 13.710 79.230 13.990 79.510 ;
        RECT 15.110 79.230 15.390 79.510 ;
        RECT 16.510 79.230 16.790 79.510 ;
        RECT 17.910 79.230 18.190 79.510 ;
        RECT 30.510 79.230 30.790 79.510 ;
        RECT 31.910 79.230 32.190 79.510 ;
        RECT 33.310 79.230 33.590 79.510 ;
        RECT 34.710 79.230 34.990 79.510 ;
        RECT 36.110 79.230 36.390 79.510 ;
        RECT 37.510 79.230 37.790 79.510 ;
        RECT 38.910 79.230 39.190 79.510 ;
        RECT 40.310 79.230 40.590 79.510 ;
        RECT 52.910 79.230 53.190 79.510 ;
        RECT 54.310 79.230 54.590 79.510 ;
        RECT 55.710 79.230 55.990 79.510 ;
        RECT 57.110 79.230 57.390 79.510 ;
        RECT 58.900 79.510 59.180 79.790 ;
        RECT 59.420 79.510 59.700 79.790 ;
        RECT 81.420 79.510 81.700 79.790 ;
        RECT 81.940 79.510 82.220 79.790 ;
        RECT 83.730 79.750 84.010 80.030 ;
        RECT 85.130 79.750 85.410 80.030 ;
        RECT 86.530 79.750 86.810 80.030 ;
        RECT 87.930 79.750 88.210 80.030 ;
        RECT 100.530 79.750 100.810 80.030 ;
        RECT 101.930 79.750 102.210 80.030 ;
        RECT 103.330 79.750 103.610 80.030 ;
        RECT 104.730 79.750 105.010 80.030 ;
        RECT 106.130 79.750 106.410 80.030 ;
        RECT 107.530 79.750 107.810 80.030 ;
        RECT 108.930 79.750 109.210 80.030 ;
        RECT 110.330 79.750 110.610 80.030 ;
        RECT 122.930 79.750 123.210 80.030 ;
        RECT 124.330 79.750 124.610 80.030 ;
        RECT 125.730 79.750 126.010 80.030 ;
        RECT 127.130 79.750 127.410 80.030 ;
        RECT 83.730 79.230 84.010 79.510 ;
        RECT 85.130 79.230 85.410 79.510 ;
        RECT 86.530 79.230 86.810 79.510 ;
        RECT 87.930 79.230 88.210 79.510 ;
        RECT 100.530 79.230 100.810 79.510 ;
        RECT 101.930 79.230 102.210 79.510 ;
        RECT 103.330 79.230 103.610 79.510 ;
        RECT 104.730 79.230 105.010 79.510 ;
        RECT 106.130 79.230 106.410 79.510 ;
        RECT 107.530 79.230 107.810 79.510 ;
        RECT 108.930 79.230 109.210 79.510 ;
        RECT 110.330 79.230 110.610 79.510 ;
        RECT 122.930 79.230 123.210 79.510 ;
        RECT 124.330 79.230 124.610 79.510 ;
        RECT 125.730 79.230 126.010 79.510 ;
        RECT 127.130 79.230 127.410 79.510 ;
        RECT 8.700 76.290 8.980 76.570 ;
        RECT 9.220 76.290 9.500 76.570 ;
        RECT 47.310 76.690 47.590 76.970 ;
        RECT 47.310 76.170 47.590 76.450 ;
        RECT 58.900 76.450 59.180 76.730 ;
        RECT 59.420 76.450 59.700 76.730 ;
        RECT 81.420 76.450 81.700 76.730 ;
        RECT 81.940 76.450 82.220 76.730 ;
        RECT 93.530 76.690 93.810 76.970 ;
        RECT 93.530 76.170 93.810 76.450 ;
        RECT 8.700 75.770 8.980 76.050 ;
        RECT 9.220 75.770 9.500 76.050 ;
        RECT 131.610 75.990 131.890 76.270 ;
        RECT 131.610 75.470 131.890 75.750 ;
        RECT 23.510 74.590 23.790 74.870 ;
        RECT 23.510 74.070 23.790 74.350 ;
        RECT 58.900 74.350 59.180 74.630 ;
        RECT 59.420 74.350 59.700 74.630 ;
        RECT 81.420 74.350 81.700 74.630 ;
        RECT 81.940 74.350 82.220 74.630 ;
        RECT 117.330 74.590 117.610 74.870 ;
        RECT 117.330 74.070 117.610 74.350 ;
        RECT 22.110 71.530 22.390 71.810 ;
        RECT 26.310 71.530 26.590 71.810 ;
        RECT 44.510 71.530 44.790 71.810 ;
        RECT 48.710 71.530 48.990 71.810 ;
        RECT 22.110 71.010 22.390 71.290 ;
        RECT 26.310 71.010 26.590 71.290 ;
        RECT 44.510 71.010 44.790 71.290 ;
        RECT 48.710 71.010 48.990 71.290 ;
        RECT 58.900 71.290 59.180 71.570 ;
        RECT 59.420 71.290 59.700 71.570 ;
        RECT 81.420 71.290 81.700 71.570 ;
        RECT 81.940 71.290 82.220 71.570 ;
        RECT 92.130 71.530 92.410 71.810 ;
        RECT 96.330 71.530 96.610 71.810 ;
        RECT 114.530 71.530 114.810 71.810 ;
        RECT 118.730 71.530 119.010 71.810 ;
        RECT 92.130 71.010 92.410 71.290 ;
        RECT 96.330 71.010 96.610 71.290 ;
        RECT 114.530 71.010 114.810 71.290 ;
        RECT 118.730 71.010 119.010 71.290 ;
        RECT 19.310 68.470 19.590 68.750 ;
        RECT 20.710 68.470 20.990 68.750 ;
        RECT 27.710 68.470 27.990 68.750 ;
        RECT 29.110 68.470 29.390 68.750 ;
        RECT 41.710 68.470 41.990 68.750 ;
        RECT 43.110 68.470 43.390 68.750 ;
        RECT 50.110 68.470 50.390 68.750 ;
        RECT 51.510 68.470 51.790 68.750 ;
        RECT 19.310 67.950 19.590 68.230 ;
        RECT 20.710 67.950 20.990 68.230 ;
        RECT 27.710 67.950 27.990 68.230 ;
        RECT 29.110 67.950 29.390 68.230 ;
        RECT 41.710 67.950 41.990 68.230 ;
        RECT 43.110 67.950 43.390 68.230 ;
        RECT 50.110 67.950 50.390 68.230 ;
        RECT 51.510 67.950 51.790 68.230 ;
        RECT 58.900 68.230 59.180 68.510 ;
        RECT 59.420 68.230 59.700 68.510 ;
        RECT 81.420 68.230 81.700 68.510 ;
        RECT 81.940 68.230 82.220 68.510 ;
        RECT 89.330 68.470 89.610 68.750 ;
        RECT 90.730 68.470 91.010 68.750 ;
        RECT 97.730 68.470 98.010 68.750 ;
        RECT 99.130 68.470 99.410 68.750 ;
        RECT 111.730 68.470 112.010 68.750 ;
        RECT 113.130 68.470 113.410 68.750 ;
        RECT 120.130 68.470 120.410 68.750 ;
        RECT 121.530 68.470 121.810 68.750 ;
        RECT 89.330 67.950 89.610 68.230 ;
        RECT 90.730 67.950 91.010 68.230 ;
        RECT 97.730 67.950 98.010 68.230 ;
        RECT 99.130 67.950 99.410 68.230 ;
        RECT 111.730 67.950 112.010 68.230 ;
        RECT 113.130 67.950 113.410 68.230 ;
        RECT 120.130 67.950 120.410 68.230 ;
        RECT 121.530 67.950 121.810 68.230 ;
        RECT 24.910 65.410 25.190 65.690 ;
        RECT 45.910 65.410 46.190 65.690 ;
        RECT 24.910 64.890 25.190 65.170 ;
        RECT 45.910 64.890 46.190 65.170 ;
        RECT 58.900 65.170 59.180 65.450 ;
        RECT 59.420 65.170 59.700 65.450 ;
        RECT 81.420 65.170 81.700 65.450 ;
        RECT 81.940 65.170 82.220 65.450 ;
        RECT 94.930 65.410 95.210 65.690 ;
        RECT 115.930 65.410 116.210 65.690 ;
        RECT 94.930 64.890 95.210 65.170 ;
        RECT 115.930 64.890 116.210 65.170 ;
        RECT 13.710 62.350 13.990 62.630 ;
        RECT 15.110 62.350 15.390 62.630 ;
        RECT 16.510 62.350 16.790 62.630 ;
        RECT 17.910 62.350 18.190 62.630 ;
        RECT 30.510 62.350 30.790 62.630 ;
        RECT 31.910 62.350 32.190 62.630 ;
        RECT 33.310 62.350 33.590 62.630 ;
        RECT 34.710 62.350 34.990 62.630 ;
        RECT 36.110 62.350 36.390 62.630 ;
        RECT 37.510 62.350 37.790 62.630 ;
        RECT 38.910 62.350 39.190 62.630 ;
        RECT 40.310 62.350 40.590 62.630 ;
        RECT 52.910 62.350 53.190 62.630 ;
        RECT 54.310 62.350 54.590 62.630 ;
        RECT 55.710 62.350 55.990 62.630 ;
        RECT 57.110 62.350 57.390 62.630 ;
        RECT 13.710 61.830 13.990 62.110 ;
        RECT 15.110 61.830 15.390 62.110 ;
        RECT 16.510 61.830 16.790 62.110 ;
        RECT 17.910 61.830 18.190 62.110 ;
        RECT 30.510 61.830 30.790 62.110 ;
        RECT 31.910 61.830 32.190 62.110 ;
        RECT 33.310 61.830 33.590 62.110 ;
        RECT 34.710 61.830 34.990 62.110 ;
        RECT 36.110 61.830 36.390 62.110 ;
        RECT 37.510 61.830 37.790 62.110 ;
        RECT 38.910 61.830 39.190 62.110 ;
        RECT 40.310 61.830 40.590 62.110 ;
        RECT 52.910 61.830 53.190 62.110 ;
        RECT 54.310 61.830 54.590 62.110 ;
        RECT 55.710 61.830 55.990 62.110 ;
        RECT 57.110 61.830 57.390 62.110 ;
        RECT 58.900 62.110 59.180 62.390 ;
        RECT 59.420 62.110 59.700 62.390 ;
        RECT 81.420 62.110 81.700 62.390 ;
        RECT 81.940 62.110 82.220 62.390 ;
        RECT 83.730 62.350 84.010 62.630 ;
        RECT 85.130 62.350 85.410 62.630 ;
        RECT 86.530 62.350 86.810 62.630 ;
        RECT 87.930 62.350 88.210 62.630 ;
        RECT 100.530 62.350 100.810 62.630 ;
        RECT 101.930 62.350 102.210 62.630 ;
        RECT 103.330 62.350 103.610 62.630 ;
        RECT 104.730 62.350 105.010 62.630 ;
        RECT 106.130 62.350 106.410 62.630 ;
        RECT 107.530 62.350 107.810 62.630 ;
        RECT 108.930 62.350 109.210 62.630 ;
        RECT 110.330 62.350 110.610 62.630 ;
        RECT 122.930 62.350 123.210 62.630 ;
        RECT 124.330 62.350 124.610 62.630 ;
        RECT 125.730 62.350 126.010 62.630 ;
        RECT 127.130 62.350 127.410 62.630 ;
        RECT 83.730 61.830 84.010 62.110 ;
        RECT 85.130 61.830 85.410 62.110 ;
        RECT 86.530 61.830 86.810 62.110 ;
        RECT 87.930 61.830 88.210 62.110 ;
        RECT 100.530 61.830 100.810 62.110 ;
        RECT 101.930 61.830 102.210 62.110 ;
        RECT 103.330 61.830 103.610 62.110 ;
        RECT 104.730 61.830 105.010 62.110 ;
        RECT 106.130 61.830 106.410 62.110 ;
        RECT 107.530 61.830 107.810 62.110 ;
        RECT 108.930 61.830 109.210 62.110 ;
        RECT 110.330 61.830 110.610 62.110 ;
        RECT 122.930 61.830 123.210 62.110 ;
        RECT 124.330 61.830 124.610 62.110 ;
        RECT 125.730 61.830 126.010 62.110 ;
        RECT 127.130 61.830 127.410 62.110 ;
        RECT 8.700 58.890 8.980 59.170 ;
        RECT 9.220 58.890 9.500 59.170 ;
        RECT 47.310 59.290 47.590 59.570 ;
        RECT 47.310 58.770 47.590 59.050 ;
        RECT 59.450 59.330 59.730 59.610 ;
        RECT 59.450 58.810 59.730 59.090 ;
        RECT 81.390 59.330 81.670 59.610 ;
        RECT 81.390 58.810 81.670 59.090 ;
        RECT 93.530 59.290 93.810 59.570 ;
        RECT 93.530 58.770 93.810 59.050 ;
        RECT 8.700 58.370 8.980 58.650 ;
        RECT 9.220 58.370 9.500 58.650 ;
        RECT 131.610 58.590 131.890 58.870 ;
        RECT 131.610 58.070 131.890 58.350 ;
        RECT 23.510 57.190 23.790 57.470 ;
        RECT 23.510 56.670 23.790 56.950 ;
        RECT 58.900 56.950 59.180 57.230 ;
        RECT 59.420 56.950 59.700 57.230 ;
        RECT 81.420 56.950 81.700 57.230 ;
        RECT 81.940 56.950 82.220 57.230 ;
        RECT 117.330 57.190 117.610 57.470 ;
        RECT 117.330 56.670 117.610 56.950 ;
        RECT 22.110 54.130 22.390 54.410 ;
        RECT 26.310 54.130 26.590 54.410 ;
        RECT 44.510 54.130 44.790 54.410 ;
        RECT 48.710 54.130 48.990 54.410 ;
        RECT 22.110 53.610 22.390 53.890 ;
        RECT 26.310 53.610 26.590 53.890 ;
        RECT 44.510 53.610 44.790 53.890 ;
        RECT 48.710 53.610 48.990 53.890 ;
        RECT 58.900 53.890 59.180 54.170 ;
        RECT 59.420 53.890 59.700 54.170 ;
        RECT 81.420 53.890 81.700 54.170 ;
        RECT 81.940 53.890 82.220 54.170 ;
        RECT 92.130 54.130 92.410 54.410 ;
        RECT 96.330 54.130 96.610 54.410 ;
        RECT 114.530 54.130 114.810 54.410 ;
        RECT 118.730 54.130 119.010 54.410 ;
        RECT 92.130 53.610 92.410 53.890 ;
        RECT 96.330 53.610 96.610 53.890 ;
        RECT 114.530 53.610 114.810 53.890 ;
        RECT 118.730 53.610 119.010 53.890 ;
        RECT 19.310 51.070 19.590 51.350 ;
        RECT 20.710 51.070 20.990 51.350 ;
        RECT 27.710 51.070 27.990 51.350 ;
        RECT 29.110 51.070 29.390 51.350 ;
        RECT 41.710 51.070 41.990 51.350 ;
        RECT 43.110 51.070 43.390 51.350 ;
        RECT 50.110 51.070 50.390 51.350 ;
        RECT 51.510 51.070 51.790 51.350 ;
        RECT 19.310 50.550 19.590 50.830 ;
        RECT 20.710 50.550 20.990 50.830 ;
        RECT 27.710 50.550 27.990 50.830 ;
        RECT 29.110 50.550 29.390 50.830 ;
        RECT 41.710 50.550 41.990 50.830 ;
        RECT 43.110 50.550 43.390 50.830 ;
        RECT 50.110 50.550 50.390 50.830 ;
        RECT 51.510 50.550 51.790 50.830 ;
        RECT 58.900 50.830 59.180 51.110 ;
        RECT 59.420 50.830 59.700 51.110 ;
        RECT 81.420 50.830 81.700 51.110 ;
        RECT 81.940 50.830 82.220 51.110 ;
        RECT 89.330 51.070 89.610 51.350 ;
        RECT 90.730 51.070 91.010 51.350 ;
        RECT 97.730 51.070 98.010 51.350 ;
        RECT 99.130 51.070 99.410 51.350 ;
        RECT 111.730 51.070 112.010 51.350 ;
        RECT 113.130 51.070 113.410 51.350 ;
        RECT 120.130 51.070 120.410 51.350 ;
        RECT 121.530 51.070 121.810 51.350 ;
        RECT 89.330 50.550 89.610 50.830 ;
        RECT 90.730 50.550 91.010 50.830 ;
        RECT 97.730 50.550 98.010 50.830 ;
        RECT 99.130 50.550 99.410 50.830 ;
        RECT 111.730 50.550 112.010 50.830 ;
        RECT 113.130 50.550 113.410 50.830 ;
        RECT 120.130 50.550 120.410 50.830 ;
        RECT 121.530 50.550 121.810 50.830 ;
        RECT 24.910 48.010 25.190 48.290 ;
        RECT 45.910 48.010 46.190 48.290 ;
        RECT 24.910 47.490 25.190 47.770 ;
        RECT 45.910 47.490 46.190 47.770 ;
        RECT 58.900 47.770 59.180 48.050 ;
        RECT 59.420 47.770 59.700 48.050 ;
        RECT 81.420 47.770 81.700 48.050 ;
        RECT 81.940 47.770 82.220 48.050 ;
        RECT 94.930 48.010 95.210 48.290 ;
        RECT 115.930 48.010 116.210 48.290 ;
        RECT 94.930 47.490 95.210 47.770 ;
        RECT 115.930 47.490 116.210 47.770 ;
        RECT 13.710 44.950 13.990 45.230 ;
        RECT 15.110 44.950 15.390 45.230 ;
        RECT 16.510 44.950 16.790 45.230 ;
        RECT 17.910 44.950 18.190 45.230 ;
        RECT 30.510 44.950 30.790 45.230 ;
        RECT 31.910 44.950 32.190 45.230 ;
        RECT 33.310 44.950 33.590 45.230 ;
        RECT 34.710 44.950 34.990 45.230 ;
        RECT 36.110 44.950 36.390 45.230 ;
        RECT 37.510 44.950 37.790 45.230 ;
        RECT 38.910 44.950 39.190 45.230 ;
        RECT 40.310 44.950 40.590 45.230 ;
        RECT 52.910 44.950 53.190 45.230 ;
        RECT 54.310 44.950 54.590 45.230 ;
        RECT 55.710 44.950 55.990 45.230 ;
        RECT 57.110 44.950 57.390 45.230 ;
        RECT 13.710 44.430 13.990 44.710 ;
        RECT 15.110 44.430 15.390 44.710 ;
        RECT 16.510 44.430 16.790 44.710 ;
        RECT 17.910 44.430 18.190 44.710 ;
        RECT 30.510 44.430 30.790 44.710 ;
        RECT 31.910 44.430 32.190 44.710 ;
        RECT 33.310 44.430 33.590 44.710 ;
        RECT 34.710 44.430 34.990 44.710 ;
        RECT 36.110 44.430 36.390 44.710 ;
        RECT 37.510 44.430 37.790 44.710 ;
        RECT 38.910 44.430 39.190 44.710 ;
        RECT 40.310 44.430 40.590 44.710 ;
        RECT 52.910 44.430 53.190 44.710 ;
        RECT 54.310 44.430 54.590 44.710 ;
        RECT 55.710 44.430 55.990 44.710 ;
        RECT 57.110 44.430 57.390 44.710 ;
        RECT 58.900 44.710 59.180 44.990 ;
        RECT 59.420 44.710 59.700 44.990 ;
        RECT 81.420 44.710 81.700 44.990 ;
        RECT 81.940 44.710 82.220 44.990 ;
        RECT 83.730 44.950 84.010 45.230 ;
        RECT 85.130 44.950 85.410 45.230 ;
        RECT 86.530 44.950 86.810 45.230 ;
        RECT 87.930 44.950 88.210 45.230 ;
        RECT 100.530 44.950 100.810 45.230 ;
        RECT 101.930 44.950 102.210 45.230 ;
        RECT 103.330 44.950 103.610 45.230 ;
        RECT 104.730 44.950 105.010 45.230 ;
        RECT 106.130 44.950 106.410 45.230 ;
        RECT 107.530 44.950 107.810 45.230 ;
        RECT 108.930 44.950 109.210 45.230 ;
        RECT 110.330 44.950 110.610 45.230 ;
        RECT 122.930 44.950 123.210 45.230 ;
        RECT 124.330 44.950 124.610 45.230 ;
        RECT 125.730 44.950 126.010 45.230 ;
        RECT 127.130 44.950 127.410 45.230 ;
        RECT 83.730 44.430 84.010 44.710 ;
        RECT 85.130 44.430 85.410 44.710 ;
        RECT 86.530 44.430 86.810 44.710 ;
        RECT 87.930 44.430 88.210 44.710 ;
        RECT 100.530 44.430 100.810 44.710 ;
        RECT 101.930 44.430 102.210 44.710 ;
        RECT 103.330 44.430 103.610 44.710 ;
        RECT 104.730 44.430 105.010 44.710 ;
        RECT 106.130 44.430 106.410 44.710 ;
        RECT 107.530 44.430 107.810 44.710 ;
        RECT 108.930 44.430 109.210 44.710 ;
        RECT 110.330 44.430 110.610 44.710 ;
        RECT 122.930 44.430 123.210 44.710 ;
        RECT 124.330 44.430 124.610 44.710 ;
        RECT 125.730 44.430 126.010 44.710 ;
        RECT 127.130 44.430 127.410 44.710 ;
        RECT 8.700 41.490 8.980 41.770 ;
        RECT 9.220 41.490 9.500 41.770 ;
        RECT 47.310 41.890 47.590 42.170 ;
        RECT 47.310 41.370 47.590 41.650 ;
        RECT 58.900 41.650 59.180 41.930 ;
        RECT 59.420 41.650 59.700 41.930 ;
        RECT 81.420 41.650 81.700 41.930 ;
        RECT 81.940 41.650 82.220 41.930 ;
        RECT 93.530 41.890 93.810 42.170 ;
        RECT 93.530 41.370 93.810 41.650 ;
        RECT 8.700 40.970 8.980 41.250 ;
        RECT 9.220 40.970 9.500 41.250 ;
        RECT 131.610 41.190 131.890 41.470 ;
        RECT 131.610 40.670 131.890 40.950 ;
        RECT 47.080 38.580 48.160 38.935 ;
        RECT 14.320 37.700 15.400 38.055 ;
        RECT 47.080 36.820 48.160 37.175 ;
        RECT 14.320 35.940 15.400 36.295 ;
        RECT 47.080 35.060 48.160 35.415 ;
        RECT 93.160 38.580 94.240 38.935 ;
        RECT 125.920 37.700 127.000 38.055 ;
        RECT 93.160 36.820 94.240 37.175 ;
        RECT 125.920 35.940 127.000 36.295 ;
        RECT 93.160 35.060 94.240 35.415 ;
        RECT 14.320 34.185 15.400 34.535 ;
        RECT 125.920 34.185 127.000 34.535 ;
        RECT 47.080 33.300 48.160 33.655 ;
        RECT 14.320 32.420 15.400 32.775 ;
        RECT 93.160 33.300 94.240 33.655 ;
        RECT 47.080 31.540 48.160 31.895 ;
        RECT 14.320 30.660 15.400 31.015 ;
        RECT 47.080 29.780 48.160 30.135 ;
        RECT 54.860 32.040 55.140 32.320 ;
        RECT 55.380 32.040 55.660 32.320 ;
        RECT 58.820 32.040 59.100 32.320 ;
        RECT 59.340 32.040 59.620 32.320 ;
        RECT 14.320 28.905 15.400 29.255 ;
        RECT 47.080 28.020 48.160 28.375 ;
        RECT 14.320 27.140 15.400 27.495 ;
        RECT 47.080 26.260 48.160 26.615 ;
        RECT 14.320 25.380 15.400 25.735 ;
        RECT 47.080 24.500 48.160 24.855 ;
        RECT 54.860 31.160 55.140 31.440 ;
        RECT 55.380 31.160 55.660 31.440 ;
        RECT 58.820 31.160 59.100 31.440 ;
        RECT 59.340 31.160 59.620 31.440 ;
        RECT 58.820 30.280 59.100 30.560 ;
        RECT 59.340 30.280 59.620 30.560 ;
        RECT 54.860 29.400 55.140 29.680 ;
        RECT 55.380 29.400 55.660 29.680 ;
        RECT 58.820 29.400 59.100 29.680 ;
        RECT 59.340 29.400 59.620 29.680 ;
        RECT 54.860 28.520 55.140 28.800 ;
        RECT 55.380 28.520 55.660 28.800 ;
        RECT 58.820 28.520 59.100 28.800 ;
        RECT 59.340 28.520 59.620 28.800 ;
        RECT 14.320 23.625 15.400 23.975 ;
        RECT 47.080 22.740 48.160 23.095 ;
        RECT 14.320 21.860 15.400 22.215 ;
        RECT 47.080 20.980 48.160 21.335 ;
        RECT 14.320 20.100 15.400 20.455 ;
        RECT 47.080 19.220 48.160 19.575 ;
        RECT 14.320 18.345 15.400 18.695 ;
        RECT 47.080 17.460 48.160 17.815 ;
        RECT 14.320 16.580 15.400 16.935 ;
        RECT 47.080 15.700 48.160 16.055 ;
        RECT 14.320 14.820 15.400 15.175 ;
        RECT 47.080 13.940 48.160 14.295 ;
        RECT 54.860 27.640 55.140 27.920 ;
        RECT 55.380 27.640 55.660 27.920 ;
        RECT 58.820 27.640 59.100 27.920 ;
        RECT 59.340 27.640 59.620 27.920 ;
        RECT 54.860 26.930 55.140 27.210 ;
        RECT 55.380 26.930 55.660 27.210 ;
        RECT 54.860 25.880 55.140 26.160 ;
        RECT 55.380 25.880 55.660 26.160 ;
        RECT 58.820 25.880 59.100 26.160 ;
        RECT 59.340 25.880 59.620 26.160 ;
        RECT 54.860 25.000 55.140 25.280 ;
        RECT 55.380 25.000 55.660 25.280 ;
        RECT 58.740 25.000 59.020 25.280 ;
        RECT 59.260 25.000 59.540 25.280 ;
        RECT 54.860 23.240 55.140 23.520 ;
        RECT 55.380 23.240 55.660 23.520 ;
        RECT 60.980 24.560 61.260 24.840 ;
        RECT 61.500 24.560 61.780 24.840 ;
        RECT 60.980 22.800 61.260 23.080 ;
        RECT 61.500 22.800 61.780 23.080 ;
        RECT 58.820 22.360 59.100 22.640 ;
        RECT 59.340 22.360 59.620 22.640 ;
        RECT 58.820 21.480 59.100 21.760 ;
        RECT 59.340 21.480 59.620 21.760 ;
        RECT 54.860 20.600 55.140 20.880 ;
        RECT 55.380 20.600 55.660 20.880 ;
        RECT 52.700 19.280 52.980 19.560 ;
        RECT 53.220 19.280 53.500 19.560 ;
        RECT 54.860 18.840 55.140 19.120 ;
        RECT 55.380 18.840 55.660 19.120 ;
        RECT 58.820 18.840 59.100 19.120 ;
        RECT 59.340 18.840 59.620 19.120 ;
        RECT 54.860 17.960 55.140 18.240 ;
        RECT 55.380 17.960 55.660 18.240 ;
        RECT 58.820 17.960 59.100 18.240 ;
        RECT 59.340 17.960 59.620 18.240 ;
        RECT 52.700 17.520 52.980 17.800 ;
        RECT 53.220 17.520 53.500 17.800 ;
        RECT 54.860 16.200 55.140 16.480 ;
        RECT 55.380 16.200 55.660 16.480 ;
        RECT 58.820 16.390 59.100 16.670 ;
        RECT 59.340 16.390 59.620 16.670 ;
        RECT 60.900 15.760 61.180 16.040 ;
        RECT 61.420 15.760 61.700 16.040 ;
        RECT 54.860 15.320 55.140 15.600 ;
        RECT 55.380 15.320 55.660 15.600 ;
        RECT 58.820 15.320 59.100 15.600 ;
        RECT 59.340 15.320 59.620 15.600 ;
        RECT 54.860 14.440 55.140 14.720 ;
        RECT 55.380 14.440 55.660 14.720 ;
        RECT 58.820 14.440 59.100 14.720 ;
        RECT 59.340 14.440 59.620 14.720 ;
        RECT 14.320 13.065 15.400 13.415 ;
        RECT 81.700 32.040 81.980 32.320 ;
        RECT 82.220 32.040 82.500 32.320 ;
        RECT 85.660 32.040 85.940 32.320 ;
        RECT 86.180 32.040 86.460 32.320 ;
        RECT 81.700 31.160 81.980 31.440 ;
        RECT 82.220 31.160 82.500 31.440 ;
        RECT 85.660 31.160 85.940 31.440 ;
        RECT 86.180 31.160 86.460 31.440 ;
        RECT 81.700 30.280 81.980 30.560 ;
        RECT 82.220 30.280 82.500 30.560 ;
        RECT 81.700 29.400 81.980 29.680 ;
        RECT 82.220 29.400 82.500 29.680 ;
        RECT 85.660 29.400 85.940 29.680 ;
        RECT 86.180 29.400 86.460 29.680 ;
        RECT 81.700 28.520 81.980 28.800 ;
        RECT 82.220 28.520 82.500 28.800 ;
        RECT 85.660 28.520 85.940 28.800 ;
        RECT 86.180 28.520 86.460 28.800 ;
        RECT 65.860 25.880 66.140 26.160 ;
        RECT 66.380 25.880 66.660 26.160 ;
        RECT 68.180 26.320 68.460 26.600 ;
        RECT 68.700 26.320 68.980 26.600 ;
        RECT 54.860 13.560 55.140 13.840 ;
        RECT 55.380 13.560 55.660 13.840 ;
        RECT 58.820 13.560 59.100 13.840 ;
        RECT 59.340 13.560 59.620 13.840 ;
        RECT 65.860 18.840 66.140 19.120 ;
        RECT 66.380 18.840 66.660 19.120 ;
        RECT 66.020 17.960 66.300 18.240 ;
        RECT 66.540 17.960 66.820 18.240 ;
        RECT 68.100 17.520 68.380 17.800 ;
        RECT 68.620 17.520 68.900 17.800 ;
        RECT 65.940 14.400 66.220 14.680 ;
        RECT 66.460 14.400 66.740 14.680 ;
        RECT 72.340 26.320 72.620 26.600 ;
        RECT 72.860 26.320 73.140 26.600 ;
        RECT 74.500 25.880 74.780 26.160 ;
        RECT 75.020 25.880 75.300 26.160 ;
        RECT 74.500 18.840 74.780 19.120 ;
        RECT 75.020 18.840 75.300 19.120 ;
        RECT 74.500 17.960 74.780 18.240 ;
        RECT 75.020 17.960 75.300 18.240 ;
        RECT 72.420 17.520 72.700 17.800 ;
        RECT 72.940 17.520 73.220 17.800 ;
        RECT 74.580 14.400 74.860 14.680 ;
        RECT 75.100 14.400 75.380 14.680 ;
        RECT 125.920 32.420 127.000 32.775 ;
        RECT 93.160 31.540 94.240 31.895 ;
        RECT 125.920 30.660 127.000 31.015 ;
        RECT 93.160 29.780 94.240 30.135 ;
        RECT 125.920 28.905 127.000 29.255 ;
        RECT 81.700 27.640 81.980 27.920 ;
        RECT 82.220 27.640 82.500 27.920 ;
        RECT 85.660 27.640 85.940 27.920 ;
        RECT 86.180 27.640 86.460 27.920 ;
        RECT 85.660 26.930 85.940 27.210 ;
        RECT 86.180 26.930 86.460 27.210 ;
        RECT 81.700 25.880 81.980 26.160 ;
        RECT 82.220 25.880 82.500 26.160 ;
        RECT 85.660 25.880 85.940 26.160 ;
        RECT 86.180 25.880 86.460 26.160 ;
        RECT 81.780 25.000 82.060 25.280 ;
        RECT 82.300 25.000 82.580 25.280 ;
        RECT 85.660 25.000 85.940 25.280 ;
        RECT 86.180 25.000 86.460 25.280 ;
        RECT 79.540 24.560 79.820 24.840 ;
        RECT 80.060 24.560 80.340 24.840 ;
        RECT 79.540 22.800 79.820 23.080 ;
        RECT 80.060 22.800 80.340 23.080 ;
        RECT 81.700 22.360 81.980 22.640 ;
        RECT 82.220 22.360 82.500 22.640 ;
        RECT 85.660 23.240 85.940 23.520 ;
        RECT 86.180 23.240 86.460 23.520 ;
        RECT 81.700 21.480 81.980 21.760 ;
        RECT 82.220 21.480 82.500 21.760 ;
        RECT 85.660 20.600 85.940 20.880 ;
        RECT 86.180 20.600 86.460 20.880 ;
        RECT 87.820 19.280 88.100 19.560 ;
        RECT 88.340 19.280 88.620 19.560 ;
        RECT 81.700 18.840 81.980 19.120 ;
        RECT 82.220 18.840 82.500 19.120 ;
        RECT 85.660 18.840 85.940 19.120 ;
        RECT 86.180 18.840 86.460 19.120 ;
        RECT 81.700 17.960 81.980 18.240 ;
        RECT 82.220 17.960 82.500 18.240 ;
        RECT 85.660 17.960 85.940 18.240 ;
        RECT 86.180 17.960 86.460 18.240 ;
        RECT 87.820 17.520 88.100 17.800 ;
        RECT 88.340 17.520 88.620 17.800 ;
        RECT 81.700 16.390 81.980 16.670 ;
        RECT 82.220 16.390 82.500 16.670 ;
        RECT 85.660 16.200 85.940 16.480 ;
        RECT 86.180 16.200 86.460 16.480 ;
        RECT 79.620 15.760 79.900 16.040 ;
        RECT 80.140 15.760 80.420 16.040 ;
        RECT 81.700 15.320 81.980 15.600 ;
        RECT 82.220 15.320 82.500 15.600 ;
        RECT 85.660 15.320 85.940 15.600 ;
        RECT 86.180 15.320 86.460 15.600 ;
        RECT 81.700 14.440 81.980 14.720 ;
        RECT 82.220 14.440 82.500 14.720 ;
        RECT 85.660 14.440 85.940 14.720 ;
        RECT 86.180 14.440 86.460 14.720 ;
        RECT 93.160 28.020 94.240 28.375 ;
        RECT 125.920 27.140 127.000 27.495 ;
        RECT 93.160 26.260 94.240 26.615 ;
        RECT 125.920 25.380 127.000 25.735 ;
        RECT 93.160 24.500 94.240 24.855 ;
        RECT 125.920 23.625 127.000 23.975 ;
        RECT 93.160 22.740 94.240 23.095 ;
        RECT 125.920 21.860 127.000 22.215 ;
        RECT 93.160 20.980 94.240 21.335 ;
        RECT 125.920 20.100 127.000 20.455 ;
        RECT 93.160 19.220 94.240 19.575 ;
        RECT 125.920 18.345 127.000 18.695 ;
        RECT 81.700 13.560 81.980 13.840 ;
        RECT 82.220 13.560 82.500 13.840 ;
        RECT 85.660 13.560 85.940 13.840 ;
        RECT 86.180 13.560 86.460 13.840 ;
        RECT 93.160 17.460 94.240 17.815 ;
        RECT 125.920 16.580 127.000 16.935 ;
        RECT 93.160 15.700 94.240 16.055 ;
        RECT 125.920 14.820 127.000 15.175 ;
        RECT 93.160 13.940 94.240 14.295 ;
        RECT 125.920 13.065 127.000 13.415 ;
        RECT 58.740 10.220 59.020 10.500 ;
        RECT 59.260 10.220 59.540 10.500 ;
        RECT 81.700 10.220 81.980 10.500 ;
        RECT 82.220 10.220 82.500 10.500 ;
        RECT 58.740 9.700 59.020 9.980 ;
        RECT 59.260 9.700 59.540 9.980 ;
        RECT 81.700 9.700 81.980 9.980 ;
        RECT 82.220 9.700 82.500 9.980 ;
        RECT 54.780 6.620 55.060 6.900 ;
        RECT 55.300 6.620 55.580 6.900 ;
        RECT 85.660 6.620 85.940 6.900 ;
        RECT 86.180 6.620 86.460 6.900 ;
        RECT 54.780 6.100 55.060 6.380 ;
        RECT 55.300 6.100 55.580 6.380 ;
        RECT 85.660 6.100 85.940 6.380 ;
        RECT 86.180 6.100 86.460 6.380 ;
        RECT 60.900 5.050 61.180 5.330 ;
        RECT 61.420 5.050 61.700 5.330 ;
        RECT 79.620 5.050 79.900 5.330 ;
        RECT 80.140 5.050 80.420 5.330 ;
        RECT 143.740 222.100 144.020 222.380 ;
        RECT 144.260 222.100 144.540 222.380 ;
        RECT 147.700 222.100 147.980 222.380 ;
        RECT 148.220 222.100 148.500 222.380 ;
        RECT 61.660 4.030 61.940 4.310 ;
        RECT 62.180 4.030 62.460 4.310 ;
        RECT 78.780 4.030 79.060 4.310 ;
        RECT 79.300 4.030 79.580 4.310 ;
        RECT 143.740 221.220 144.020 221.500 ;
        RECT 144.260 221.220 144.540 221.500 ;
        RECT 147.700 221.220 147.980 221.500 ;
        RECT 148.220 221.220 148.500 221.500 ;
        RECT 147.700 220.340 147.980 220.620 ;
        RECT 148.220 220.340 148.500 220.620 ;
        RECT 143.740 219.460 144.020 219.740 ;
        RECT 144.260 219.460 144.540 219.740 ;
        RECT 147.700 219.460 147.980 219.740 ;
        RECT 148.220 219.460 148.500 219.740 ;
        RECT 143.740 218.580 144.020 218.860 ;
        RECT 144.260 218.580 144.540 218.860 ;
        RECT 141.580 218.140 141.860 218.420 ;
        RECT 142.100 218.140 142.380 218.420 ;
        RECT 141.580 214.620 141.860 214.900 ;
        RECT 142.100 214.620 142.380 214.900 ;
        RECT 143.740 214.180 144.020 214.460 ;
        RECT 144.260 214.180 144.540 214.460 ;
        RECT 147.700 215.940 147.980 216.220 ;
        RECT 148.220 215.940 148.500 216.220 ;
        RECT 147.700 215.060 147.980 215.340 ;
        RECT 148.220 215.060 148.500 215.340 ;
        RECT 143.740 213.300 144.020 213.580 ;
        RECT 144.260 213.300 144.540 213.580 ;
        RECT 141.580 209.340 141.860 209.620 ;
        RECT 142.100 209.340 142.380 209.620 ;
        RECT 143.740 210.660 144.020 210.940 ;
        RECT 144.260 210.660 144.540 210.940 ;
        RECT 147.700 210.660 147.980 210.940 ;
        RECT 148.220 210.660 148.500 210.940 ;
        RECT 147.700 209.780 147.980 210.060 ;
        RECT 148.220 209.780 148.500 210.060 ;
        RECT 143.740 208.900 144.020 209.180 ;
        RECT 144.260 208.900 144.540 209.180 ;
        RECT 147.700 208.900 147.980 209.180 ;
        RECT 148.220 208.900 148.500 209.180 ;
        RECT 143.740 208.020 144.020 208.300 ;
        RECT 144.260 208.020 144.540 208.300 ;
        RECT 141.580 204.060 141.860 204.340 ;
        RECT 142.100 204.060 142.380 204.340 ;
        RECT 143.740 205.380 144.020 205.660 ;
        RECT 144.260 205.380 144.540 205.660 ;
        RECT 147.700 205.380 147.980 205.660 ;
        RECT 148.220 205.380 148.500 205.660 ;
        RECT 149.860 216.380 150.140 216.660 ;
        RECT 150.380 216.380 150.660 216.660 ;
        RECT 149.860 212.860 150.140 213.140 ;
        RECT 150.380 212.860 150.660 213.140 ;
        RECT 149.860 211.100 150.140 211.380 ;
        RECT 150.380 211.100 150.660 211.380 ;
        RECT 149.860 207.580 150.140 207.860 ;
        RECT 150.380 207.580 150.660 207.860 ;
        RECT 149.860 205.820 150.140 206.100 ;
        RECT 150.380 205.820 150.660 206.100 ;
        RECT 143.740 201.860 144.020 202.140 ;
        RECT 144.260 201.860 144.540 202.140 ;
        RECT 147.700 201.860 147.980 202.140 ;
        RECT 148.220 201.860 148.500 202.140 ;
        RECT 143.740 200.100 144.020 200.380 ;
        RECT 144.260 200.100 144.540 200.380 ;
        RECT 147.700 200.100 147.980 200.380 ;
        RECT 148.220 200.100 148.500 200.380 ;
        RECT 143.740 199.220 144.020 199.500 ;
        RECT 144.260 199.220 144.540 199.500 ;
        RECT 147.700 199.220 147.980 199.500 ;
        RECT 148.220 199.220 148.500 199.500 ;
        RECT 141.580 198.780 141.860 199.060 ;
        RECT 142.100 198.780 142.380 199.060 ;
        RECT 147.700 197.460 147.980 197.740 ;
        RECT 148.220 197.460 148.500 197.740 ;
        RECT 143.740 196.580 144.020 196.860 ;
        RECT 144.260 196.580 144.540 196.860 ;
        RECT 147.700 196.580 147.980 196.860 ;
        RECT 148.220 196.580 148.500 196.860 ;
        RECT 147.700 195.700 147.980 195.980 ;
        RECT 148.220 195.700 148.500 195.980 ;
        RECT 143.740 194.820 144.020 195.100 ;
        RECT 144.260 194.820 144.540 195.100 ;
        RECT 147.700 194.820 147.980 195.100 ;
        RECT 148.220 194.820 148.500 195.100 ;
        RECT 143.740 193.940 144.020 194.220 ;
        RECT 144.260 193.940 144.540 194.220 ;
        RECT 141.580 193.500 141.860 193.780 ;
        RECT 142.100 193.500 142.380 193.780 ;
        RECT 141.580 189.980 141.860 190.260 ;
        RECT 142.100 189.980 142.380 190.260 ;
        RECT 143.740 189.540 144.020 189.820 ;
        RECT 144.260 189.540 144.540 189.820 ;
        RECT 147.700 191.300 147.980 191.580 ;
        RECT 148.220 191.300 148.500 191.580 ;
        RECT 147.700 190.420 147.980 190.700 ;
        RECT 148.220 190.420 148.500 190.700 ;
        RECT 143.740 188.660 144.020 188.940 ;
        RECT 144.260 188.660 144.540 188.940 ;
        RECT 141.580 184.700 141.860 184.980 ;
        RECT 142.100 184.700 142.380 184.980 ;
        RECT 143.740 186.020 144.020 186.300 ;
        RECT 144.260 186.020 144.540 186.300 ;
        RECT 147.700 186.020 147.980 186.300 ;
        RECT 148.220 186.020 148.500 186.300 ;
        RECT 147.700 185.140 147.980 185.420 ;
        RECT 148.220 185.140 148.500 185.420 ;
        RECT 143.740 184.260 144.020 184.540 ;
        RECT 144.260 184.260 144.540 184.540 ;
        RECT 147.700 184.260 147.980 184.540 ;
        RECT 148.220 184.260 148.500 184.540 ;
        RECT 143.740 183.380 144.020 183.660 ;
        RECT 144.260 183.380 144.540 183.660 ;
        RECT 141.580 179.420 141.860 179.700 ;
        RECT 142.100 179.420 142.380 179.700 ;
        RECT 143.740 180.740 144.020 181.020 ;
        RECT 144.260 180.740 144.540 181.020 ;
        RECT 147.700 180.740 147.980 181.020 ;
        RECT 148.220 180.740 148.500 181.020 ;
        RECT 149.860 191.740 150.140 192.020 ;
        RECT 150.380 191.740 150.660 192.020 ;
        RECT 149.860 188.220 150.140 188.500 ;
        RECT 150.380 188.220 150.660 188.500 ;
        RECT 149.860 186.460 150.140 186.740 ;
        RECT 150.380 186.460 150.660 186.740 ;
        RECT 149.860 182.940 150.140 183.220 ;
        RECT 150.380 182.940 150.660 183.220 ;
        RECT 149.860 181.180 150.140 181.460 ;
        RECT 150.380 181.180 150.660 181.460 ;
        RECT 143.740 177.220 144.020 177.500 ;
        RECT 144.260 177.220 144.540 177.500 ;
        RECT 147.700 177.220 147.980 177.500 ;
        RECT 148.220 177.220 148.500 177.500 ;
        RECT 143.740 175.460 144.020 175.740 ;
        RECT 144.260 175.460 144.540 175.740 ;
        RECT 147.700 175.460 147.980 175.740 ;
        RECT 148.220 175.460 148.500 175.740 ;
        RECT 143.740 174.580 144.020 174.860 ;
        RECT 144.260 174.580 144.540 174.860 ;
        RECT 147.700 174.580 147.980 174.860 ;
        RECT 148.220 174.580 148.500 174.860 ;
        RECT 141.580 174.140 141.860 174.420 ;
        RECT 142.100 174.140 142.380 174.420 ;
        RECT 147.700 172.820 147.980 173.100 ;
        RECT 148.220 172.820 148.500 173.100 ;
        RECT 143.740 171.940 144.020 172.220 ;
        RECT 144.260 171.940 144.540 172.220 ;
        RECT 147.700 171.940 147.980 172.220 ;
        RECT 148.220 171.940 148.500 172.220 ;
        RECT 147.700 171.060 147.980 171.340 ;
        RECT 148.220 171.060 148.500 171.340 ;
        RECT 143.740 170.180 144.020 170.460 ;
        RECT 144.260 170.180 144.540 170.460 ;
        RECT 147.700 170.180 147.980 170.460 ;
        RECT 148.220 170.180 148.500 170.460 ;
        RECT 143.740 169.300 144.020 169.580 ;
        RECT 144.260 169.300 144.540 169.580 ;
        RECT 141.580 168.860 141.860 169.140 ;
        RECT 142.100 168.860 142.380 169.140 ;
        RECT 141.580 165.340 141.860 165.620 ;
        RECT 142.100 165.340 142.380 165.620 ;
        RECT 143.740 164.900 144.020 165.180 ;
        RECT 144.260 164.900 144.540 165.180 ;
        RECT 147.700 166.660 147.980 166.940 ;
        RECT 148.220 166.660 148.500 166.940 ;
        RECT 147.700 165.780 147.980 166.060 ;
        RECT 148.220 165.780 148.500 166.060 ;
        RECT 143.740 164.020 144.020 164.300 ;
        RECT 144.260 164.020 144.540 164.300 ;
        RECT 141.580 160.060 141.860 160.340 ;
        RECT 142.100 160.060 142.380 160.340 ;
        RECT 143.740 161.380 144.020 161.660 ;
        RECT 144.260 161.380 144.540 161.660 ;
        RECT 147.700 161.380 147.980 161.660 ;
        RECT 148.220 161.380 148.500 161.660 ;
        RECT 147.700 160.500 147.980 160.780 ;
        RECT 148.220 160.500 148.500 160.780 ;
        RECT 143.740 159.620 144.020 159.900 ;
        RECT 144.260 159.620 144.540 159.900 ;
        RECT 147.700 159.620 147.980 159.900 ;
        RECT 148.220 159.620 148.500 159.900 ;
        RECT 143.740 158.740 144.020 159.020 ;
        RECT 144.260 158.740 144.540 159.020 ;
        RECT 141.580 154.780 141.860 155.060 ;
        RECT 142.100 154.780 142.380 155.060 ;
        RECT 143.740 156.100 144.020 156.380 ;
        RECT 144.260 156.100 144.540 156.380 ;
        RECT 147.700 156.100 147.980 156.380 ;
        RECT 148.220 156.100 148.500 156.380 ;
        RECT 149.860 167.100 150.140 167.380 ;
        RECT 150.380 167.100 150.660 167.380 ;
        RECT 149.860 163.580 150.140 163.860 ;
        RECT 150.380 163.580 150.660 163.860 ;
        RECT 149.860 161.820 150.140 162.100 ;
        RECT 150.380 161.820 150.660 162.100 ;
        RECT 149.860 158.300 150.140 158.580 ;
        RECT 150.380 158.300 150.660 158.580 ;
        RECT 149.860 156.540 150.140 156.820 ;
        RECT 150.380 156.540 150.660 156.820 ;
        RECT 143.740 152.580 144.020 152.860 ;
        RECT 144.260 152.580 144.540 152.860 ;
        RECT 147.700 152.580 147.980 152.860 ;
        RECT 148.220 152.580 148.500 152.860 ;
        RECT 143.740 150.820 144.020 151.100 ;
        RECT 144.260 150.820 144.540 151.100 ;
        RECT 147.700 150.820 147.980 151.100 ;
        RECT 148.220 150.820 148.500 151.100 ;
        RECT 143.740 149.940 144.020 150.220 ;
        RECT 144.260 149.940 144.540 150.220 ;
        RECT 147.700 149.940 147.980 150.220 ;
        RECT 148.220 149.940 148.500 150.220 ;
        RECT 141.580 149.500 141.860 149.780 ;
        RECT 142.100 149.500 142.380 149.780 ;
        RECT 147.700 148.180 147.980 148.460 ;
        RECT 148.220 148.180 148.500 148.460 ;
        RECT 143.740 147.300 144.020 147.580 ;
        RECT 144.260 147.300 144.540 147.580 ;
        RECT 147.700 147.300 147.980 147.580 ;
        RECT 148.220 147.300 148.500 147.580 ;
        RECT 147.700 146.420 147.980 146.700 ;
        RECT 148.220 146.420 148.500 146.700 ;
        RECT 143.740 145.540 144.020 145.820 ;
        RECT 144.260 145.540 144.540 145.820 ;
        RECT 147.700 145.540 147.980 145.820 ;
        RECT 148.220 145.540 148.500 145.820 ;
        RECT 143.740 144.660 144.020 144.940 ;
        RECT 144.260 144.660 144.540 144.940 ;
        RECT 141.580 144.220 141.860 144.500 ;
        RECT 142.100 144.220 142.380 144.500 ;
        RECT 141.580 140.700 141.860 140.980 ;
        RECT 142.100 140.700 142.380 140.980 ;
        RECT 143.740 140.260 144.020 140.540 ;
        RECT 144.260 140.260 144.540 140.540 ;
        RECT 147.700 142.020 147.980 142.300 ;
        RECT 148.220 142.020 148.500 142.300 ;
        RECT 147.700 141.140 147.980 141.420 ;
        RECT 148.220 141.140 148.500 141.420 ;
        RECT 143.740 139.380 144.020 139.660 ;
        RECT 144.260 139.380 144.540 139.660 ;
        RECT 141.580 135.420 141.860 135.700 ;
        RECT 142.100 135.420 142.380 135.700 ;
        RECT 143.740 136.740 144.020 137.020 ;
        RECT 144.260 136.740 144.540 137.020 ;
        RECT 147.700 136.740 147.980 137.020 ;
        RECT 148.220 136.740 148.500 137.020 ;
        RECT 147.700 135.860 147.980 136.140 ;
        RECT 148.220 135.860 148.500 136.140 ;
        RECT 143.740 134.980 144.020 135.260 ;
        RECT 144.260 134.980 144.540 135.260 ;
        RECT 147.700 134.980 147.980 135.260 ;
        RECT 148.220 134.980 148.500 135.260 ;
        RECT 143.740 134.100 144.020 134.380 ;
        RECT 144.260 134.100 144.540 134.380 ;
        RECT 141.580 130.140 141.860 130.420 ;
        RECT 142.100 130.140 142.380 130.420 ;
        RECT 143.740 131.460 144.020 131.740 ;
        RECT 144.260 131.460 144.540 131.740 ;
        RECT 147.700 131.460 147.980 131.740 ;
        RECT 148.220 131.460 148.500 131.740 ;
        RECT 149.860 142.460 150.140 142.740 ;
        RECT 150.380 142.460 150.660 142.740 ;
        RECT 149.860 138.940 150.140 139.220 ;
        RECT 150.380 138.940 150.660 139.220 ;
        RECT 149.860 137.180 150.140 137.460 ;
        RECT 150.380 137.180 150.660 137.460 ;
        RECT 149.860 133.660 150.140 133.940 ;
        RECT 150.380 133.660 150.660 133.940 ;
        RECT 149.860 131.900 150.140 132.180 ;
        RECT 150.380 131.900 150.660 132.180 ;
        RECT 143.740 127.940 144.020 128.220 ;
        RECT 144.260 127.940 144.540 128.220 ;
        RECT 147.700 127.940 147.980 128.220 ;
        RECT 148.220 127.940 148.500 128.220 ;
        RECT 143.740 126.180 144.020 126.460 ;
        RECT 144.260 126.180 144.540 126.460 ;
        RECT 147.700 126.180 147.980 126.460 ;
        RECT 148.220 126.180 148.500 126.460 ;
        RECT 143.740 125.300 144.020 125.580 ;
        RECT 144.260 125.300 144.540 125.580 ;
        RECT 147.700 125.300 147.980 125.580 ;
        RECT 148.220 125.300 148.500 125.580 ;
        RECT 141.580 124.860 141.860 125.140 ;
        RECT 142.100 124.860 142.380 125.140 ;
        RECT 147.700 123.540 147.980 123.820 ;
        RECT 148.220 123.540 148.500 123.820 ;
        RECT 143.740 122.660 144.020 122.940 ;
        RECT 144.260 122.660 144.540 122.940 ;
        RECT 147.700 122.660 147.980 122.940 ;
        RECT 148.220 122.660 148.500 122.940 ;
        RECT 147.700 121.780 147.980 122.060 ;
        RECT 148.220 121.780 148.500 122.060 ;
        RECT 143.740 120.900 144.020 121.180 ;
        RECT 144.260 120.900 144.540 121.180 ;
        RECT 147.700 120.900 147.980 121.180 ;
        RECT 148.220 120.900 148.500 121.180 ;
        RECT 143.740 120.020 144.020 120.300 ;
        RECT 144.260 120.020 144.540 120.300 ;
        RECT 141.580 119.580 141.860 119.860 ;
        RECT 142.100 119.580 142.380 119.860 ;
        RECT 141.580 116.060 141.860 116.340 ;
        RECT 142.100 116.060 142.380 116.340 ;
        RECT 143.740 115.620 144.020 115.900 ;
        RECT 144.260 115.620 144.540 115.900 ;
        RECT 147.700 117.380 147.980 117.660 ;
        RECT 148.220 117.380 148.500 117.660 ;
        RECT 147.700 116.500 147.980 116.780 ;
        RECT 148.220 116.500 148.500 116.780 ;
        RECT 143.740 114.740 144.020 115.020 ;
        RECT 144.260 114.740 144.540 115.020 ;
        RECT 141.580 110.780 141.860 111.060 ;
        RECT 142.100 110.780 142.380 111.060 ;
        RECT 143.740 112.100 144.020 112.380 ;
        RECT 144.260 112.100 144.540 112.380 ;
        RECT 147.700 112.100 147.980 112.380 ;
        RECT 148.220 112.100 148.500 112.380 ;
        RECT 147.700 111.220 147.980 111.500 ;
        RECT 148.220 111.220 148.500 111.500 ;
        RECT 143.740 110.340 144.020 110.620 ;
        RECT 144.260 110.340 144.540 110.620 ;
        RECT 147.700 110.340 147.980 110.620 ;
        RECT 148.220 110.340 148.500 110.620 ;
        RECT 143.740 109.460 144.020 109.740 ;
        RECT 144.260 109.460 144.540 109.740 ;
        RECT 141.580 105.500 141.860 105.780 ;
        RECT 142.100 105.500 142.380 105.780 ;
        RECT 143.740 106.820 144.020 107.100 ;
        RECT 144.260 106.820 144.540 107.100 ;
        RECT 147.700 106.820 147.980 107.100 ;
        RECT 148.220 106.820 148.500 107.100 ;
        RECT 149.860 117.820 150.140 118.100 ;
        RECT 150.380 117.820 150.660 118.100 ;
        RECT 149.860 114.300 150.140 114.580 ;
        RECT 150.380 114.300 150.660 114.580 ;
        RECT 149.860 112.540 150.140 112.820 ;
        RECT 150.380 112.540 150.660 112.820 ;
        RECT 149.860 109.020 150.140 109.300 ;
        RECT 150.380 109.020 150.660 109.300 ;
        RECT 149.860 107.260 150.140 107.540 ;
        RECT 150.380 107.260 150.660 107.540 ;
        RECT 143.740 103.300 144.020 103.580 ;
        RECT 144.260 103.300 144.540 103.580 ;
        RECT 147.700 103.300 147.980 103.580 ;
        RECT 148.220 103.300 148.500 103.580 ;
        RECT 143.740 101.540 144.020 101.820 ;
        RECT 144.260 101.540 144.540 101.820 ;
        RECT 147.700 101.540 147.980 101.820 ;
        RECT 148.220 101.540 148.500 101.820 ;
        RECT 143.740 100.660 144.020 100.940 ;
        RECT 144.260 100.660 144.540 100.940 ;
        RECT 147.700 100.660 147.980 100.940 ;
        RECT 148.220 100.660 148.500 100.940 ;
        RECT 141.580 100.220 141.860 100.500 ;
        RECT 142.100 100.220 142.380 100.500 ;
        RECT 147.700 98.900 147.980 99.180 ;
        RECT 148.220 98.900 148.500 99.180 ;
        RECT 143.740 98.020 144.020 98.300 ;
        RECT 144.260 98.020 144.540 98.300 ;
        RECT 147.700 98.020 147.980 98.300 ;
        RECT 148.220 98.020 148.500 98.300 ;
        RECT 147.700 97.140 147.980 97.420 ;
        RECT 148.220 97.140 148.500 97.420 ;
        RECT 143.740 96.260 144.020 96.540 ;
        RECT 144.260 96.260 144.540 96.540 ;
        RECT 147.700 96.260 147.980 96.540 ;
        RECT 148.220 96.260 148.500 96.540 ;
        RECT 143.740 95.380 144.020 95.660 ;
        RECT 144.260 95.380 144.540 95.660 ;
        RECT 141.580 94.940 141.860 95.220 ;
        RECT 142.100 94.940 142.380 95.220 ;
        RECT 141.580 91.420 141.860 91.700 ;
        RECT 142.100 91.420 142.380 91.700 ;
        RECT 143.740 90.980 144.020 91.260 ;
        RECT 144.260 90.980 144.540 91.260 ;
        RECT 147.700 92.740 147.980 93.020 ;
        RECT 148.220 92.740 148.500 93.020 ;
        RECT 147.700 91.860 147.980 92.140 ;
        RECT 148.220 91.860 148.500 92.140 ;
        RECT 143.740 90.100 144.020 90.380 ;
        RECT 144.260 90.100 144.540 90.380 ;
        RECT 141.580 86.140 141.860 86.420 ;
        RECT 142.100 86.140 142.380 86.420 ;
        RECT 143.740 87.460 144.020 87.740 ;
        RECT 144.260 87.460 144.540 87.740 ;
        RECT 147.700 87.460 147.980 87.740 ;
        RECT 148.220 87.460 148.500 87.740 ;
        RECT 147.700 86.580 147.980 86.860 ;
        RECT 148.220 86.580 148.500 86.860 ;
        RECT 143.740 85.700 144.020 85.980 ;
        RECT 144.260 85.700 144.540 85.980 ;
        RECT 147.700 85.700 147.980 85.980 ;
        RECT 148.220 85.700 148.500 85.980 ;
        RECT 143.740 84.820 144.020 85.100 ;
        RECT 144.260 84.820 144.540 85.100 ;
        RECT 141.580 80.860 141.860 81.140 ;
        RECT 142.100 80.860 142.380 81.140 ;
        RECT 143.740 82.180 144.020 82.460 ;
        RECT 144.260 82.180 144.540 82.460 ;
        RECT 147.700 82.180 147.980 82.460 ;
        RECT 148.220 82.180 148.500 82.460 ;
        RECT 149.860 93.180 150.140 93.460 ;
        RECT 150.380 93.180 150.660 93.460 ;
        RECT 149.860 89.660 150.140 89.940 ;
        RECT 150.380 89.660 150.660 89.940 ;
        RECT 149.860 87.900 150.140 88.180 ;
        RECT 150.380 87.900 150.660 88.180 ;
        RECT 149.860 84.380 150.140 84.660 ;
        RECT 150.380 84.380 150.660 84.660 ;
        RECT 149.860 82.620 150.140 82.900 ;
        RECT 150.380 82.620 150.660 82.900 ;
        RECT 143.740 78.660 144.020 78.940 ;
        RECT 144.260 78.660 144.540 78.940 ;
        RECT 147.700 78.660 147.980 78.940 ;
        RECT 148.220 78.660 148.500 78.940 ;
        RECT 143.740 76.900 144.020 77.180 ;
        RECT 144.260 76.900 144.540 77.180 ;
        RECT 147.700 76.900 147.980 77.180 ;
        RECT 148.220 76.900 148.500 77.180 ;
        RECT 143.740 76.020 144.020 76.300 ;
        RECT 144.260 76.020 144.540 76.300 ;
        RECT 147.700 76.020 147.980 76.300 ;
        RECT 148.220 76.020 148.500 76.300 ;
        RECT 141.580 75.580 141.860 75.860 ;
        RECT 142.100 75.580 142.380 75.860 ;
        RECT 147.700 74.260 147.980 74.540 ;
        RECT 148.220 74.260 148.500 74.540 ;
        RECT 143.740 73.380 144.020 73.660 ;
        RECT 144.260 73.380 144.540 73.660 ;
        RECT 147.700 73.380 147.980 73.660 ;
        RECT 148.220 73.380 148.500 73.660 ;
        RECT 147.700 72.500 147.980 72.780 ;
        RECT 148.220 72.500 148.500 72.780 ;
        RECT 143.740 71.620 144.020 71.900 ;
        RECT 144.260 71.620 144.540 71.900 ;
        RECT 147.700 71.620 147.980 71.900 ;
        RECT 148.220 71.620 148.500 71.900 ;
        RECT 143.740 70.740 144.020 71.020 ;
        RECT 144.260 70.740 144.540 71.020 ;
        RECT 141.580 70.300 141.860 70.580 ;
        RECT 142.100 70.300 142.380 70.580 ;
        RECT 141.580 66.780 141.860 67.060 ;
        RECT 142.100 66.780 142.380 67.060 ;
        RECT 143.740 66.340 144.020 66.620 ;
        RECT 144.260 66.340 144.540 66.620 ;
        RECT 147.700 68.100 147.980 68.380 ;
        RECT 148.220 68.100 148.500 68.380 ;
        RECT 147.700 67.220 147.980 67.500 ;
        RECT 148.220 67.220 148.500 67.500 ;
        RECT 143.740 65.460 144.020 65.740 ;
        RECT 144.260 65.460 144.540 65.740 ;
        RECT 141.580 61.500 141.860 61.780 ;
        RECT 142.100 61.500 142.380 61.780 ;
        RECT 143.740 62.820 144.020 63.100 ;
        RECT 144.260 62.820 144.540 63.100 ;
        RECT 147.700 62.820 147.980 63.100 ;
        RECT 148.220 62.820 148.500 63.100 ;
        RECT 147.700 61.940 147.980 62.220 ;
        RECT 148.220 61.940 148.500 62.220 ;
        RECT 143.740 61.060 144.020 61.340 ;
        RECT 144.260 61.060 144.540 61.340 ;
        RECT 147.700 61.060 147.980 61.340 ;
        RECT 148.220 61.060 148.500 61.340 ;
        RECT 143.740 60.180 144.020 60.460 ;
        RECT 144.260 60.180 144.540 60.460 ;
        RECT 141.580 56.220 141.860 56.500 ;
        RECT 142.100 56.220 142.380 56.500 ;
        RECT 143.740 57.540 144.020 57.820 ;
        RECT 144.260 57.540 144.540 57.820 ;
        RECT 147.700 57.540 147.980 57.820 ;
        RECT 148.220 57.540 148.500 57.820 ;
        RECT 149.860 68.540 150.140 68.820 ;
        RECT 150.380 68.540 150.660 68.820 ;
        RECT 149.860 65.020 150.140 65.300 ;
        RECT 150.380 65.020 150.660 65.300 ;
        RECT 149.860 63.260 150.140 63.540 ;
        RECT 150.380 63.260 150.660 63.540 ;
        RECT 149.860 59.740 150.140 60.020 ;
        RECT 150.380 59.740 150.660 60.020 ;
        RECT 149.860 57.980 150.140 58.260 ;
        RECT 150.380 57.980 150.660 58.260 ;
        RECT 143.740 54.020 144.020 54.300 ;
        RECT 144.260 54.020 144.540 54.300 ;
        RECT 147.700 54.020 147.980 54.300 ;
        RECT 148.220 54.020 148.500 54.300 ;
        RECT 143.740 52.260 144.020 52.540 ;
        RECT 144.260 52.260 144.540 52.540 ;
        RECT 147.700 52.260 147.980 52.540 ;
        RECT 148.220 52.260 148.500 52.540 ;
        RECT 143.740 51.380 144.020 51.660 ;
        RECT 144.260 51.380 144.540 51.660 ;
        RECT 147.700 51.380 147.980 51.660 ;
        RECT 148.220 51.380 148.500 51.660 ;
        RECT 141.580 50.940 141.860 51.220 ;
        RECT 142.100 50.940 142.380 51.220 ;
        RECT 147.700 49.620 147.980 49.900 ;
        RECT 148.220 49.620 148.500 49.900 ;
        RECT 143.740 48.740 144.020 49.020 ;
        RECT 144.260 48.740 144.540 49.020 ;
        RECT 147.700 48.740 147.980 49.020 ;
        RECT 148.220 48.740 148.500 49.020 ;
        RECT 147.700 47.860 147.980 48.140 ;
        RECT 148.220 47.860 148.500 48.140 ;
        RECT 143.740 46.980 144.020 47.260 ;
        RECT 144.260 46.980 144.540 47.260 ;
        RECT 147.700 46.980 147.980 47.260 ;
        RECT 148.220 46.980 148.500 47.260 ;
        RECT 143.740 46.100 144.020 46.380 ;
        RECT 144.260 46.100 144.540 46.380 ;
        RECT 141.580 45.660 141.860 45.940 ;
        RECT 142.100 45.660 142.380 45.940 ;
        RECT 141.580 42.140 141.860 42.420 ;
        RECT 142.100 42.140 142.380 42.420 ;
        RECT 143.740 41.700 144.020 41.980 ;
        RECT 144.260 41.700 144.540 41.980 ;
        RECT 147.700 43.460 147.980 43.740 ;
        RECT 148.220 43.460 148.500 43.740 ;
        RECT 147.700 42.580 147.980 42.860 ;
        RECT 148.220 42.580 148.500 42.860 ;
        RECT 143.740 40.820 144.020 41.100 ;
        RECT 144.260 40.820 144.540 41.100 ;
        RECT 141.580 36.860 141.860 37.140 ;
        RECT 142.100 36.860 142.380 37.140 ;
        RECT 143.740 38.180 144.020 38.460 ;
        RECT 144.260 38.180 144.540 38.460 ;
        RECT 147.700 38.180 147.980 38.460 ;
        RECT 148.220 38.180 148.500 38.460 ;
        RECT 147.700 37.300 147.980 37.580 ;
        RECT 148.220 37.300 148.500 37.580 ;
        RECT 143.740 36.420 144.020 36.700 ;
        RECT 144.260 36.420 144.540 36.700 ;
        RECT 147.700 36.420 147.980 36.700 ;
        RECT 148.220 36.420 148.500 36.700 ;
        RECT 143.740 35.540 144.020 35.820 ;
        RECT 144.260 35.540 144.540 35.820 ;
        RECT 141.580 31.580 141.860 31.860 ;
        RECT 142.100 31.580 142.380 31.860 ;
        RECT 143.740 32.900 144.020 33.180 ;
        RECT 144.260 32.900 144.540 33.180 ;
        RECT 147.700 32.900 147.980 33.180 ;
        RECT 148.220 32.900 148.500 33.180 ;
        RECT 149.860 43.900 150.140 44.180 ;
        RECT 150.380 43.900 150.660 44.180 ;
        RECT 149.860 40.380 150.140 40.660 ;
        RECT 150.380 40.380 150.660 40.660 ;
        RECT 149.860 38.620 150.140 38.900 ;
        RECT 150.380 38.620 150.660 38.900 ;
        RECT 149.860 35.100 150.140 35.380 ;
        RECT 150.380 35.100 150.660 35.380 ;
        RECT 149.860 33.340 150.140 33.620 ;
        RECT 150.380 33.340 150.660 33.620 ;
        RECT 143.740 29.380 144.020 29.660 ;
        RECT 144.260 29.380 144.540 29.660 ;
        RECT 147.700 29.380 147.980 29.660 ;
        RECT 148.220 29.380 148.500 29.660 ;
        RECT 143.740 27.620 144.020 27.900 ;
        RECT 144.260 27.620 144.540 27.900 ;
        RECT 147.700 27.620 147.980 27.900 ;
        RECT 148.220 27.620 148.500 27.900 ;
        RECT 143.740 26.740 144.020 27.020 ;
        RECT 144.260 26.740 144.540 27.020 ;
        RECT 147.700 26.740 147.980 27.020 ;
        RECT 148.220 26.740 148.500 27.020 ;
        RECT 141.580 26.300 141.860 26.580 ;
        RECT 142.100 26.300 142.380 26.580 ;
        RECT 147.700 24.980 147.980 25.260 ;
        RECT 148.220 24.980 148.500 25.260 ;
        RECT 143.740 24.100 144.020 24.380 ;
        RECT 144.260 24.100 144.540 24.380 ;
        RECT 147.700 24.100 147.980 24.380 ;
        RECT 148.220 24.100 148.500 24.380 ;
        RECT 143.740 22.340 144.020 22.620 ;
        RECT 144.260 22.340 144.540 22.620 ;
        RECT 147.700 22.340 147.980 22.620 ;
        RECT 148.220 22.340 148.500 22.620 ;
        RECT 147.700 21.460 147.980 21.740 ;
        RECT 148.220 21.460 148.500 21.740 ;
        RECT 143.740 18.820 144.020 19.100 ;
        RECT 144.260 18.820 144.540 19.100 ;
        RECT 147.700 18.820 147.980 19.100 ;
        RECT 148.220 18.820 148.500 19.100 ;
        RECT 143.740 17.060 144.020 17.340 ;
        RECT 144.260 17.060 144.540 17.340 ;
        RECT 147.700 17.060 147.980 17.340 ;
        RECT 148.220 17.060 148.500 17.340 ;
        RECT 143.740 15.300 144.020 15.580 ;
        RECT 144.260 15.300 144.540 15.580 ;
        RECT 147.700 15.300 147.980 15.580 ;
        RECT 148.220 15.300 148.500 15.580 ;
        RECT 143.740 14.420 144.020 14.700 ;
        RECT 144.260 14.420 144.540 14.700 ;
        RECT 143.740 11.780 144.020 12.060 ;
        RECT 144.260 11.780 144.540 12.060 ;
        RECT 147.700 11.780 147.980 12.060 ;
        RECT 148.220 11.780 148.500 12.060 ;
        RECT 143.740 10.020 144.020 10.300 ;
        RECT 144.260 10.020 144.540 10.300 ;
        RECT 147.700 10.020 147.980 10.300 ;
        RECT 148.220 10.020 148.500 10.300 ;
        RECT 143.740 9.140 144.020 9.420 ;
        RECT 144.260 9.140 144.540 9.420 ;
        RECT 147.700 9.140 147.980 9.420 ;
        RECT 148.220 9.140 148.500 9.420 ;
        RECT 143.740 6.500 144.020 6.780 ;
        RECT 144.260 6.500 144.540 6.780 ;
        RECT 147.700 6.500 147.980 6.780 ;
        RECT 148.220 6.500 148.500 6.780 ;
        RECT 143.740 4.740 144.020 5.020 ;
        RECT 144.260 4.740 144.540 5.020 ;
        RECT 147.700 4.740 147.980 5.020 ;
        RECT 148.220 4.740 148.500 5.020 ;
        RECT 143.740 3.860 144.020 4.140 ;
        RECT 144.260 3.860 144.540 4.140 ;
        RECT 147.700 3.860 147.980 4.140 ;
        RECT 148.220 3.860 148.500 4.140 ;
        RECT 143.740 2.980 144.020 3.260 ;
        RECT 144.260 2.980 144.540 3.260 ;
        RECT 147.700 2.980 147.980 3.260 ;
        RECT 148.220 2.980 148.500 3.260 ;
      LAYER met1 ;
        RECT 24.580 221.190 25.500 222.110 ;
        RECT 27.540 221.190 28.460 222.110 ;
        RECT 49.780 221.190 50.700 222.110 ;
        RECT 52.740 221.190 53.660 222.110 ;
        RECT 74.980 221.190 75.900 222.110 ;
        RECT 77.940 221.190 78.860 222.110 ;
        RECT 100.180 221.190 101.100 222.110 ;
        RECT 103.140 221.190 104.060 222.110 ;
        RECT 143.680 222.070 144.600 222.410 ;
        RECT 147.640 222.070 148.560 222.410 ;
        RECT 143.680 221.190 144.600 221.530 ;
        RECT 147.640 221.190 148.560 221.530 ;
        RECT 147.640 220.610 148.560 220.650 ;
        RECT 147.640 220.310 149.320 220.610 ;
        RECT 143.680 219.430 144.600 219.770 ;
        RECT 147.640 219.430 148.560 219.770 ;
        RECT 143.680 218.850 144.600 218.890 ;
        RECT 143.680 218.550 145.360 218.850 ;
        RECT 21.700 217.590 22.620 218.510 ;
        RECT 30.420 217.590 31.340 218.510 ;
        RECT 46.900 217.590 47.820 218.510 ;
        RECT 55.620 217.590 56.540 218.510 ;
        RECT 72.100 217.590 73.020 218.510 ;
        RECT 80.820 217.590 81.740 218.510 ;
        RECT 97.300 217.590 98.220 218.510 ;
        RECT 106.020 217.590 106.940 218.510 ;
        RECT 122.500 217.590 123.420 218.510 ;
        RECT 141.520 218.110 142.440 218.450 ;
        RECT 17.740 213.990 18.660 214.910 ;
        RECT 34.380 213.990 35.300 214.910 ;
        RECT 42.940 213.990 43.860 214.910 ;
        RECT 59.580 213.990 60.500 214.910 ;
        RECT 68.140 213.990 69.060 214.910 ;
        RECT 84.780 213.990 85.700 214.910 ;
        RECT 93.340 213.990 94.260 214.910 ;
        RECT 109.980 213.990 110.900 214.910 ;
        RECT 118.540 213.990 119.460 214.910 ;
        RECT 141.520 214.890 142.440 214.930 ;
        RECT 140.920 214.590 142.440 214.890 ;
        RECT 17.740 210.800 18.660 211.140 ;
        RECT 21.700 210.800 22.620 211.140 ;
        RECT 30.500 210.800 31.420 211.140 ;
        RECT 34.460 210.800 35.380 211.140 ;
        RECT 42.940 210.800 43.860 211.140 ;
        RECT 46.900 210.800 47.820 211.140 ;
        RECT 55.700 210.800 56.620 211.140 ;
        RECT 59.660 210.800 60.580 211.140 ;
        RECT 68.140 210.800 69.060 211.140 ;
        RECT 72.100 210.800 73.020 211.140 ;
        RECT 80.900 210.800 81.820 211.140 ;
        RECT 84.860 210.800 85.780 211.140 ;
        RECT 93.340 210.800 94.260 211.140 ;
        RECT 97.300 210.800 98.220 211.140 ;
        RECT 106.100 210.800 107.020 211.140 ;
        RECT 110.060 210.800 110.980 211.140 ;
        RECT 17.740 209.920 18.660 210.260 ;
        RECT 21.700 209.920 22.620 210.260 ;
        RECT 30.500 209.920 31.420 210.260 ;
        RECT 34.460 209.920 35.380 210.260 ;
        RECT 42.940 209.920 43.860 210.260 ;
        RECT 46.900 209.920 47.820 210.260 ;
        RECT 55.700 209.920 56.620 210.260 ;
        RECT 59.660 209.920 60.580 210.260 ;
        RECT 68.140 209.920 69.060 210.260 ;
        RECT 72.100 209.920 73.020 210.260 ;
        RECT 80.900 209.920 81.820 210.260 ;
        RECT 84.860 209.920 85.780 210.260 ;
        RECT 93.340 209.920 94.260 210.260 ;
        RECT 97.300 209.920 98.220 210.260 ;
        RECT 106.100 209.920 107.020 210.260 ;
        RECT 110.060 209.920 110.980 210.260 ;
        RECT 21.700 209.230 22.620 209.570 ;
        RECT 30.340 209.340 31.260 209.380 ;
        RECT 32.020 209.340 32.320 209.380 ;
        RECT 30.340 209.040 32.320 209.340 ;
        RECT 46.900 209.230 47.820 209.570 ;
        RECT 55.540 209.340 56.460 209.380 ;
        RECT 57.220 209.340 57.520 209.380 ;
        RECT 55.540 209.040 57.520 209.340 ;
        RECT 72.100 209.230 73.020 209.570 ;
        RECT 80.740 209.340 81.660 209.380 ;
        RECT 82.420 209.340 82.720 209.380 ;
        RECT 80.740 209.040 82.720 209.340 ;
        RECT 97.300 209.230 98.220 209.570 ;
        RECT 105.940 209.040 106.860 209.380 ;
        RECT 118.540 209.040 119.460 209.380 ;
        RECT 122.500 209.040 123.420 209.380 ;
        RECT 17.740 208.160 18.660 208.500 ;
        RECT 21.700 208.160 22.620 208.500 ;
        RECT 30.500 208.160 31.420 208.500 ;
        RECT 4.000 207.140 4.340 207.450 ;
        RECT 17.740 207.280 18.660 207.620 ;
        RECT 15.580 207.140 16.500 207.180 ;
        RECT 4.000 206.840 16.500 207.140 ;
        RECT 4.000 206.530 4.340 206.840 ;
        RECT 32.020 206.540 32.320 209.040 ;
        RECT 34.460 208.160 35.380 208.500 ;
        RECT 42.940 208.160 43.860 208.500 ;
        RECT 46.900 208.160 47.820 208.500 ;
        RECT 55.700 208.160 56.620 208.500 ;
        RECT 34.460 207.280 35.380 207.620 ;
        RECT 42.940 207.280 43.860 207.620 ;
        RECT 36.460 206.840 37.380 207.180 ;
        RECT 40.780 207.140 41.700 207.180 ;
        RECT 40.480 206.840 41.700 207.140 ;
        RECT 40.480 206.540 40.780 206.840 ;
        RECT 32.020 206.240 40.780 206.540 ;
        RECT 57.220 206.540 57.520 209.040 ;
        RECT 59.660 208.160 60.580 208.500 ;
        RECT 68.140 208.160 69.060 208.500 ;
        RECT 72.100 208.160 73.020 208.500 ;
        RECT 80.900 208.160 81.820 208.500 ;
        RECT 59.660 207.280 60.580 207.620 ;
        RECT 68.140 207.280 69.060 207.620 ;
        RECT 61.660 206.840 62.580 207.180 ;
        RECT 65.980 207.140 66.900 207.180 ;
        RECT 65.680 206.840 66.900 207.140 ;
        RECT 65.680 206.540 65.980 206.840 ;
        RECT 57.220 206.240 65.980 206.540 ;
        RECT 82.420 206.540 82.720 209.040 ;
        RECT 84.860 208.160 85.780 208.500 ;
        RECT 93.340 208.160 94.260 208.500 ;
        RECT 97.300 208.160 98.220 208.500 ;
        RECT 106.100 208.160 107.020 208.500 ;
        RECT 110.060 208.160 110.980 208.500 ;
        RECT 118.540 208.160 119.460 208.500 ;
        RECT 122.500 208.160 123.420 208.500 ;
        RECT 84.860 207.280 85.780 207.620 ;
        RECT 93.340 207.280 94.260 207.620 ;
        RECT 110.060 207.280 110.980 207.620 ;
        RECT 86.860 206.840 87.780 207.180 ;
        RECT 91.180 207.140 92.100 207.180 ;
        RECT 90.880 206.840 92.100 207.140 ;
        RECT 112.060 206.840 112.980 207.180 ;
        RECT 116.380 207.030 117.300 207.370 ;
        RECT 90.880 206.540 91.180 206.840 ;
        RECT 82.420 206.240 91.180 206.540 ;
        RECT 118.540 206.400 119.460 206.740 ;
        RECT 122.500 206.400 123.420 206.740 ;
        RECT 118.540 205.520 119.460 205.860 ;
        RECT 124.740 205.080 125.660 205.420 ;
        RECT 17.740 204.640 18.660 204.980 ;
        RECT 21.700 204.640 22.620 204.980 ;
        RECT 30.500 204.640 31.420 204.980 ;
        RECT 34.460 204.640 35.380 204.980 ;
        RECT 42.940 204.640 43.860 204.980 ;
        RECT 46.900 204.640 47.820 204.980 ;
        RECT 55.700 204.640 56.620 204.980 ;
        RECT 59.660 204.640 60.580 204.980 ;
        RECT 68.140 204.640 69.060 204.980 ;
        RECT 72.100 204.640 73.020 204.980 ;
        RECT 80.900 204.640 81.820 204.980 ;
        RECT 84.860 204.640 85.780 204.980 ;
        RECT 93.340 204.640 94.260 204.980 ;
        RECT 97.300 204.640 98.220 204.980 ;
        RECT 106.100 204.640 107.020 204.980 ;
        RECT 110.060 204.640 110.980 204.980 ;
        RECT 124.660 203.320 125.580 203.660 ;
        RECT 17.740 202.880 18.660 203.220 ;
        RECT 21.700 202.880 22.620 203.220 ;
        RECT 30.500 202.880 31.420 203.220 ;
        RECT 34.460 202.880 35.380 203.220 ;
        RECT 42.940 202.880 43.860 203.220 ;
        RECT 46.900 202.880 47.820 203.220 ;
        RECT 55.700 202.880 56.620 203.220 ;
        RECT 59.660 202.880 60.580 203.220 ;
        RECT 68.140 202.880 69.060 203.220 ;
        RECT 72.100 202.880 73.020 203.220 ;
        RECT 80.900 202.880 81.820 203.220 ;
        RECT 84.860 202.880 85.780 203.220 ;
        RECT 93.340 202.880 94.260 203.220 ;
        RECT 97.300 202.880 98.220 203.220 ;
        RECT 106.100 202.880 107.020 203.220 ;
        RECT 110.060 202.880 110.980 203.220 ;
        RECT 118.540 202.880 119.460 203.220 ;
        RECT 122.500 202.880 123.420 203.220 ;
        RECT 21.700 202.000 22.620 202.340 ;
        RECT 30.500 202.000 31.420 202.340 ;
        RECT 46.900 202.000 47.820 202.340 ;
        RECT 55.700 202.000 56.620 202.340 ;
        RECT 72.100 202.000 73.020 202.340 ;
        RECT 80.900 202.000 81.820 202.340 ;
        RECT 97.300 202.000 98.220 202.340 ;
        RECT 106.100 202.000 107.020 202.340 ;
        RECT 118.540 202.300 119.460 202.340 ;
        RECT 117.760 202.000 119.460 202.300 ;
        RECT 122.500 202.000 123.420 202.340 ;
        RECT 15.580 201.860 16.500 201.900 ;
        RECT 36.620 201.860 37.540 201.900 ;
        RECT 15.580 201.560 17.260 201.860 ;
        RECT 16.960 195.260 17.260 201.560 ;
        RECT 35.860 201.560 37.540 201.860 ;
        RECT 40.780 201.860 41.700 201.900 ;
        RECT 61.820 201.860 62.740 201.900 ;
        RECT 40.780 201.560 42.460 201.860 ;
        RECT 17.740 199.360 18.660 199.700 ;
        RECT 21.700 199.360 22.620 199.700 ;
        RECT 30.500 199.360 31.420 199.700 ;
        RECT 34.460 199.360 35.380 199.700 ;
        RECT 17.740 197.600 18.660 197.940 ;
        RECT 21.700 197.600 22.620 197.940 ;
        RECT 30.500 197.600 31.420 197.940 ;
        RECT 34.460 197.600 35.380 197.940 ;
        RECT 23.860 196.580 24.780 196.620 ;
        RECT 28.340 196.580 29.260 196.620 ;
        RECT 23.860 196.280 25.540 196.580 ;
        RECT 17.740 195.840 18.660 196.180 ;
        RECT 21.700 195.840 22.620 196.180 ;
        RECT 17.740 195.260 18.660 195.300 ;
        RECT 16.960 194.960 18.660 195.260 ;
        RECT 23.860 193.060 24.780 193.100 ;
        RECT 23.080 192.760 24.780 193.060 ;
        RECT 17.740 192.320 18.660 192.660 ;
        RECT 21.700 192.320 22.620 192.660 ;
        RECT 17.740 191.440 18.660 191.780 ;
        RECT 21.700 191.440 22.620 191.780 ;
        RECT 15.580 191.000 16.500 191.340 ;
        RECT 17.740 188.800 18.660 189.140 ;
        RECT 17.740 187.920 18.660 188.260 ;
        RECT 21.700 187.920 22.620 188.260 ;
        RECT 17.740 185.280 18.660 185.620 ;
        RECT 17.740 184.400 18.660 184.740 ;
        RECT 21.700 184.400 22.620 184.740 ;
        RECT 20.910 182.290 21.250 183.210 ;
        RECT 17.740 181.760 18.660 182.100 ;
        RECT 21.700 181.760 22.620 182.100 ;
        RECT 17.740 180.880 18.660 181.220 ;
        RECT 21.700 180.880 22.620 181.220 ;
        RECT 17.740 178.240 18.660 178.580 ;
        RECT 17.740 177.360 18.660 177.700 ;
        RECT 21.700 177.360 22.620 177.700 ;
        RECT 15.580 175.460 16.500 175.500 ;
        RECT 15.580 175.160 17.260 175.460 ;
        RECT 20.035 175.250 20.375 176.170 ;
        RECT 15.660 168.080 16.580 168.420 ;
        RECT 15.580 159.620 16.500 159.660 ;
        RECT 14.980 159.320 16.500 159.620 ;
        RECT 14.980 154.340 15.280 159.320 ;
        RECT 15.580 155.800 16.500 156.140 ;
        RECT 16.960 154.780 17.260 175.160 ;
        RECT 17.740 174.720 18.660 175.060 ;
        RECT 21.700 174.720 22.620 175.060 ;
        RECT 17.740 173.840 18.660 174.180 ;
        RECT 21.700 173.840 22.620 174.180 ;
        RECT 17.740 171.200 18.660 171.540 ;
        RECT 17.740 170.320 18.660 170.660 ;
        RECT 21.700 170.320 22.620 170.660 ;
        RECT 19.235 168.210 19.575 169.130 ;
        RECT 21.700 168.860 22.620 168.900 ;
        RECT 23.080 168.860 23.380 192.760 ;
        RECT 21.700 168.560 23.380 168.860 ;
        RECT 17.740 167.680 18.660 168.020 ;
        RECT 21.700 167.680 22.620 168.020 ;
        RECT 17.740 166.800 18.660 167.140 ;
        RECT 21.700 166.800 22.620 167.140 ;
        RECT 17.740 164.160 18.660 164.500 ;
        RECT 17.740 163.280 18.660 163.620 ;
        RECT 21.700 163.280 22.620 163.620 ;
        RECT 17.740 160.640 18.660 160.980 ;
        RECT 21.700 160.640 22.620 160.980 ;
        RECT 23.860 159.320 24.780 159.660 ;
        RECT 17.740 155.360 18.660 155.700 ;
        RECT 21.700 155.360 22.620 155.700 ;
        RECT 17.740 154.780 18.660 154.820 ;
        RECT 16.960 154.480 18.660 154.780 ;
        RECT 15.580 154.340 16.500 154.380 ;
        RECT 14.980 154.040 16.500 154.340 ;
        RECT 14.980 142.020 15.280 154.040 ;
        RECT 15.740 150.820 16.660 150.860 ;
        RECT 15.660 150.520 17.260 150.820 ;
        RECT 15.660 150.480 16.580 150.520 ;
        RECT 15.740 145.540 16.660 145.580 ;
        RECT 16.960 145.540 17.260 150.520 ;
        RECT 17.740 150.080 18.660 150.420 ;
        RECT 21.700 150.080 22.620 150.420 ;
        RECT 17.740 148.320 18.660 148.660 ;
        RECT 21.700 148.320 22.620 148.660 ;
        RECT 21.700 147.440 22.620 147.780 ;
        RECT 17.740 146.560 18.660 146.900 ;
        RECT 17.740 145.680 18.660 146.020 ;
        RECT 15.740 145.240 17.260 145.540 ;
        RECT 17.740 143.040 18.660 143.380 ;
        RECT 21.700 143.340 22.620 143.380 ;
        RECT 25.240 143.340 25.540 196.280 ;
        RECT 21.700 143.040 25.540 143.340 ;
        RECT 27.580 196.280 29.260 196.580 ;
        RECT 27.580 143.340 27.880 196.280 ;
        RECT 30.500 195.840 31.420 196.180 ;
        RECT 34.460 195.840 35.380 196.180 ;
        RECT 34.460 195.260 35.380 195.300 ;
        RECT 35.860 195.260 36.160 201.560 ;
        RECT 34.460 194.960 36.160 195.260 ;
        RECT 42.160 195.260 42.460 201.560 ;
        RECT 61.060 201.560 62.740 201.860 ;
        RECT 65.980 201.860 66.900 201.900 ;
        RECT 87.020 201.860 87.940 201.900 ;
        RECT 65.980 201.560 67.660 201.860 ;
        RECT 42.940 199.360 43.860 199.700 ;
        RECT 46.900 199.360 47.820 199.700 ;
        RECT 55.700 199.360 56.620 199.700 ;
        RECT 59.660 199.360 60.580 199.700 ;
        RECT 42.940 197.600 43.860 197.940 ;
        RECT 46.900 197.600 47.820 197.940 ;
        RECT 55.700 197.600 56.620 197.940 ;
        RECT 59.660 197.600 60.580 197.940 ;
        RECT 49.060 196.580 49.980 196.620 ;
        RECT 53.540 196.580 54.460 196.620 ;
        RECT 49.060 196.280 50.740 196.580 ;
        RECT 42.940 195.840 43.860 196.180 ;
        RECT 46.900 195.840 47.820 196.180 ;
        RECT 42.940 195.260 43.860 195.300 ;
        RECT 42.160 194.960 43.860 195.260 ;
        RECT 28.340 193.060 29.260 193.100 ;
        RECT 49.060 193.060 49.980 193.100 ;
        RECT 28.340 192.760 30.040 193.060 ;
        RECT 29.740 168.860 30.040 192.760 ;
        RECT 48.280 192.760 49.980 193.060 ;
        RECT 30.500 192.320 31.420 192.660 ;
        RECT 34.460 192.320 35.380 192.660 ;
        RECT 42.940 192.320 43.860 192.660 ;
        RECT 46.900 192.320 47.820 192.660 ;
        RECT 30.500 191.440 31.420 191.780 ;
        RECT 34.460 191.440 35.380 191.780 ;
        RECT 42.940 191.440 43.860 191.780 ;
        RECT 46.900 191.440 47.820 191.780 ;
        RECT 36.460 191.000 37.380 191.340 ;
        RECT 40.780 191.000 41.700 191.340 ;
        RECT 34.460 188.800 35.380 189.140 ;
        RECT 42.940 188.800 43.860 189.140 ;
        RECT 30.500 187.920 31.420 188.260 ;
        RECT 34.460 187.920 35.380 188.260 ;
        RECT 42.940 187.920 43.860 188.260 ;
        RECT 46.900 187.920 47.820 188.260 ;
        RECT 34.460 185.280 35.380 185.620 ;
        RECT 42.940 185.280 43.860 185.620 ;
        RECT 30.500 184.400 31.420 184.740 ;
        RECT 34.460 184.400 35.380 184.740 ;
        RECT 42.940 184.400 43.860 184.740 ;
        RECT 46.900 184.400 47.820 184.740 ;
        RECT 31.870 182.290 32.210 183.210 ;
        RECT 46.110 182.290 46.450 183.210 ;
        RECT 30.500 181.760 31.420 182.100 ;
        RECT 34.460 181.760 35.380 182.100 ;
        RECT 42.940 181.760 43.860 182.100 ;
        RECT 46.900 181.760 47.820 182.100 ;
        RECT 30.500 180.880 31.420 181.220 ;
        RECT 34.460 180.880 35.380 181.220 ;
        RECT 42.940 180.880 43.860 181.220 ;
        RECT 46.900 180.880 47.820 181.220 ;
        RECT 34.460 178.240 35.380 178.580 ;
        RECT 42.940 178.240 43.860 178.580 ;
        RECT 30.500 177.360 31.420 177.700 ;
        RECT 34.460 177.360 35.380 177.700 ;
        RECT 42.940 177.360 43.860 177.700 ;
        RECT 46.900 177.360 47.820 177.700 ;
        RECT 32.745 175.250 33.085 176.170 ;
        RECT 36.620 175.460 37.540 175.500 ;
        RECT 35.860 175.160 37.540 175.460 ;
        RECT 40.780 175.460 41.700 175.500 ;
        RECT 40.780 175.160 42.460 175.460 ;
        RECT 45.235 175.250 45.575 176.170 ;
        RECT 30.500 174.720 31.420 175.060 ;
        RECT 34.460 174.720 35.380 175.060 ;
        RECT 30.500 173.840 31.420 174.180 ;
        RECT 34.460 173.840 35.380 174.180 ;
        RECT 34.460 171.200 35.380 171.540 ;
        RECT 30.500 170.320 31.420 170.660 ;
        RECT 34.460 170.320 35.380 170.660 ;
        RECT 30.500 168.860 31.420 168.900 ;
        RECT 29.740 168.560 31.420 168.860 ;
        RECT 33.545 168.210 33.885 169.130 ;
        RECT 30.500 167.680 31.420 168.020 ;
        RECT 34.460 167.680 35.380 168.020 ;
        RECT 30.500 166.800 31.420 167.140 ;
        RECT 34.460 166.800 35.380 167.140 ;
        RECT 34.460 164.160 35.380 164.500 ;
        RECT 30.500 163.280 31.420 163.620 ;
        RECT 34.460 163.280 35.380 163.620 ;
        RECT 30.500 160.640 31.420 160.980 ;
        RECT 34.460 160.640 35.380 160.980 ;
        RECT 28.180 159.320 29.100 159.660 ;
        RECT 30.500 155.360 31.420 155.700 ;
        RECT 34.460 155.360 35.380 155.700 ;
        RECT 34.460 154.780 35.380 154.820 ;
        RECT 35.860 154.780 36.160 175.160 ;
        RECT 36.540 168.080 37.460 168.420 ;
        RECT 40.860 168.080 41.780 168.420 ;
        RECT 36.620 159.620 37.540 159.660 ;
        RECT 40.780 159.620 41.700 159.660 ;
        RECT 36.620 159.320 38.140 159.620 ;
        RECT 36.460 155.800 37.380 156.140 ;
        RECT 34.460 154.480 36.160 154.780 ;
        RECT 36.620 154.340 37.540 154.380 ;
        RECT 37.840 154.340 38.140 159.320 ;
        RECT 36.620 154.040 38.140 154.340 ;
        RECT 36.460 150.820 37.380 150.860 ;
        RECT 35.860 150.520 37.460 150.820 ;
        RECT 30.500 150.080 31.420 150.420 ;
        RECT 34.460 150.080 35.380 150.420 ;
        RECT 30.500 148.320 31.420 148.660 ;
        RECT 34.460 148.320 35.380 148.660 ;
        RECT 30.500 147.440 31.420 147.780 ;
        RECT 34.460 146.560 35.380 146.900 ;
        RECT 34.460 145.680 35.380 146.020 ;
        RECT 35.860 145.540 36.160 150.520 ;
        RECT 36.540 150.480 37.460 150.520 ;
        RECT 36.460 145.540 37.380 145.580 ;
        RECT 35.860 145.240 37.380 145.540 ;
        RECT 30.500 143.340 31.420 143.380 ;
        RECT 27.580 143.040 31.420 143.340 ;
        RECT 34.460 143.040 35.380 143.380 ;
        RECT 21.780 143.000 22.700 143.040 ;
        RECT 30.420 143.000 31.340 143.040 ;
        RECT 21.700 142.160 22.620 142.500 ;
        RECT 30.500 142.160 31.420 142.500 ;
        RECT 15.580 142.020 16.500 142.060 ;
        RECT 36.620 142.020 37.540 142.060 ;
        RECT 37.840 142.020 38.140 154.040 ;
        RECT 14.980 141.720 16.580 142.020 ;
        RECT 15.660 141.680 16.580 141.720 ;
        RECT 36.540 141.720 38.140 142.020 ;
        RECT 40.180 159.320 41.700 159.620 ;
        RECT 40.180 154.340 40.480 159.320 ;
        RECT 40.780 155.800 41.700 156.140 ;
        RECT 42.160 154.780 42.460 175.160 ;
        RECT 42.940 174.720 43.860 175.060 ;
        RECT 46.900 174.720 47.820 175.060 ;
        RECT 42.940 173.840 43.860 174.180 ;
        RECT 46.900 173.840 47.820 174.180 ;
        RECT 42.940 171.200 43.860 171.540 ;
        RECT 42.940 170.320 43.860 170.660 ;
        RECT 46.900 170.320 47.820 170.660 ;
        RECT 44.435 168.210 44.775 169.130 ;
        RECT 46.900 168.860 47.820 168.900 ;
        RECT 48.280 168.860 48.580 192.760 ;
        RECT 46.900 168.560 48.580 168.860 ;
        RECT 42.940 167.680 43.860 168.020 ;
        RECT 46.900 167.680 47.820 168.020 ;
        RECT 42.940 166.800 43.860 167.140 ;
        RECT 46.900 166.800 47.820 167.140 ;
        RECT 42.940 164.160 43.860 164.500 ;
        RECT 42.940 163.280 43.860 163.620 ;
        RECT 46.900 163.280 47.820 163.620 ;
        RECT 42.940 160.640 43.860 160.980 ;
        RECT 46.900 160.640 47.820 160.980 ;
        RECT 49.060 159.320 49.980 159.660 ;
        RECT 42.940 155.360 43.860 155.700 ;
        RECT 46.900 155.360 47.820 155.700 ;
        RECT 42.940 154.780 43.860 154.820 ;
        RECT 42.160 154.480 43.860 154.780 ;
        RECT 40.780 154.340 41.700 154.380 ;
        RECT 40.180 154.040 41.700 154.340 ;
        RECT 40.180 142.020 40.480 154.040 ;
        RECT 40.940 150.820 41.860 150.860 ;
        RECT 40.860 150.520 42.460 150.820 ;
        RECT 40.860 150.480 41.780 150.520 ;
        RECT 40.940 145.540 41.860 145.580 ;
        RECT 42.160 145.540 42.460 150.520 ;
        RECT 42.940 150.080 43.860 150.420 ;
        RECT 46.900 150.080 47.820 150.420 ;
        RECT 42.940 148.320 43.860 148.660 ;
        RECT 46.900 148.320 47.820 148.660 ;
        RECT 46.900 147.440 47.820 147.780 ;
        RECT 42.940 146.560 43.860 146.900 ;
        RECT 42.940 145.680 43.860 146.020 ;
        RECT 40.940 145.240 42.460 145.540 ;
        RECT 42.940 143.040 43.860 143.380 ;
        RECT 46.900 143.340 47.820 143.380 ;
        RECT 50.440 143.340 50.740 196.280 ;
        RECT 46.900 143.040 50.740 143.340 ;
        RECT 52.780 196.280 54.460 196.580 ;
        RECT 52.780 143.340 53.080 196.280 ;
        RECT 55.700 195.840 56.620 196.180 ;
        RECT 59.660 195.840 60.580 196.180 ;
        RECT 59.660 195.260 60.580 195.300 ;
        RECT 61.060 195.260 61.360 201.560 ;
        RECT 59.660 194.960 61.360 195.260 ;
        RECT 67.360 195.260 67.660 201.560 ;
        RECT 86.260 201.560 87.940 201.860 ;
        RECT 91.180 201.860 92.100 201.900 ;
        RECT 112.220 201.860 113.140 201.900 ;
        RECT 91.180 201.560 92.860 201.860 ;
        RECT 68.140 199.360 69.060 199.700 ;
        RECT 72.100 199.360 73.020 199.700 ;
        RECT 80.900 199.360 81.820 199.700 ;
        RECT 84.860 199.360 85.780 199.700 ;
        RECT 68.140 197.600 69.060 197.940 ;
        RECT 72.100 197.600 73.020 197.940 ;
        RECT 80.900 197.600 81.820 197.940 ;
        RECT 84.860 197.600 85.780 197.940 ;
        RECT 74.260 196.580 75.180 196.620 ;
        RECT 78.740 196.580 79.660 196.620 ;
        RECT 74.260 196.280 75.940 196.580 ;
        RECT 68.140 195.840 69.060 196.180 ;
        RECT 72.100 195.840 73.020 196.180 ;
        RECT 68.140 195.260 69.060 195.300 ;
        RECT 67.360 194.960 69.060 195.260 ;
        RECT 53.540 193.060 54.460 193.100 ;
        RECT 74.260 193.060 75.180 193.100 ;
        RECT 53.540 192.760 55.240 193.060 ;
        RECT 54.940 168.860 55.240 192.760 ;
        RECT 73.480 192.760 75.180 193.060 ;
        RECT 55.700 192.320 56.620 192.660 ;
        RECT 59.660 192.320 60.580 192.660 ;
        RECT 68.140 192.320 69.060 192.660 ;
        RECT 72.100 192.320 73.020 192.660 ;
        RECT 55.700 191.440 56.620 191.780 ;
        RECT 59.660 191.440 60.580 191.780 ;
        RECT 68.140 191.440 69.060 191.780 ;
        RECT 72.100 191.440 73.020 191.780 ;
        RECT 61.660 191.000 62.580 191.340 ;
        RECT 65.980 191.000 66.900 191.340 ;
        RECT 59.660 188.800 60.580 189.140 ;
        RECT 68.140 188.800 69.060 189.140 ;
        RECT 55.700 187.920 56.620 188.260 ;
        RECT 59.660 187.920 60.580 188.260 ;
        RECT 68.140 187.920 69.060 188.260 ;
        RECT 72.100 187.920 73.020 188.260 ;
        RECT 59.660 185.280 60.580 185.620 ;
        RECT 68.140 185.280 69.060 185.620 ;
        RECT 55.700 184.400 56.620 184.740 ;
        RECT 59.660 184.400 60.580 184.740 ;
        RECT 68.140 184.400 69.060 184.740 ;
        RECT 72.100 184.400 73.020 184.740 ;
        RECT 57.070 182.290 57.410 183.210 ;
        RECT 71.310 182.290 71.650 183.210 ;
        RECT 55.700 181.760 56.620 182.100 ;
        RECT 59.660 181.760 60.580 182.100 ;
        RECT 68.140 181.760 69.060 182.100 ;
        RECT 72.100 181.760 73.020 182.100 ;
        RECT 55.700 180.880 56.620 181.220 ;
        RECT 59.660 180.880 60.580 181.220 ;
        RECT 68.140 180.880 69.060 181.220 ;
        RECT 72.100 180.880 73.020 181.220 ;
        RECT 59.660 178.240 60.580 178.580 ;
        RECT 68.140 178.240 69.060 178.580 ;
        RECT 55.700 177.360 56.620 177.700 ;
        RECT 59.660 177.360 60.580 177.700 ;
        RECT 68.140 177.360 69.060 177.700 ;
        RECT 72.100 177.360 73.020 177.700 ;
        RECT 57.945 175.250 58.285 176.170 ;
        RECT 61.820 175.460 62.740 175.500 ;
        RECT 61.060 175.160 62.740 175.460 ;
        RECT 65.980 175.460 66.900 175.500 ;
        RECT 65.980 175.160 67.660 175.460 ;
        RECT 70.435 175.250 70.775 176.170 ;
        RECT 55.700 174.720 56.620 175.060 ;
        RECT 59.660 174.720 60.580 175.060 ;
        RECT 55.700 173.840 56.620 174.180 ;
        RECT 59.660 173.840 60.580 174.180 ;
        RECT 59.660 171.200 60.580 171.540 ;
        RECT 55.700 170.320 56.620 170.660 ;
        RECT 59.660 170.320 60.580 170.660 ;
        RECT 55.700 168.860 56.620 168.900 ;
        RECT 54.940 168.560 56.620 168.860 ;
        RECT 58.745 168.210 59.085 169.130 ;
        RECT 55.700 167.680 56.620 168.020 ;
        RECT 59.660 167.680 60.580 168.020 ;
        RECT 55.700 166.800 56.620 167.140 ;
        RECT 59.660 166.800 60.580 167.140 ;
        RECT 59.660 164.160 60.580 164.500 ;
        RECT 55.700 163.280 56.620 163.620 ;
        RECT 59.660 163.280 60.580 163.620 ;
        RECT 55.700 160.640 56.620 160.980 ;
        RECT 59.660 160.640 60.580 160.980 ;
        RECT 53.380 159.320 54.300 159.660 ;
        RECT 55.700 155.360 56.620 155.700 ;
        RECT 59.660 155.360 60.580 155.700 ;
        RECT 59.660 154.780 60.580 154.820 ;
        RECT 61.060 154.780 61.360 175.160 ;
        RECT 61.740 168.080 62.660 168.420 ;
        RECT 66.060 168.080 66.980 168.420 ;
        RECT 61.820 159.620 62.740 159.660 ;
        RECT 65.980 159.620 66.900 159.660 ;
        RECT 61.820 159.320 63.340 159.620 ;
        RECT 61.660 155.800 62.580 156.140 ;
        RECT 59.660 154.480 61.360 154.780 ;
        RECT 61.820 154.340 62.740 154.380 ;
        RECT 63.040 154.340 63.340 159.320 ;
        RECT 61.820 154.040 63.340 154.340 ;
        RECT 61.660 150.820 62.580 150.860 ;
        RECT 61.060 150.520 62.660 150.820 ;
        RECT 55.700 150.080 56.620 150.420 ;
        RECT 59.660 150.080 60.580 150.420 ;
        RECT 55.700 148.320 56.620 148.660 ;
        RECT 59.660 148.320 60.580 148.660 ;
        RECT 55.700 147.440 56.620 147.780 ;
        RECT 59.660 146.560 60.580 146.900 ;
        RECT 59.660 145.680 60.580 146.020 ;
        RECT 61.060 145.540 61.360 150.520 ;
        RECT 61.740 150.480 62.660 150.520 ;
        RECT 61.660 145.540 62.580 145.580 ;
        RECT 61.060 145.240 62.580 145.540 ;
        RECT 55.700 143.340 56.620 143.380 ;
        RECT 52.780 143.040 56.620 143.340 ;
        RECT 59.660 143.040 60.580 143.380 ;
        RECT 46.980 143.000 47.900 143.040 ;
        RECT 55.620 143.000 56.540 143.040 ;
        RECT 46.900 142.160 47.820 142.500 ;
        RECT 55.700 142.160 56.620 142.500 ;
        RECT 40.780 142.020 41.700 142.060 ;
        RECT 61.820 142.020 62.740 142.060 ;
        RECT 63.040 142.020 63.340 154.040 ;
        RECT 40.180 141.720 41.780 142.020 ;
        RECT 36.540 141.680 37.460 141.720 ;
        RECT 40.860 141.680 41.780 141.720 ;
        RECT 61.740 141.720 63.340 142.020 ;
        RECT 65.380 159.320 66.900 159.620 ;
        RECT 65.380 154.340 65.680 159.320 ;
        RECT 65.980 155.800 66.900 156.140 ;
        RECT 67.360 154.780 67.660 175.160 ;
        RECT 68.140 174.720 69.060 175.060 ;
        RECT 72.100 174.720 73.020 175.060 ;
        RECT 68.140 173.840 69.060 174.180 ;
        RECT 72.100 173.840 73.020 174.180 ;
        RECT 68.140 171.200 69.060 171.540 ;
        RECT 68.140 170.320 69.060 170.660 ;
        RECT 72.100 170.320 73.020 170.660 ;
        RECT 69.635 168.210 69.975 169.130 ;
        RECT 72.100 168.860 73.020 168.900 ;
        RECT 73.480 168.860 73.780 192.760 ;
        RECT 72.100 168.560 73.780 168.860 ;
        RECT 68.140 167.680 69.060 168.020 ;
        RECT 72.100 167.680 73.020 168.020 ;
        RECT 68.140 166.800 69.060 167.140 ;
        RECT 72.100 166.800 73.020 167.140 ;
        RECT 68.140 164.160 69.060 164.500 ;
        RECT 68.140 163.280 69.060 163.620 ;
        RECT 72.100 163.280 73.020 163.620 ;
        RECT 68.140 160.640 69.060 160.980 ;
        RECT 72.100 160.640 73.020 160.980 ;
        RECT 74.260 159.320 75.180 159.660 ;
        RECT 68.140 155.360 69.060 155.700 ;
        RECT 72.100 155.360 73.020 155.700 ;
        RECT 68.140 154.780 69.060 154.820 ;
        RECT 67.360 154.480 69.060 154.780 ;
        RECT 65.980 154.340 66.900 154.380 ;
        RECT 65.380 154.040 66.900 154.340 ;
        RECT 65.380 142.020 65.680 154.040 ;
        RECT 66.140 150.820 67.060 150.860 ;
        RECT 66.060 150.520 67.660 150.820 ;
        RECT 66.060 150.480 66.980 150.520 ;
        RECT 66.140 145.540 67.060 145.580 ;
        RECT 67.360 145.540 67.660 150.520 ;
        RECT 68.140 150.080 69.060 150.420 ;
        RECT 72.100 150.080 73.020 150.420 ;
        RECT 68.140 148.320 69.060 148.660 ;
        RECT 72.100 148.320 73.020 148.660 ;
        RECT 72.100 147.440 73.020 147.780 ;
        RECT 68.140 146.560 69.060 146.900 ;
        RECT 68.140 145.680 69.060 146.020 ;
        RECT 66.140 145.240 67.660 145.540 ;
        RECT 68.140 143.040 69.060 143.380 ;
        RECT 72.100 143.340 73.020 143.380 ;
        RECT 75.640 143.340 75.940 196.280 ;
        RECT 72.100 143.040 75.940 143.340 ;
        RECT 77.980 196.280 79.660 196.580 ;
        RECT 77.980 143.340 78.280 196.280 ;
        RECT 80.900 195.840 81.820 196.180 ;
        RECT 84.860 195.840 85.780 196.180 ;
        RECT 84.860 195.260 85.780 195.300 ;
        RECT 86.260 195.260 86.560 201.560 ;
        RECT 84.860 194.960 86.560 195.260 ;
        RECT 92.560 195.260 92.860 201.560 ;
        RECT 111.460 201.560 113.140 201.860 ;
        RECT 93.340 199.360 94.260 199.700 ;
        RECT 97.300 199.360 98.220 199.700 ;
        RECT 106.100 199.360 107.020 199.700 ;
        RECT 110.060 199.360 110.980 199.700 ;
        RECT 109.980 198.480 110.900 198.820 ;
        RECT 93.340 197.600 94.260 197.940 ;
        RECT 97.300 197.600 98.220 197.940 ;
        RECT 106.100 197.600 107.020 197.940 ;
        RECT 110.060 197.600 110.980 197.940 ;
        RECT 99.460 196.580 100.380 196.620 ;
        RECT 103.940 196.580 104.860 196.620 ;
        RECT 99.460 196.280 101.140 196.580 ;
        RECT 93.340 195.840 94.260 196.180 ;
        RECT 97.300 195.840 98.220 196.180 ;
        RECT 93.340 195.260 94.260 195.300 ;
        RECT 92.560 194.960 94.260 195.260 ;
        RECT 78.740 193.060 79.660 193.100 ;
        RECT 99.460 193.060 100.380 193.100 ;
        RECT 78.740 192.760 80.440 193.060 ;
        RECT 80.140 168.860 80.440 192.760 ;
        RECT 98.680 192.760 100.380 193.060 ;
        RECT 80.900 192.320 81.820 192.660 ;
        RECT 84.860 192.320 85.780 192.660 ;
        RECT 93.340 192.320 94.260 192.660 ;
        RECT 97.300 192.320 98.220 192.660 ;
        RECT 80.900 191.440 81.820 191.780 ;
        RECT 84.860 191.440 85.780 191.780 ;
        RECT 93.340 191.440 94.260 191.780 ;
        RECT 97.300 191.440 98.220 191.780 ;
        RECT 86.860 191.000 87.780 191.340 ;
        RECT 91.180 191.000 92.100 191.340 ;
        RECT 84.860 188.800 85.780 189.140 ;
        RECT 93.340 188.800 94.260 189.140 ;
        RECT 80.900 187.920 81.820 188.260 ;
        RECT 84.860 187.920 85.780 188.260 ;
        RECT 93.340 187.920 94.260 188.260 ;
        RECT 97.300 187.920 98.220 188.260 ;
        RECT 84.860 185.280 85.780 185.620 ;
        RECT 93.340 185.280 94.260 185.620 ;
        RECT 80.900 184.400 81.820 184.740 ;
        RECT 84.860 184.400 85.780 184.740 ;
        RECT 93.340 184.400 94.260 184.740 ;
        RECT 97.300 184.400 98.220 184.740 ;
        RECT 82.270 182.290 82.610 183.210 ;
        RECT 96.510 182.290 96.850 183.210 ;
        RECT 80.900 181.760 81.820 182.100 ;
        RECT 84.860 181.760 85.780 182.100 ;
        RECT 93.340 181.760 94.260 182.100 ;
        RECT 97.300 181.760 98.220 182.100 ;
        RECT 80.900 180.880 81.820 181.220 ;
        RECT 84.860 180.880 85.780 181.220 ;
        RECT 93.340 180.880 94.260 181.220 ;
        RECT 97.300 180.880 98.220 181.220 ;
        RECT 84.860 178.240 85.780 178.580 ;
        RECT 93.340 178.240 94.260 178.580 ;
        RECT 80.900 177.360 81.820 177.700 ;
        RECT 84.860 177.360 85.780 177.700 ;
        RECT 93.340 177.360 94.260 177.700 ;
        RECT 97.300 177.360 98.220 177.700 ;
        RECT 83.145 175.250 83.485 176.170 ;
        RECT 87.020 175.460 87.940 175.500 ;
        RECT 86.260 175.160 87.940 175.460 ;
        RECT 91.180 175.460 92.100 175.500 ;
        RECT 91.180 175.160 92.860 175.460 ;
        RECT 95.635 175.250 95.975 176.170 ;
        RECT 80.900 174.720 81.820 175.060 ;
        RECT 84.860 174.720 85.780 175.060 ;
        RECT 80.900 173.840 81.820 174.180 ;
        RECT 84.860 173.840 85.780 174.180 ;
        RECT 84.860 171.200 85.780 171.540 ;
        RECT 80.900 170.320 81.820 170.660 ;
        RECT 84.860 170.320 85.780 170.660 ;
        RECT 80.900 168.860 81.820 168.900 ;
        RECT 80.140 168.560 81.820 168.860 ;
        RECT 83.945 168.210 84.285 169.130 ;
        RECT 80.900 167.680 81.820 168.020 ;
        RECT 84.860 167.680 85.780 168.020 ;
        RECT 80.900 166.800 81.820 167.140 ;
        RECT 84.860 166.800 85.780 167.140 ;
        RECT 84.860 164.160 85.780 164.500 ;
        RECT 80.900 163.280 81.820 163.620 ;
        RECT 84.860 163.280 85.780 163.620 ;
        RECT 80.900 160.640 81.820 160.980 ;
        RECT 84.860 160.640 85.780 160.980 ;
        RECT 78.580 159.320 79.500 159.660 ;
        RECT 80.900 155.360 81.820 155.700 ;
        RECT 84.860 155.360 85.780 155.700 ;
        RECT 84.860 154.780 85.780 154.820 ;
        RECT 86.260 154.780 86.560 175.160 ;
        RECT 86.940 168.080 87.860 168.420 ;
        RECT 91.260 168.080 92.180 168.420 ;
        RECT 87.020 159.620 87.940 159.660 ;
        RECT 91.180 159.620 92.100 159.660 ;
        RECT 87.020 159.320 88.540 159.620 ;
        RECT 86.860 155.800 87.780 156.140 ;
        RECT 84.860 154.480 86.560 154.780 ;
        RECT 87.020 154.340 87.940 154.380 ;
        RECT 88.240 154.340 88.540 159.320 ;
        RECT 87.020 154.040 88.540 154.340 ;
        RECT 86.860 150.820 87.780 150.860 ;
        RECT 86.260 150.520 87.860 150.820 ;
        RECT 80.900 150.080 81.820 150.420 ;
        RECT 84.860 150.080 85.780 150.420 ;
        RECT 80.900 148.320 81.820 148.660 ;
        RECT 84.860 148.320 85.780 148.660 ;
        RECT 80.900 147.440 81.820 147.780 ;
        RECT 84.860 146.560 85.780 146.900 ;
        RECT 84.860 145.680 85.780 146.020 ;
        RECT 86.260 145.540 86.560 150.520 ;
        RECT 86.940 150.480 87.860 150.520 ;
        RECT 86.860 145.540 87.780 145.580 ;
        RECT 86.260 145.240 87.780 145.540 ;
        RECT 80.900 143.340 81.820 143.380 ;
        RECT 77.980 143.040 81.820 143.340 ;
        RECT 84.860 143.040 85.780 143.380 ;
        RECT 72.180 143.000 73.100 143.040 ;
        RECT 80.820 143.000 81.740 143.040 ;
        RECT 72.100 142.160 73.020 142.500 ;
        RECT 80.900 142.160 81.820 142.500 ;
        RECT 65.980 142.020 66.900 142.060 ;
        RECT 87.020 142.020 87.940 142.060 ;
        RECT 88.240 142.020 88.540 154.040 ;
        RECT 65.380 141.720 66.980 142.020 ;
        RECT 61.740 141.680 62.660 141.720 ;
        RECT 66.060 141.680 66.980 141.720 ;
        RECT 86.940 141.720 88.540 142.020 ;
        RECT 90.580 159.320 92.100 159.620 ;
        RECT 90.580 154.340 90.880 159.320 ;
        RECT 91.180 155.800 92.100 156.140 ;
        RECT 92.560 154.780 92.860 175.160 ;
        RECT 93.340 174.720 94.260 175.060 ;
        RECT 97.300 174.720 98.220 175.060 ;
        RECT 93.340 173.840 94.260 174.180 ;
        RECT 97.300 173.840 98.220 174.180 ;
        RECT 93.340 171.200 94.260 171.540 ;
        RECT 93.340 170.320 94.260 170.660 ;
        RECT 97.300 170.320 98.220 170.660 ;
        RECT 94.835 168.210 95.175 169.130 ;
        RECT 97.300 168.860 98.220 168.900 ;
        RECT 98.680 168.860 98.980 192.760 ;
        RECT 97.300 168.560 98.980 168.860 ;
        RECT 93.340 167.680 94.260 168.020 ;
        RECT 97.300 167.680 98.220 168.020 ;
        RECT 93.340 166.800 94.260 167.140 ;
        RECT 97.300 166.800 98.220 167.140 ;
        RECT 93.340 164.160 94.260 164.500 ;
        RECT 93.340 163.280 94.260 163.620 ;
        RECT 97.300 163.280 98.220 163.620 ;
        RECT 93.340 160.640 94.260 160.980 ;
        RECT 97.300 160.640 98.220 160.980 ;
        RECT 99.460 159.320 100.380 159.660 ;
        RECT 93.340 155.360 94.260 155.700 ;
        RECT 97.300 155.360 98.220 155.700 ;
        RECT 93.340 154.780 94.260 154.820 ;
        RECT 92.560 154.480 94.260 154.780 ;
        RECT 91.180 154.340 92.100 154.380 ;
        RECT 90.580 154.040 92.100 154.340 ;
        RECT 90.580 142.020 90.880 154.040 ;
        RECT 91.340 150.820 92.260 150.860 ;
        RECT 91.260 150.520 92.860 150.820 ;
        RECT 91.260 150.480 92.180 150.520 ;
        RECT 91.340 145.540 92.260 145.580 ;
        RECT 92.560 145.540 92.860 150.520 ;
        RECT 93.340 150.080 94.260 150.420 ;
        RECT 97.300 150.080 98.220 150.420 ;
        RECT 93.340 148.320 94.260 148.660 ;
        RECT 97.300 148.320 98.220 148.660 ;
        RECT 97.300 147.440 98.220 147.780 ;
        RECT 93.340 146.560 94.260 146.900 ;
        RECT 93.340 145.680 94.260 146.020 ;
        RECT 91.340 145.240 92.860 145.540 ;
        RECT 93.340 143.040 94.260 143.380 ;
        RECT 97.300 143.340 98.220 143.380 ;
        RECT 100.840 143.340 101.140 196.280 ;
        RECT 97.300 143.040 101.140 143.340 ;
        RECT 103.180 196.280 104.860 196.580 ;
        RECT 103.180 143.340 103.480 196.280 ;
        RECT 106.100 195.840 107.020 196.180 ;
        RECT 110.060 195.840 110.980 196.180 ;
        RECT 110.060 195.260 110.980 195.300 ;
        RECT 111.460 195.260 111.760 201.560 ;
        RECT 116.380 198.340 117.300 198.380 ;
        RECT 117.760 198.340 118.060 202.000 ;
        RECT 118.540 199.360 119.460 199.700 ;
        RECT 122.500 199.360 123.420 199.700 ;
        RECT 140.920 199.050 141.220 214.590 ;
        RECT 143.680 214.150 144.600 214.490 ;
        RECT 143.680 213.570 144.600 213.610 ;
        RECT 145.060 213.570 145.360 218.550 ;
        RECT 149.020 216.650 149.320 220.310 ;
        RECT 149.800 216.650 150.720 216.690 ;
        RECT 149.020 216.350 150.720 216.650 ;
        RECT 147.640 215.910 148.560 216.250 ;
        RECT 147.640 215.030 148.560 215.370 ;
        RECT 143.680 213.270 145.360 213.570 ;
        RECT 149.800 213.130 150.720 213.170 ;
        RECT 149.800 212.830 151.480 213.130 ;
        RECT 149.800 211.370 150.720 211.410 ;
        RECT 149.020 211.070 150.720 211.370 ;
        RECT 143.680 210.630 144.600 210.970 ;
        RECT 147.640 210.630 148.560 210.970 ;
        RECT 147.640 210.050 148.560 210.090 ;
        RECT 149.020 210.050 149.320 211.070 ;
        RECT 147.640 209.750 149.320 210.050 ;
        RECT 141.520 209.610 142.440 209.650 ;
        RECT 141.520 209.310 143.200 209.610 ;
        RECT 142.900 208.290 143.200 209.310 ;
        RECT 143.680 208.870 144.600 209.210 ;
        RECT 147.640 208.870 148.560 209.210 ;
        RECT 143.680 208.290 144.600 208.330 ;
        RECT 142.900 207.990 144.600 208.290 ;
        RECT 149.020 206.090 149.320 209.750 ;
        RECT 149.800 207.850 150.720 207.890 ;
        RECT 151.180 207.850 151.480 212.830 ;
        RECT 149.800 207.550 151.480 207.850 ;
        RECT 149.800 206.090 150.720 206.130 ;
        RECT 149.020 205.790 150.720 206.090 ;
        RECT 143.680 205.350 144.600 205.690 ;
        RECT 147.640 205.350 148.560 205.690 ;
        RECT 141.520 204.330 142.440 204.370 ;
        RECT 141.520 204.030 142.600 204.330 ;
        RECT 142.300 203.730 143.200 204.030 ;
        RECT 142.900 199.490 143.200 203.730 ;
        RECT 143.680 201.830 144.600 202.170 ;
        RECT 147.640 201.830 148.560 202.170 ;
        RECT 143.680 200.070 144.600 200.410 ;
        RECT 147.640 200.070 148.560 200.410 ;
        RECT 143.680 199.490 144.600 199.530 ;
        RECT 142.900 199.190 144.600 199.490 ;
        RECT 147.640 199.190 148.560 199.530 ;
        RECT 141.520 199.050 142.440 199.090 ;
        RECT 140.920 198.750 142.440 199.050 ;
        RECT 110.060 194.960 111.760 195.260 ;
        RECT 115.780 198.040 118.060 198.340 ;
        RECT 112.060 194.520 112.980 194.860 ;
        RECT 103.940 193.060 104.860 193.100 ;
        RECT 103.940 192.760 105.640 193.060 ;
        RECT 105.340 168.860 105.640 192.760 ;
        RECT 106.100 192.320 107.020 192.660 ;
        RECT 110.060 192.320 110.980 192.660 ;
        RECT 106.100 191.440 107.020 191.780 ;
        RECT 110.060 191.440 110.980 191.780 ;
        RECT 112.060 191.000 112.980 191.340 ;
        RECT 110.060 188.800 110.980 189.140 ;
        RECT 106.100 187.920 107.020 188.260 ;
        RECT 110.060 187.920 110.980 188.260 ;
        RECT 115.780 186.020 116.080 198.040 ;
        RECT 118.540 197.600 119.460 197.940 ;
        RECT 122.500 197.600 123.420 197.940 ;
        RECT 147.640 197.730 148.560 197.770 ;
        RECT 151.180 197.730 151.480 207.550 ;
        RECT 147.640 197.430 151.480 197.730 ;
        RECT 143.680 196.550 144.600 196.890 ;
        RECT 147.640 196.550 148.560 196.890 ;
        RECT 147.640 195.970 148.560 196.010 ;
        RECT 147.640 195.670 149.320 195.970 ;
        RECT 143.680 194.790 144.600 195.130 ;
        RECT 147.640 194.790 148.560 195.130 ;
        RECT 143.680 194.210 144.600 194.250 ;
        RECT 143.680 193.910 145.360 194.210 ;
        RECT 141.520 193.470 142.440 193.810 ;
        RECT 141.520 190.250 142.440 190.290 ;
        RECT 140.920 189.950 142.440 190.250 ;
        RECT 116.540 187.780 117.460 187.820 ;
        RECT 116.540 187.480 118.060 187.780 ;
        RECT 116.380 186.020 117.300 186.060 ;
        RECT 115.780 185.720 117.300 186.020 ;
        RECT 110.060 185.280 110.980 185.620 ;
        RECT 106.100 184.400 107.020 184.740 ;
        RECT 110.060 184.400 110.980 184.740 ;
        RECT 107.470 182.290 107.810 183.210 ;
        RECT 106.100 181.760 107.020 182.100 ;
        RECT 110.060 181.760 110.980 182.100 ;
        RECT 106.100 180.880 107.020 181.220 ;
        RECT 110.060 180.880 110.980 181.220 ;
        RECT 110.060 178.240 110.980 178.580 ;
        RECT 106.100 177.360 107.020 177.700 ;
        RECT 110.060 177.360 110.980 177.700 ;
        RECT 108.345 175.250 108.685 176.170 ;
        RECT 112.220 175.460 113.140 175.500 ;
        RECT 111.460 175.160 113.140 175.460 ;
        RECT 106.100 174.720 107.020 175.060 ;
        RECT 110.060 174.720 110.980 175.060 ;
        RECT 106.100 173.840 107.020 174.180 ;
        RECT 110.060 173.840 110.980 174.180 ;
        RECT 110.060 171.200 110.980 171.540 ;
        RECT 106.100 170.320 107.020 170.660 ;
        RECT 110.060 170.320 110.980 170.660 ;
        RECT 106.100 168.860 107.020 168.900 ;
        RECT 105.340 168.560 107.020 168.860 ;
        RECT 109.145 168.210 109.485 169.130 ;
        RECT 106.100 167.680 107.020 168.020 ;
        RECT 110.060 167.680 110.980 168.020 ;
        RECT 106.100 166.800 107.020 167.140 ;
        RECT 110.060 166.800 110.980 167.140 ;
        RECT 110.060 164.160 110.980 164.500 ;
        RECT 106.100 163.280 107.020 163.620 ;
        RECT 110.060 163.280 110.980 163.620 ;
        RECT 106.100 160.640 107.020 160.980 ;
        RECT 110.060 160.640 110.980 160.980 ;
        RECT 103.780 159.320 104.700 159.660 ;
        RECT 106.100 155.360 107.020 155.700 ;
        RECT 110.060 155.360 110.980 155.700 ;
        RECT 110.060 154.780 110.980 154.820 ;
        RECT 111.460 154.780 111.760 175.160 ;
        RECT 112.140 168.080 113.060 168.420 ;
        RECT 112.220 159.620 113.140 159.660 ;
        RECT 112.220 159.320 113.740 159.620 ;
        RECT 112.060 155.800 112.980 156.140 ;
        RECT 110.060 154.480 111.760 154.780 ;
        RECT 112.220 154.340 113.140 154.380 ;
        RECT 113.440 154.340 113.740 159.320 ;
        RECT 112.220 154.040 113.740 154.340 ;
        RECT 112.060 150.820 112.980 150.860 ;
        RECT 111.460 150.520 113.060 150.820 ;
        RECT 106.100 150.080 107.020 150.420 ;
        RECT 110.060 150.080 110.980 150.420 ;
        RECT 106.100 148.320 107.020 148.660 ;
        RECT 110.060 148.320 110.980 148.660 ;
        RECT 106.100 147.440 107.020 147.780 ;
        RECT 110.060 146.560 110.980 146.900 ;
        RECT 110.060 145.680 110.980 146.020 ;
        RECT 111.460 145.540 111.760 150.520 ;
        RECT 112.140 150.480 113.060 150.520 ;
        RECT 112.060 145.540 112.980 145.580 ;
        RECT 111.460 145.240 112.980 145.540 ;
        RECT 106.100 143.340 107.020 143.380 ;
        RECT 103.180 143.040 107.020 143.340 ;
        RECT 110.060 143.040 110.980 143.380 ;
        RECT 97.380 143.000 98.300 143.040 ;
        RECT 106.020 143.000 106.940 143.040 ;
        RECT 97.300 142.160 98.220 142.500 ;
        RECT 106.100 142.160 107.020 142.500 ;
        RECT 91.180 142.020 92.100 142.060 ;
        RECT 112.220 142.020 113.140 142.060 ;
        RECT 113.440 142.020 113.740 154.040 ;
        RECT 90.580 141.720 92.180 142.020 ;
        RECT 86.940 141.680 87.860 141.720 ;
        RECT 91.260 141.680 92.180 141.720 ;
        RECT 112.140 141.720 113.740 142.020 ;
        RECT 115.780 142.020 116.080 185.720 ;
        RECT 116.380 182.500 117.460 182.540 ;
        RECT 117.760 182.500 118.060 187.480 ;
        RECT 122.500 186.160 123.420 186.500 ;
        RECT 118.540 185.280 119.460 185.620 ;
        RECT 122.500 184.400 123.420 184.740 ;
        RECT 116.380 182.200 118.060 182.500 ;
        RECT 122.500 181.760 123.420 182.100 ;
        RECT 122.500 180.880 123.420 181.220 ;
        RECT 122.500 180.300 123.420 180.340 ;
        RECT 122.500 180.000 124.180 180.300 ;
        RECT 122.500 178.240 123.420 178.580 ;
        RECT 122.500 177.360 123.420 177.700 ;
        RECT 122.500 174.720 123.420 175.060 ;
        RECT 122.500 173.840 123.420 174.180 ;
        RECT 118.540 172.960 119.460 173.300 ;
        RECT 118.540 172.080 119.460 172.420 ;
        RECT 122.500 172.080 123.420 172.420 ;
        RECT 122.500 170.320 123.420 170.660 ;
        RECT 118.540 169.440 119.460 169.780 ;
        RECT 122.500 169.440 123.420 169.780 ;
        RECT 118.540 168.560 119.460 168.900 ;
        RECT 122.500 168.560 123.420 168.900 ;
        RECT 118.620 166.990 119.540 167.330 ;
        RECT 123.880 166.660 124.180 180.000 ;
        RECT 124.660 176.920 125.580 177.260 ;
        RECT 140.920 174.410 141.220 189.950 ;
        RECT 143.680 189.510 144.600 189.850 ;
        RECT 143.680 188.930 144.600 188.970 ;
        RECT 145.060 188.930 145.360 193.910 ;
        RECT 149.020 192.010 149.320 195.670 ;
        RECT 149.800 192.010 150.720 192.050 ;
        RECT 149.020 191.710 150.720 192.010 ;
        RECT 147.640 191.270 148.560 191.610 ;
        RECT 147.640 190.390 148.560 190.730 ;
        RECT 143.680 188.630 145.360 188.930 ;
        RECT 149.800 188.490 150.720 188.530 ;
        RECT 149.800 188.190 151.480 188.490 ;
        RECT 149.800 186.730 150.720 186.770 ;
        RECT 149.020 186.430 150.720 186.730 ;
        RECT 143.680 185.990 144.600 186.330 ;
        RECT 147.640 185.990 148.560 186.330 ;
        RECT 147.640 185.410 148.560 185.450 ;
        RECT 149.020 185.410 149.320 186.430 ;
        RECT 147.640 185.110 149.320 185.410 ;
        RECT 141.520 184.970 142.440 185.010 ;
        RECT 141.520 184.670 143.200 184.970 ;
        RECT 142.900 183.650 143.200 184.670 ;
        RECT 143.680 184.230 144.600 184.570 ;
        RECT 147.640 184.230 148.560 184.570 ;
        RECT 143.680 183.650 144.600 183.690 ;
        RECT 142.900 183.350 144.600 183.650 ;
        RECT 149.020 181.450 149.320 185.110 ;
        RECT 149.800 183.210 150.720 183.250 ;
        RECT 151.180 183.210 151.480 188.190 ;
        RECT 149.800 182.910 151.480 183.210 ;
        RECT 149.800 181.450 150.720 181.490 ;
        RECT 149.020 181.150 150.720 181.450 ;
        RECT 143.680 180.710 144.600 181.050 ;
        RECT 147.640 180.710 148.560 181.050 ;
        RECT 141.520 179.690 142.440 179.730 ;
        RECT 141.520 179.390 142.600 179.690 ;
        RECT 142.300 179.090 143.200 179.390 ;
        RECT 142.900 174.850 143.200 179.090 ;
        RECT 143.680 177.190 144.600 177.530 ;
        RECT 147.640 177.190 148.560 177.530 ;
        RECT 143.680 175.430 144.600 175.770 ;
        RECT 147.640 175.430 148.560 175.770 ;
        RECT 143.680 174.850 144.600 174.890 ;
        RECT 142.900 174.550 144.600 174.850 ;
        RECT 147.640 174.550 148.560 174.890 ;
        RECT 141.520 174.410 142.440 174.450 ;
        RECT 140.920 174.110 142.440 174.410 ;
        RECT 147.640 173.090 148.560 173.130 ;
        RECT 151.180 173.090 151.480 182.910 ;
        RECT 147.640 172.790 151.480 173.090 ;
        RECT 143.680 171.910 144.600 172.250 ;
        RECT 147.640 171.910 148.560 172.250 ;
        RECT 147.640 171.330 148.560 171.370 ;
        RECT 147.640 171.030 149.320 171.330 ;
        RECT 143.680 170.150 144.600 170.490 ;
        RECT 147.640 170.150 148.560 170.490 ;
        RECT 143.680 169.570 144.600 169.610 ;
        RECT 143.680 169.270 145.360 169.570 ;
        RECT 141.520 168.830 142.440 169.170 ;
        RECT 124.660 166.660 125.580 166.700 ;
        RECT 123.880 166.360 125.580 166.660 ;
        RECT 118.540 165.920 119.460 166.260 ;
        RECT 122.500 165.920 123.420 166.260 ;
        RECT 122.500 165.040 123.420 165.380 ;
        RECT 123.880 163.140 124.180 166.360 ;
        RECT 141.520 165.610 142.440 165.650 ;
        RECT 140.920 165.310 142.440 165.610 ;
        RECT 124.660 163.140 125.580 163.180 ;
        RECT 123.880 162.840 125.580 163.140 ;
        RECT 122.500 162.400 123.420 162.740 ;
        RECT 122.500 161.520 123.420 161.860 ;
        RECT 122.500 158.880 123.420 159.220 ;
        RECT 122.500 158.000 123.420 158.340 ;
        RECT 124.660 157.560 125.580 157.900 ;
        RECT 116.540 156.100 117.460 156.140 ;
        RECT 116.540 155.800 118.060 156.100 ;
        RECT 116.380 150.820 117.460 150.860 ;
        RECT 117.760 150.820 118.060 155.800 ;
        RECT 122.500 155.360 123.420 155.700 ;
        RECT 122.500 154.480 123.420 154.820 ;
        RECT 118.540 153.600 119.460 153.940 ;
        RECT 116.380 150.520 118.060 150.820 ;
        RECT 140.920 149.770 141.220 165.310 ;
        RECT 143.680 164.870 144.600 165.210 ;
        RECT 143.680 164.290 144.600 164.330 ;
        RECT 145.060 164.290 145.360 169.270 ;
        RECT 149.020 167.370 149.320 171.030 ;
        RECT 149.800 167.370 150.720 167.410 ;
        RECT 149.020 167.070 150.720 167.370 ;
        RECT 147.640 166.630 148.560 166.970 ;
        RECT 147.640 165.750 148.560 166.090 ;
        RECT 143.680 163.990 145.360 164.290 ;
        RECT 149.800 163.850 150.720 163.890 ;
        RECT 149.800 163.550 151.480 163.850 ;
        RECT 149.800 162.090 150.720 162.130 ;
        RECT 149.020 161.790 150.720 162.090 ;
        RECT 143.680 161.350 144.600 161.690 ;
        RECT 147.640 161.350 148.560 161.690 ;
        RECT 147.640 160.770 148.560 160.810 ;
        RECT 149.020 160.770 149.320 161.790 ;
        RECT 147.640 160.470 149.320 160.770 ;
        RECT 141.520 160.330 142.440 160.370 ;
        RECT 141.520 160.030 143.200 160.330 ;
        RECT 142.900 159.010 143.200 160.030 ;
        RECT 143.680 159.590 144.600 159.930 ;
        RECT 147.640 159.590 148.560 159.930 ;
        RECT 143.680 159.010 144.600 159.050 ;
        RECT 142.900 158.710 144.600 159.010 ;
        RECT 149.020 156.810 149.320 160.470 ;
        RECT 149.800 158.570 150.720 158.610 ;
        RECT 151.180 158.570 151.480 163.550 ;
        RECT 149.800 158.270 151.480 158.570 ;
        RECT 149.800 156.810 150.720 156.850 ;
        RECT 149.020 156.510 150.720 156.810 ;
        RECT 143.680 156.070 144.600 156.410 ;
        RECT 147.640 156.070 148.560 156.410 ;
        RECT 141.520 155.050 142.440 155.090 ;
        RECT 141.520 154.750 142.600 155.050 ;
        RECT 142.300 154.450 143.200 154.750 ;
        RECT 142.900 150.210 143.200 154.450 ;
        RECT 143.680 152.550 144.600 152.890 ;
        RECT 147.640 152.550 148.560 152.890 ;
        RECT 143.680 150.790 144.600 151.130 ;
        RECT 147.640 150.790 148.560 151.130 ;
        RECT 143.680 150.210 144.600 150.250 ;
        RECT 142.900 149.910 144.600 150.210 ;
        RECT 147.640 149.910 148.560 150.250 ;
        RECT 141.520 149.770 142.440 149.810 ;
        RECT 140.920 149.470 142.440 149.770 ;
        RECT 147.640 148.450 148.560 148.490 ;
        RECT 151.180 148.450 151.480 158.270 ;
        RECT 147.640 148.150 151.480 148.450 ;
        RECT 143.680 147.270 144.600 147.610 ;
        RECT 147.640 147.270 148.560 147.610 ;
        RECT 147.640 146.690 148.560 146.730 ;
        RECT 147.640 146.390 149.320 146.690 ;
        RECT 143.680 145.510 144.600 145.850 ;
        RECT 147.640 145.510 148.560 145.850 ;
        RECT 143.680 144.930 144.600 144.970 ;
        RECT 143.680 144.630 145.360 144.930 ;
        RECT 141.520 144.190 142.440 144.530 ;
        RECT 122.500 142.160 123.420 142.500 ;
        RECT 116.380 142.020 117.300 142.060 ;
        RECT 115.780 141.720 117.300 142.020 ;
        RECT 112.140 141.680 113.060 141.720 ;
        RECT 118.540 141.280 119.460 141.620 ;
        RECT 141.520 140.970 142.440 141.010 ;
        RECT 17.740 140.400 18.660 140.740 ;
        RECT 21.700 140.400 22.620 140.740 ;
        RECT 30.500 140.400 31.420 140.740 ;
        RECT 34.460 140.400 35.380 140.740 ;
        RECT 42.940 140.400 43.860 140.740 ;
        RECT 46.900 140.400 47.820 140.740 ;
        RECT 55.700 140.400 56.620 140.740 ;
        RECT 59.660 140.400 60.580 140.740 ;
        RECT 68.140 140.400 69.060 140.740 ;
        RECT 72.100 140.400 73.020 140.740 ;
        RECT 80.900 140.400 81.820 140.740 ;
        RECT 84.860 140.400 85.780 140.740 ;
        RECT 93.340 140.400 94.260 140.740 ;
        RECT 97.300 140.400 98.220 140.740 ;
        RECT 106.100 140.400 107.020 140.740 ;
        RECT 110.060 140.400 110.980 140.740 ;
        RECT 118.540 140.400 119.460 140.740 ;
        RECT 122.500 140.400 123.420 140.740 ;
        RECT 140.920 140.670 142.440 140.970 ;
        RECT 17.740 139.520 18.660 139.860 ;
        RECT 21.700 139.520 22.620 139.860 ;
        RECT 30.500 139.520 31.420 139.860 ;
        RECT 34.460 139.520 35.380 139.860 ;
        RECT 42.940 139.520 43.860 139.860 ;
        RECT 46.900 139.520 47.820 139.860 ;
        RECT 55.700 139.520 56.620 139.860 ;
        RECT 59.660 139.520 60.580 139.860 ;
        RECT 68.140 139.520 69.060 139.860 ;
        RECT 72.100 139.520 73.020 139.860 ;
        RECT 80.900 139.520 81.820 139.860 ;
        RECT 84.860 139.520 85.780 139.860 ;
        RECT 93.340 139.520 94.260 139.860 ;
        RECT 97.300 139.520 98.220 139.860 ;
        RECT 106.100 139.520 107.020 139.860 ;
        RECT 110.060 139.520 110.980 139.860 ;
        RECT 118.540 139.520 119.460 139.860 ;
        RECT 122.500 139.520 123.420 139.860 ;
        RECT 72.020 135.350 72.360 135.960 ;
        RECT 72.020 135.040 72.440 135.350 ;
        RECT 65.120 128.560 65.460 129.170 ;
        RECT 65.120 128.250 65.540 128.560 ;
        RECT 63.320 127.590 63.660 128.200 ;
        RECT 63.320 127.280 63.740 127.590 ;
        RECT 61.520 126.620 61.860 127.230 ;
        RECT 61.520 126.310 61.940 126.620 ;
        RECT 60.620 119.830 60.960 120.440 ;
        RECT 60.620 119.520 61.040 119.830 ;
        RECT 12.240 110.130 58.120 110.510 ;
        RECT 8.640 93.110 9.560 94.030 ;
        RECT 12.240 93.190 12.620 110.130 ;
        RECT 12.940 93.190 13.320 110.130 ;
        RECT 13.640 97.870 14.020 110.130 ;
        RECT 13.680 96.570 14.020 97.490 ;
        RECT 13.640 93.190 14.020 96.270 ;
        RECT 14.340 93.190 14.720 110.130 ;
        RECT 15.040 97.870 15.420 110.130 ;
        RECT 15.080 96.570 15.420 97.490 ;
        RECT 15.040 93.190 15.420 96.270 ;
        RECT 15.740 93.190 16.120 110.130 ;
        RECT 16.440 97.870 16.820 110.130 ;
        RECT 16.480 96.570 16.820 97.490 ;
        RECT 16.440 93.190 16.820 96.270 ;
        RECT 17.140 93.190 17.520 110.130 ;
        RECT 17.840 97.870 18.220 110.130 ;
        RECT 17.880 96.570 18.220 97.490 ;
        RECT 17.840 93.190 18.220 96.270 ;
        RECT 18.540 93.190 18.920 110.130 ;
        RECT 19.240 103.990 19.620 110.130 ;
        RECT 19.280 102.690 19.620 103.610 ;
        RECT 19.240 93.190 19.620 102.390 ;
        RECT 19.940 93.190 20.320 110.130 ;
        RECT 20.640 103.990 21.020 110.130 ;
        RECT 20.680 102.690 21.020 103.610 ;
        RECT 20.640 93.190 21.020 102.390 ;
        RECT 21.340 93.190 21.720 110.130 ;
        RECT 22.040 107.050 22.420 110.130 ;
        RECT 22.080 105.750 22.420 106.670 ;
        RECT 22.040 93.190 22.420 105.450 ;
        RECT 22.740 93.190 23.120 110.130 ;
        RECT 23.480 108.810 23.820 109.730 ;
        RECT 23.440 93.190 23.820 108.510 ;
        RECT 24.140 93.190 24.520 110.130 ;
        RECT 24.840 100.930 25.220 110.130 ;
        RECT 24.880 99.630 25.220 100.550 ;
        RECT 24.840 93.190 25.220 99.330 ;
        RECT 25.540 93.190 25.920 110.130 ;
        RECT 26.240 107.050 26.620 110.130 ;
        RECT 26.280 105.750 26.620 106.670 ;
        RECT 26.240 93.190 26.620 105.450 ;
        RECT 26.940 93.190 27.320 110.130 ;
        RECT 27.640 103.990 28.020 110.130 ;
        RECT 27.680 102.690 28.020 103.610 ;
        RECT 27.640 93.190 28.020 102.390 ;
        RECT 28.340 93.190 28.720 110.130 ;
        RECT 29.040 103.990 29.420 110.130 ;
        RECT 29.080 102.690 29.420 103.610 ;
        RECT 29.040 93.190 29.420 102.390 ;
        RECT 29.740 93.190 30.120 110.130 ;
        RECT 30.440 97.870 30.820 110.130 ;
        RECT 30.480 96.570 30.820 97.490 ;
        RECT 30.440 93.190 30.820 96.270 ;
        RECT 31.140 93.190 31.520 110.130 ;
        RECT 31.840 97.870 32.220 110.130 ;
        RECT 31.880 96.570 32.220 97.490 ;
        RECT 31.840 93.190 32.220 96.270 ;
        RECT 32.540 93.190 32.920 110.130 ;
        RECT 33.240 97.870 33.620 110.130 ;
        RECT 33.280 96.570 33.620 97.490 ;
        RECT 33.240 93.190 33.620 96.270 ;
        RECT 33.940 93.190 34.320 110.130 ;
        RECT 34.640 97.870 35.020 110.130 ;
        RECT 34.680 96.570 35.020 97.490 ;
        RECT 34.640 93.190 35.020 96.270 ;
        RECT 35.340 93.190 35.720 110.130 ;
        RECT 36.040 97.870 36.420 110.130 ;
        RECT 36.080 96.570 36.420 97.490 ;
        RECT 36.040 93.190 36.420 96.270 ;
        RECT 36.740 93.190 37.120 110.130 ;
        RECT 37.440 97.870 37.820 110.130 ;
        RECT 37.480 96.570 37.820 97.490 ;
        RECT 37.440 93.190 37.820 96.270 ;
        RECT 38.140 93.190 38.520 110.130 ;
        RECT 38.840 97.870 39.220 110.130 ;
        RECT 38.880 96.570 39.220 97.490 ;
        RECT 38.840 93.190 39.220 96.270 ;
        RECT 39.540 93.190 39.920 110.130 ;
        RECT 40.240 97.870 40.620 110.130 ;
        RECT 40.280 96.570 40.620 97.490 ;
        RECT 40.240 93.190 40.620 96.270 ;
        RECT 40.940 93.190 41.320 110.130 ;
        RECT 41.640 103.990 42.020 110.130 ;
        RECT 41.680 102.690 42.020 103.610 ;
        RECT 41.640 93.190 42.020 102.390 ;
        RECT 42.340 93.190 42.720 110.130 ;
        RECT 43.040 103.990 43.420 110.130 ;
        RECT 43.080 102.690 43.420 103.610 ;
        RECT 43.040 93.190 43.420 102.390 ;
        RECT 43.740 93.190 44.120 110.130 ;
        RECT 44.440 107.050 44.820 110.130 ;
        RECT 44.480 105.750 44.820 106.670 ;
        RECT 44.440 93.190 44.820 105.450 ;
        RECT 45.140 93.190 45.520 110.130 ;
        RECT 45.840 100.930 46.220 110.130 ;
        RECT 45.880 99.630 46.220 100.550 ;
        RECT 45.840 93.190 46.220 99.330 ;
        RECT 46.540 93.190 46.920 110.130 ;
        RECT 47.240 94.810 47.620 110.130 ;
        RECT 47.280 93.510 47.620 94.430 ;
        RECT 47.940 93.190 48.320 110.130 ;
        RECT 48.640 107.050 49.020 110.130 ;
        RECT 48.680 105.750 49.020 106.670 ;
        RECT 48.640 93.190 49.020 105.450 ;
        RECT 49.340 93.190 49.720 110.130 ;
        RECT 50.040 103.990 50.420 110.130 ;
        RECT 50.080 102.690 50.420 103.610 ;
        RECT 50.040 93.190 50.420 102.390 ;
        RECT 50.740 93.190 51.120 110.130 ;
        RECT 51.440 103.990 51.820 110.130 ;
        RECT 51.480 102.690 51.820 103.610 ;
        RECT 51.440 93.190 51.820 102.390 ;
        RECT 52.140 93.190 52.520 110.130 ;
        RECT 52.840 97.870 53.220 110.130 ;
        RECT 52.880 96.570 53.220 97.490 ;
        RECT 52.840 93.190 53.220 96.270 ;
        RECT 53.540 93.190 53.920 110.130 ;
        RECT 54.240 97.870 54.620 110.130 ;
        RECT 54.280 96.570 54.620 97.490 ;
        RECT 54.240 93.190 54.620 96.270 ;
        RECT 54.940 93.190 55.320 110.130 ;
        RECT 55.640 97.870 56.020 110.130 ;
        RECT 55.680 96.570 56.020 97.490 ;
        RECT 55.640 93.190 56.020 96.270 ;
        RECT 56.340 93.190 56.720 110.130 ;
        RECT 57.040 97.870 57.420 110.130 ;
        RECT 57.080 96.570 57.420 97.490 ;
        RECT 57.040 93.190 57.420 96.270 ;
        RECT 57.740 93.190 58.120 110.130 ;
        RECT 60.660 110.210 61.040 119.520 ;
        RECT 61.560 110.210 61.940 126.310 ;
        RECT 62.420 120.800 62.760 121.410 ;
        RECT 62.420 120.490 62.840 120.800 ;
        RECT 62.460 110.210 62.840 120.490 ;
        RECT 63.360 110.210 63.740 127.280 ;
        RECT 64.220 121.770 64.560 122.380 ;
        RECT 64.220 121.460 64.640 121.770 ;
        RECT 64.260 110.210 64.640 121.460 ;
        RECT 65.160 110.210 65.540 128.250 ;
        RECT 68.720 125.650 69.060 126.260 ;
        RECT 68.720 125.340 69.140 125.650 ;
        RECT 67.820 124.680 68.160 125.290 ;
        RECT 67.820 124.370 68.240 124.680 ;
        RECT 66.920 123.710 67.260 124.320 ;
        RECT 66.920 123.400 67.340 123.710 ;
        RECT 66.020 122.740 66.360 123.350 ;
        RECT 66.020 122.430 66.440 122.740 ;
        RECT 66.060 110.210 66.440 122.430 ;
        RECT 66.960 110.210 67.340 123.400 ;
        RECT 67.860 110.210 68.240 124.370 ;
        RECT 68.760 110.210 69.140 125.340 ;
        RECT 72.060 110.210 72.440 135.040 ;
        RECT 72.920 134.380 73.260 134.990 ;
        RECT 72.920 134.070 73.340 134.380 ;
        RECT 72.960 110.210 73.340 134.070 ;
        RECT 73.820 133.410 74.160 134.020 ;
        RECT 73.820 133.100 74.240 133.410 ;
        RECT 73.860 110.210 74.240 133.100 ;
        RECT 74.720 132.440 75.060 133.050 ;
        RECT 74.720 132.130 75.140 132.440 ;
        RECT 74.760 110.210 75.140 132.130 ;
        RECT 75.620 131.470 75.960 132.080 ;
        RECT 75.620 131.160 76.040 131.470 ;
        RECT 75.660 110.210 76.040 131.160 ;
        RECT 77.420 130.500 77.760 131.110 ;
        RECT 77.420 130.190 77.840 130.500 ;
        RECT 76.520 118.860 76.860 119.470 ;
        RECT 76.520 118.550 76.940 118.860 ;
        RECT 76.560 110.210 76.940 118.550 ;
        RECT 77.460 110.210 77.840 130.190 ;
        RECT 79.220 129.530 79.560 130.140 ;
        RECT 79.220 129.220 79.640 129.530 ;
        RECT 78.320 117.890 78.660 118.500 ;
        RECT 78.320 117.580 78.740 117.890 ;
        RECT 78.360 110.210 78.740 117.580 ;
        RECT 79.260 110.210 79.640 129.220 ;
        RECT 140.920 125.130 141.220 140.670 ;
        RECT 143.680 140.230 144.600 140.570 ;
        RECT 143.680 139.650 144.600 139.690 ;
        RECT 145.060 139.650 145.360 144.630 ;
        RECT 149.020 142.730 149.320 146.390 ;
        RECT 149.800 142.730 150.720 142.770 ;
        RECT 149.020 142.430 150.720 142.730 ;
        RECT 147.640 141.990 148.560 142.330 ;
        RECT 147.640 141.110 148.560 141.450 ;
        RECT 143.680 139.350 145.360 139.650 ;
        RECT 149.800 139.210 150.720 139.250 ;
        RECT 149.800 138.910 151.480 139.210 ;
        RECT 149.800 137.450 150.720 137.490 ;
        RECT 149.020 137.150 150.720 137.450 ;
        RECT 143.680 136.710 144.600 137.050 ;
        RECT 147.640 136.710 148.560 137.050 ;
        RECT 147.640 136.130 148.560 136.170 ;
        RECT 149.020 136.130 149.320 137.150 ;
        RECT 147.640 135.830 149.320 136.130 ;
        RECT 141.520 135.690 142.440 135.730 ;
        RECT 141.520 135.390 143.200 135.690 ;
        RECT 142.900 134.370 143.200 135.390 ;
        RECT 143.680 134.950 144.600 135.290 ;
        RECT 147.640 134.950 148.560 135.290 ;
        RECT 143.680 134.370 144.600 134.410 ;
        RECT 142.900 134.070 144.600 134.370 ;
        RECT 149.020 132.170 149.320 135.830 ;
        RECT 149.800 133.930 150.720 133.970 ;
        RECT 151.180 133.930 151.480 138.910 ;
        RECT 149.800 133.630 151.480 133.930 ;
        RECT 149.800 132.170 150.720 132.210 ;
        RECT 149.020 131.870 150.720 132.170 ;
        RECT 143.680 131.430 144.600 131.770 ;
        RECT 147.640 131.430 148.560 131.770 ;
        RECT 141.520 130.410 142.440 130.450 ;
        RECT 141.520 130.110 142.600 130.410 ;
        RECT 142.300 129.810 143.200 130.110 ;
        RECT 142.900 125.570 143.200 129.810 ;
        RECT 143.680 127.910 144.600 128.250 ;
        RECT 147.640 127.910 148.560 128.250 ;
        RECT 143.680 126.150 144.600 126.490 ;
        RECT 147.640 126.150 148.560 126.490 ;
        RECT 143.680 125.570 144.600 125.610 ;
        RECT 142.900 125.270 144.600 125.570 ;
        RECT 147.640 125.270 148.560 125.610 ;
        RECT 141.520 125.130 142.440 125.170 ;
        RECT 140.920 124.830 142.440 125.130 ;
        RECT 147.640 123.810 148.560 123.850 ;
        RECT 151.180 123.810 151.480 133.630 ;
        RECT 147.640 123.510 151.480 123.810 ;
        RECT 143.680 122.630 144.600 122.970 ;
        RECT 147.640 122.630 148.560 122.970 ;
        RECT 147.640 122.050 148.560 122.090 ;
        RECT 147.640 121.750 149.320 122.050 ;
        RECT 143.680 120.870 144.600 121.210 ;
        RECT 147.640 120.870 148.560 121.210 ;
        RECT 143.680 120.290 144.600 120.330 ;
        RECT 143.680 119.990 145.360 120.290 ;
        RECT 141.520 119.550 142.440 119.890 ;
        RECT 80.120 116.920 80.460 117.530 ;
        RECT 80.120 116.610 80.540 116.920 ;
        RECT 80.160 110.210 80.540 116.610 ;
        RECT 141.520 116.330 142.440 116.370 ;
        RECT 140.920 116.030 142.440 116.330 ;
        RECT 60.660 109.730 60.960 110.210 ;
        RECT 58.840 109.120 59.760 109.460 ;
        RECT 60.660 108.810 61.000 109.730 ;
        RECT 60.660 106.670 60.960 108.810 ;
        RECT 58.840 106.060 59.760 106.400 ;
        RECT 60.660 105.750 61.000 106.670 ;
        RECT 60.660 103.610 60.960 105.750 ;
        RECT 58.840 103.000 59.760 103.340 ;
        RECT 60.660 102.690 61.000 103.610 ;
        RECT 60.660 100.550 60.960 102.690 ;
        RECT 58.840 99.940 59.760 100.280 ;
        RECT 60.660 99.630 61.000 100.550 ;
        RECT 60.660 97.490 60.960 99.630 ;
        RECT 58.840 96.880 59.760 97.220 ;
        RECT 60.660 96.570 61.000 97.490 ;
        RECT 60.660 94.430 60.960 96.570 ;
        RECT 58.840 93.820 59.760 94.160 ;
        RECT 60.660 93.510 61.000 94.430 ;
        RECT 12.240 93.110 58.120 93.190 ;
        RECT 8.640 92.810 58.120 93.110 ;
        RECT 12.240 92.730 58.120 92.810 ;
        RECT 8.640 75.710 9.560 76.630 ;
        RECT 12.240 75.790 12.620 92.730 ;
        RECT 12.940 75.790 13.320 92.730 ;
        RECT 13.640 80.470 14.020 92.730 ;
        RECT 13.680 79.170 14.020 80.090 ;
        RECT 13.640 75.790 14.020 78.870 ;
        RECT 14.340 75.790 14.720 92.730 ;
        RECT 15.040 80.470 15.420 92.730 ;
        RECT 15.080 79.170 15.420 80.090 ;
        RECT 15.040 75.790 15.420 78.870 ;
        RECT 15.740 75.790 16.120 92.730 ;
        RECT 16.440 80.470 16.820 92.730 ;
        RECT 16.480 79.170 16.820 80.090 ;
        RECT 16.440 75.790 16.820 78.870 ;
        RECT 17.140 75.790 17.520 92.730 ;
        RECT 17.840 80.470 18.220 92.730 ;
        RECT 17.880 79.170 18.220 80.090 ;
        RECT 17.840 75.790 18.220 78.870 ;
        RECT 18.540 75.790 18.920 92.730 ;
        RECT 19.240 86.590 19.620 92.730 ;
        RECT 19.280 85.290 19.620 86.210 ;
        RECT 19.240 75.790 19.620 84.990 ;
        RECT 19.940 75.790 20.320 92.730 ;
        RECT 20.640 86.590 21.020 92.730 ;
        RECT 20.680 85.290 21.020 86.210 ;
        RECT 20.640 75.790 21.020 84.990 ;
        RECT 21.340 75.790 21.720 92.730 ;
        RECT 22.040 89.650 22.420 92.730 ;
        RECT 22.080 88.350 22.420 89.270 ;
        RECT 22.040 75.790 22.420 88.050 ;
        RECT 22.740 75.790 23.120 92.730 ;
        RECT 23.480 91.410 23.820 92.330 ;
        RECT 23.440 75.790 23.820 91.110 ;
        RECT 24.140 75.790 24.520 92.730 ;
        RECT 24.840 83.530 25.220 92.730 ;
        RECT 24.880 82.230 25.220 83.150 ;
        RECT 24.840 75.790 25.220 81.930 ;
        RECT 25.540 75.790 25.920 92.730 ;
        RECT 26.240 89.650 26.620 92.730 ;
        RECT 26.280 88.350 26.620 89.270 ;
        RECT 26.240 75.790 26.620 88.050 ;
        RECT 26.940 75.790 27.320 92.730 ;
        RECT 27.640 86.590 28.020 92.730 ;
        RECT 27.680 85.290 28.020 86.210 ;
        RECT 27.640 75.790 28.020 84.990 ;
        RECT 28.340 75.790 28.720 92.730 ;
        RECT 29.040 86.590 29.420 92.730 ;
        RECT 29.080 85.290 29.420 86.210 ;
        RECT 29.040 75.790 29.420 84.990 ;
        RECT 29.740 75.790 30.120 92.730 ;
        RECT 30.440 80.470 30.820 92.730 ;
        RECT 30.480 79.170 30.820 80.090 ;
        RECT 30.440 75.790 30.820 78.870 ;
        RECT 31.140 75.790 31.520 92.730 ;
        RECT 31.840 80.470 32.220 92.730 ;
        RECT 31.880 79.170 32.220 80.090 ;
        RECT 31.840 75.790 32.220 78.870 ;
        RECT 32.540 75.790 32.920 92.730 ;
        RECT 33.240 80.470 33.620 92.730 ;
        RECT 33.280 79.170 33.620 80.090 ;
        RECT 33.240 75.790 33.620 78.870 ;
        RECT 33.940 75.790 34.320 92.730 ;
        RECT 34.640 80.470 35.020 92.730 ;
        RECT 34.680 79.170 35.020 80.090 ;
        RECT 34.640 75.790 35.020 78.870 ;
        RECT 35.340 75.790 35.720 92.730 ;
        RECT 36.040 80.470 36.420 92.730 ;
        RECT 36.080 79.170 36.420 80.090 ;
        RECT 36.040 75.790 36.420 78.870 ;
        RECT 36.740 75.790 37.120 92.730 ;
        RECT 37.440 80.470 37.820 92.730 ;
        RECT 37.480 79.170 37.820 80.090 ;
        RECT 37.440 75.790 37.820 78.870 ;
        RECT 38.140 75.790 38.520 92.730 ;
        RECT 38.840 80.470 39.220 92.730 ;
        RECT 38.880 79.170 39.220 80.090 ;
        RECT 38.840 75.790 39.220 78.870 ;
        RECT 39.540 75.790 39.920 92.730 ;
        RECT 40.240 80.470 40.620 92.730 ;
        RECT 40.280 79.170 40.620 80.090 ;
        RECT 40.240 75.790 40.620 78.870 ;
        RECT 40.940 75.790 41.320 92.730 ;
        RECT 41.640 86.590 42.020 92.730 ;
        RECT 41.680 85.290 42.020 86.210 ;
        RECT 41.640 75.790 42.020 84.990 ;
        RECT 42.340 75.790 42.720 92.730 ;
        RECT 43.040 86.590 43.420 92.730 ;
        RECT 43.080 85.290 43.420 86.210 ;
        RECT 43.040 75.790 43.420 84.990 ;
        RECT 43.740 75.790 44.120 92.730 ;
        RECT 44.440 89.650 44.820 92.730 ;
        RECT 44.480 88.350 44.820 89.270 ;
        RECT 44.440 75.790 44.820 88.050 ;
        RECT 45.140 75.790 45.520 92.730 ;
        RECT 45.840 83.530 46.220 92.730 ;
        RECT 45.880 82.230 46.220 83.150 ;
        RECT 45.840 75.790 46.220 81.930 ;
        RECT 46.540 75.790 46.920 92.730 ;
        RECT 47.240 77.410 47.620 92.730 ;
        RECT 47.280 76.110 47.620 77.030 ;
        RECT 47.940 75.790 48.320 92.730 ;
        RECT 48.640 89.650 49.020 92.730 ;
        RECT 48.680 88.350 49.020 89.270 ;
        RECT 48.640 75.790 49.020 88.050 ;
        RECT 49.340 75.790 49.720 92.730 ;
        RECT 50.040 86.590 50.420 92.730 ;
        RECT 50.080 85.290 50.420 86.210 ;
        RECT 50.040 75.790 50.420 84.990 ;
        RECT 50.740 75.790 51.120 92.730 ;
        RECT 51.440 86.590 51.820 92.730 ;
        RECT 51.480 85.290 51.820 86.210 ;
        RECT 51.440 75.790 51.820 84.990 ;
        RECT 52.140 75.790 52.520 92.730 ;
        RECT 52.840 80.470 53.220 92.730 ;
        RECT 52.880 79.170 53.220 80.090 ;
        RECT 52.840 75.790 53.220 78.870 ;
        RECT 53.540 75.790 53.920 92.730 ;
        RECT 54.240 80.470 54.620 92.730 ;
        RECT 54.280 79.170 54.620 80.090 ;
        RECT 54.240 75.790 54.620 78.870 ;
        RECT 54.940 75.790 55.320 92.730 ;
        RECT 55.640 80.470 56.020 92.730 ;
        RECT 55.680 79.170 56.020 80.090 ;
        RECT 55.640 75.790 56.020 78.870 ;
        RECT 56.340 75.790 56.720 92.730 ;
        RECT 57.040 80.470 57.420 92.730 ;
        RECT 57.080 79.170 57.420 80.090 ;
        RECT 57.040 75.790 57.420 78.870 ;
        RECT 57.740 75.790 58.120 92.730 ;
        RECT 58.840 91.720 59.760 92.060 ;
        RECT 58.840 88.660 59.760 89.000 ;
        RECT 58.840 85.600 59.760 85.940 ;
        RECT 58.840 82.540 59.760 82.880 ;
        RECT 58.840 79.480 59.760 79.820 ;
        RECT 58.840 76.420 59.760 76.760 ;
        RECT 12.240 75.710 58.120 75.790 ;
        RECT 8.640 75.410 58.120 75.710 ;
        RECT 12.240 75.330 58.120 75.410 ;
        RECT 8.640 58.310 9.560 59.230 ;
        RECT 12.240 58.390 12.620 75.330 ;
        RECT 12.940 58.390 13.320 75.330 ;
        RECT 13.640 63.070 14.020 75.330 ;
        RECT 13.680 61.770 14.020 62.690 ;
        RECT 13.640 58.390 14.020 61.470 ;
        RECT 14.340 58.390 14.720 75.330 ;
        RECT 15.040 63.070 15.420 75.330 ;
        RECT 15.080 61.770 15.420 62.690 ;
        RECT 15.040 58.390 15.420 61.470 ;
        RECT 15.740 58.390 16.120 75.330 ;
        RECT 16.440 63.070 16.820 75.330 ;
        RECT 16.480 61.770 16.820 62.690 ;
        RECT 16.440 58.390 16.820 61.470 ;
        RECT 17.140 58.390 17.520 75.330 ;
        RECT 17.840 63.070 18.220 75.330 ;
        RECT 17.880 61.770 18.220 62.690 ;
        RECT 17.840 58.390 18.220 61.470 ;
        RECT 18.540 58.390 18.920 75.330 ;
        RECT 19.240 69.190 19.620 75.330 ;
        RECT 19.280 67.890 19.620 68.810 ;
        RECT 19.240 58.390 19.620 67.590 ;
        RECT 19.940 58.390 20.320 75.330 ;
        RECT 20.640 69.190 21.020 75.330 ;
        RECT 20.680 67.890 21.020 68.810 ;
        RECT 20.640 58.390 21.020 67.590 ;
        RECT 21.340 58.390 21.720 75.330 ;
        RECT 22.040 72.250 22.420 75.330 ;
        RECT 22.080 70.950 22.420 71.870 ;
        RECT 22.040 58.390 22.420 70.650 ;
        RECT 22.740 58.390 23.120 75.330 ;
        RECT 23.480 74.010 23.820 74.930 ;
        RECT 23.440 58.390 23.820 73.710 ;
        RECT 24.140 58.390 24.520 75.330 ;
        RECT 24.840 66.130 25.220 75.330 ;
        RECT 24.880 64.830 25.220 65.750 ;
        RECT 24.840 58.390 25.220 64.530 ;
        RECT 25.540 58.390 25.920 75.330 ;
        RECT 26.240 72.250 26.620 75.330 ;
        RECT 26.280 70.950 26.620 71.870 ;
        RECT 26.240 58.390 26.620 70.650 ;
        RECT 26.940 58.390 27.320 75.330 ;
        RECT 27.640 69.190 28.020 75.330 ;
        RECT 27.680 67.890 28.020 68.810 ;
        RECT 27.640 58.390 28.020 67.590 ;
        RECT 28.340 58.390 28.720 75.330 ;
        RECT 29.040 69.190 29.420 75.330 ;
        RECT 29.080 67.890 29.420 68.810 ;
        RECT 29.040 58.390 29.420 67.590 ;
        RECT 29.740 58.390 30.120 75.330 ;
        RECT 30.440 63.070 30.820 75.330 ;
        RECT 30.480 61.770 30.820 62.690 ;
        RECT 30.440 58.390 30.820 61.470 ;
        RECT 31.140 58.390 31.520 75.330 ;
        RECT 31.840 63.070 32.220 75.330 ;
        RECT 31.880 61.770 32.220 62.690 ;
        RECT 31.840 58.390 32.220 61.470 ;
        RECT 32.540 58.390 32.920 75.330 ;
        RECT 33.240 63.070 33.620 75.330 ;
        RECT 33.280 61.770 33.620 62.690 ;
        RECT 33.240 58.390 33.620 61.470 ;
        RECT 33.940 58.390 34.320 75.330 ;
        RECT 34.640 63.070 35.020 75.330 ;
        RECT 34.680 61.770 35.020 62.690 ;
        RECT 34.640 58.390 35.020 61.470 ;
        RECT 35.340 58.390 35.720 75.330 ;
        RECT 36.040 63.070 36.420 75.330 ;
        RECT 36.080 61.770 36.420 62.690 ;
        RECT 36.040 58.390 36.420 61.470 ;
        RECT 36.740 58.390 37.120 75.330 ;
        RECT 37.440 63.070 37.820 75.330 ;
        RECT 37.480 61.770 37.820 62.690 ;
        RECT 37.440 58.390 37.820 61.470 ;
        RECT 38.140 58.390 38.520 75.330 ;
        RECT 38.840 63.070 39.220 75.330 ;
        RECT 38.880 61.770 39.220 62.690 ;
        RECT 38.840 58.390 39.220 61.470 ;
        RECT 39.540 58.390 39.920 75.330 ;
        RECT 40.240 63.070 40.620 75.330 ;
        RECT 40.280 61.770 40.620 62.690 ;
        RECT 40.240 58.390 40.620 61.470 ;
        RECT 40.940 58.390 41.320 75.330 ;
        RECT 41.640 69.190 42.020 75.330 ;
        RECT 41.680 67.890 42.020 68.810 ;
        RECT 41.640 58.390 42.020 67.590 ;
        RECT 42.340 58.390 42.720 75.330 ;
        RECT 43.040 69.190 43.420 75.330 ;
        RECT 43.080 67.890 43.420 68.810 ;
        RECT 43.040 58.390 43.420 67.590 ;
        RECT 43.740 58.390 44.120 75.330 ;
        RECT 44.440 72.250 44.820 75.330 ;
        RECT 44.480 70.950 44.820 71.870 ;
        RECT 44.440 58.390 44.820 70.650 ;
        RECT 45.140 58.390 45.520 75.330 ;
        RECT 45.840 66.130 46.220 75.330 ;
        RECT 45.880 64.830 46.220 65.750 ;
        RECT 45.840 58.390 46.220 64.530 ;
        RECT 46.540 58.390 46.920 75.330 ;
        RECT 47.240 60.010 47.620 75.330 ;
        RECT 47.280 58.710 47.620 59.630 ;
        RECT 47.940 58.390 48.320 75.330 ;
        RECT 48.640 72.250 49.020 75.330 ;
        RECT 48.680 70.950 49.020 71.870 ;
        RECT 48.640 58.390 49.020 70.650 ;
        RECT 49.340 58.390 49.720 75.330 ;
        RECT 50.040 69.190 50.420 75.330 ;
        RECT 50.080 67.890 50.420 68.810 ;
        RECT 50.040 58.390 50.420 67.590 ;
        RECT 50.740 58.390 51.120 75.330 ;
        RECT 51.440 69.190 51.820 75.330 ;
        RECT 51.480 67.890 51.820 68.810 ;
        RECT 51.440 58.390 51.820 67.590 ;
        RECT 52.140 58.390 52.520 75.330 ;
        RECT 52.840 63.070 53.220 75.330 ;
        RECT 52.880 61.770 53.220 62.690 ;
        RECT 52.840 58.390 53.220 61.470 ;
        RECT 53.540 58.390 53.920 75.330 ;
        RECT 54.240 63.070 54.620 75.330 ;
        RECT 54.280 61.770 54.620 62.690 ;
        RECT 54.240 58.390 54.620 61.470 ;
        RECT 54.940 58.390 55.320 75.330 ;
        RECT 55.640 63.070 56.020 75.330 ;
        RECT 55.680 61.770 56.020 62.690 ;
        RECT 55.640 58.390 56.020 61.470 ;
        RECT 56.340 58.390 56.720 75.330 ;
        RECT 57.040 63.070 57.420 75.330 ;
        RECT 57.080 61.770 57.420 62.690 ;
        RECT 57.040 58.390 57.420 61.470 ;
        RECT 57.740 59.360 58.120 75.330 ;
        RECT 58.840 74.320 59.760 74.660 ;
        RECT 58.840 71.260 59.760 71.600 ;
        RECT 58.840 68.200 59.760 68.540 ;
        RECT 58.840 65.140 59.760 65.480 ;
        RECT 58.840 62.080 59.760 62.420 ;
        RECT 59.420 59.360 59.760 59.670 ;
        RECT 57.740 59.020 59.760 59.360 ;
        RECT 57.740 58.390 58.120 59.020 ;
        RECT 59.420 58.750 59.760 59.020 ;
        RECT 12.240 58.310 58.120 58.390 ;
        RECT 8.640 58.010 58.120 58.310 ;
        RECT 12.240 57.930 58.120 58.010 ;
        RECT 8.640 40.910 9.560 41.830 ;
        RECT 12.240 40.990 12.620 57.930 ;
        RECT 12.940 40.990 13.320 57.930 ;
        RECT 13.640 45.670 14.020 57.930 ;
        RECT 13.680 44.370 14.020 45.290 ;
        RECT 13.640 40.990 14.020 44.070 ;
        RECT 14.340 40.990 14.720 57.930 ;
        RECT 15.040 45.670 15.420 57.930 ;
        RECT 15.080 44.370 15.420 45.290 ;
        RECT 15.040 40.990 15.420 44.070 ;
        RECT 15.740 40.990 16.120 57.930 ;
        RECT 16.440 45.670 16.820 57.930 ;
        RECT 16.480 44.370 16.820 45.290 ;
        RECT 16.440 40.990 16.820 44.070 ;
        RECT 17.140 40.990 17.520 57.930 ;
        RECT 17.840 45.670 18.220 57.930 ;
        RECT 17.880 44.370 18.220 45.290 ;
        RECT 17.840 40.990 18.220 44.070 ;
        RECT 18.540 40.990 18.920 57.930 ;
        RECT 19.240 51.790 19.620 57.930 ;
        RECT 19.280 50.490 19.620 51.410 ;
        RECT 19.240 40.990 19.620 50.190 ;
        RECT 19.940 40.990 20.320 57.930 ;
        RECT 20.640 51.790 21.020 57.930 ;
        RECT 20.680 50.490 21.020 51.410 ;
        RECT 20.640 40.990 21.020 50.190 ;
        RECT 21.340 40.990 21.720 57.930 ;
        RECT 22.040 54.850 22.420 57.930 ;
        RECT 22.080 53.550 22.420 54.470 ;
        RECT 22.040 40.990 22.420 53.250 ;
        RECT 22.740 40.990 23.120 57.930 ;
        RECT 23.480 56.610 23.820 57.530 ;
        RECT 23.440 40.990 23.820 56.310 ;
        RECT 24.140 40.990 24.520 57.930 ;
        RECT 24.840 48.730 25.220 57.930 ;
        RECT 24.880 47.430 25.220 48.350 ;
        RECT 24.840 40.990 25.220 47.130 ;
        RECT 25.540 40.990 25.920 57.930 ;
        RECT 26.240 54.850 26.620 57.930 ;
        RECT 26.280 53.550 26.620 54.470 ;
        RECT 26.240 40.990 26.620 53.250 ;
        RECT 26.940 40.990 27.320 57.930 ;
        RECT 27.640 51.790 28.020 57.930 ;
        RECT 27.680 50.490 28.020 51.410 ;
        RECT 27.640 40.990 28.020 50.190 ;
        RECT 28.340 40.990 28.720 57.930 ;
        RECT 29.040 51.790 29.420 57.930 ;
        RECT 29.080 50.490 29.420 51.410 ;
        RECT 29.040 40.990 29.420 50.190 ;
        RECT 29.740 40.990 30.120 57.930 ;
        RECT 30.440 45.670 30.820 57.930 ;
        RECT 30.480 44.370 30.820 45.290 ;
        RECT 30.440 40.990 30.820 44.070 ;
        RECT 31.140 40.990 31.520 57.930 ;
        RECT 31.840 45.670 32.220 57.930 ;
        RECT 31.880 44.370 32.220 45.290 ;
        RECT 31.840 40.990 32.220 44.070 ;
        RECT 32.540 40.990 32.920 57.930 ;
        RECT 33.240 45.670 33.620 57.930 ;
        RECT 33.280 44.370 33.620 45.290 ;
        RECT 33.240 40.990 33.620 44.070 ;
        RECT 33.940 40.990 34.320 57.930 ;
        RECT 34.640 45.670 35.020 57.930 ;
        RECT 34.680 44.370 35.020 45.290 ;
        RECT 34.640 40.990 35.020 44.070 ;
        RECT 35.340 40.990 35.720 57.930 ;
        RECT 36.040 45.670 36.420 57.930 ;
        RECT 36.080 44.370 36.420 45.290 ;
        RECT 36.040 40.990 36.420 44.070 ;
        RECT 36.740 40.990 37.120 57.930 ;
        RECT 37.440 45.670 37.820 57.930 ;
        RECT 37.480 44.370 37.820 45.290 ;
        RECT 37.440 40.990 37.820 44.070 ;
        RECT 38.140 40.990 38.520 57.930 ;
        RECT 38.840 45.670 39.220 57.930 ;
        RECT 38.880 44.370 39.220 45.290 ;
        RECT 38.840 40.990 39.220 44.070 ;
        RECT 39.540 40.990 39.920 57.930 ;
        RECT 40.240 45.670 40.620 57.930 ;
        RECT 40.280 44.370 40.620 45.290 ;
        RECT 40.240 40.990 40.620 44.070 ;
        RECT 40.940 40.990 41.320 57.930 ;
        RECT 41.640 51.790 42.020 57.930 ;
        RECT 41.680 50.490 42.020 51.410 ;
        RECT 41.640 40.990 42.020 50.190 ;
        RECT 42.340 40.990 42.720 57.930 ;
        RECT 43.040 51.790 43.420 57.930 ;
        RECT 43.080 50.490 43.420 51.410 ;
        RECT 43.040 40.990 43.420 50.190 ;
        RECT 43.740 40.990 44.120 57.930 ;
        RECT 44.440 54.850 44.820 57.930 ;
        RECT 44.480 53.550 44.820 54.470 ;
        RECT 44.440 40.990 44.820 53.250 ;
        RECT 45.140 40.990 45.520 57.930 ;
        RECT 45.840 48.730 46.220 57.930 ;
        RECT 45.880 47.430 46.220 48.350 ;
        RECT 45.840 40.990 46.220 47.130 ;
        RECT 46.540 40.990 46.920 57.930 ;
        RECT 47.240 42.610 47.620 57.930 ;
        RECT 47.280 41.310 47.620 42.230 ;
        RECT 47.940 40.990 48.320 57.930 ;
        RECT 48.640 54.850 49.020 57.930 ;
        RECT 48.680 53.550 49.020 54.470 ;
        RECT 48.640 40.990 49.020 53.250 ;
        RECT 49.340 40.990 49.720 57.930 ;
        RECT 50.040 51.790 50.420 57.930 ;
        RECT 50.080 50.490 50.420 51.410 ;
        RECT 50.040 40.990 50.420 50.190 ;
        RECT 50.740 40.990 51.120 57.930 ;
        RECT 51.440 51.790 51.820 57.930 ;
        RECT 51.480 50.490 51.820 51.410 ;
        RECT 51.440 40.990 51.820 50.190 ;
        RECT 52.140 40.990 52.520 57.930 ;
        RECT 52.840 45.670 53.220 57.930 ;
        RECT 52.880 44.370 53.220 45.290 ;
        RECT 52.840 40.990 53.220 44.070 ;
        RECT 53.540 40.990 53.920 57.930 ;
        RECT 54.240 45.670 54.620 57.930 ;
        RECT 54.280 44.370 54.620 45.290 ;
        RECT 54.240 40.990 54.620 44.070 ;
        RECT 54.940 40.990 55.320 57.930 ;
        RECT 55.640 45.670 56.020 57.930 ;
        RECT 55.680 44.370 56.020 45.290 ;
        RECT 55.640 40.990 56.020 44.070 ;
        RECT 56.340 40.990 56.720 57.930 ;
        RECT 57.040 45.670 57.420 57.930 ;
        RECT 57.080 44.370 57.420 45.290 ;
        RECT 57.040 40.990 57.420 44.070 ;
        RECT 57.740 40.990 58.120 57.930 ;
        RECT 61.560 57.530 61.860 110.210 ;
        RECT 62.460 62.690 62.760 110.210 ;
        RECT 63.360 80.090 63.660 110.210 ;
        RECT 64.260 92.330 64.560 110.210 ;
        RECT 64.260 91.410 64.600 92.330 ;
        RECT 64.260 89.270 64.560 91.410 ;
        RECT 64.260 88.350 64.600 89.270 ;
        RECT 64.260 83.150 64.560 88.350 ;
        RECT 65.160 86.210 65.460 110.210 ;
        RECT 65.160 85.290 65.500 86.210 ;
        RECT 64.260 82.230 64.600 83.150 ;
        RECT 63.360 79.170 63.700 80.090 ;
        RECT 64.260 77.030 64.560 82.230 ;
        RECT 64.260 76.110 64.600 77.030 ;
        RECT 66.060 68.810 66.360 110.210 ;
        RECT 66.960 71.870 67.260 110.210 ;
        RECT 66.960 70.950 67.300 71.870 ;
        RECT 66.060 67.890 66.400 68.810 ;
        RECT 67.860 65.750 68.160 110.210 ;
        RECT 68.760 74.930 69.060 110.210 ;
        RECT 72.060 74.930 72.360 110.210 ;
        RECT 68.760 74.010 69.100 74.930 ;
        RECT 72.020 74.010 72.360 74.930 ;
        RECT 72.960 65.750 73.260 110.210 ;
        RECT 73.860 71.870 74.160 110.210 ;
        RECT 73.820 70.950 74.160 71.870 ;
        RECT 74.760 68.810 75.060 110.210 ;
        RECT 75.660 86.210 75.960 110.210 ;
        RECT 76.560 92.330 76.860 110.210 ;
        RECT 76.520 91.410 76.860 92.330 ;
        RECT 76.560 89.270 76.860 91.410 ;
        RECT 76.520 88.350 76.860 89.270 ;
        RECT 75.620 85.290 75.960 86.210 ;
        RECT 76.560 83.150 76.860 88.350 ;
        RECT 76.520 82.230 76.860 83.150 ;
        RECT 76.560 77.030 76.860 82.230 ;
        RECT 77.460 80.090 77.760 110.210 ;
        RECT 77.420 79.170 77.760 80.090 ;
        RECT 76.520 76.110 76.860 77.030 ;
        RECT 74.720 67.890 75.060 68.810 ;
        RECT 67.860 64.830 68.200 65.750 ;
        RECT 72.920 64.830 73.260 65.750 ;
        RECT 78.360 62.690 78.660 110.210 ;
        RECT 62.460 61.770 62.800 62.690 ;
        RECT 78.320 61.770 78.660 62.690 ;
        RECT 79.260 57.530 79.560 110.210 ;
        RECT 80.160 109.730 80.460 110.210 ;
        RECT 80.120 108.810 80.460 109.730 ;
        RECT 83.000 110.130 128.880 110.510 ;
        RECT 81.360 109.120 82.280 109.460 ;
        RECT 80.160 106.670 80.460 108.810 ;
        RECT 80.120 105.750 80.460 106.670 ;
        RECT 81.360 106.060 82.280 106.400 ;
        RECT 80.160 103.610 80.460 105.750 ;
        RECT 80.120 102.690 80.460 103.610 ;
        RECT 81.360 103.000 82.280 103.340 ;
        RECT 80.160 100.550 80.460 102.690 ;
        RECT 80.120 99.630 80.460 100.550 ;
        RECT 81.360 99.940 82.280 100.280 ;
        RECT 80.160 97.490 80.460 99.630 ;
        RECT 80.120 96.570 80.460 97.490 ;
        RECT 81.360 96.880 82.280 97.220 ;
        RECT 80.160 94.430 80.460 96.570 ;
        RECT 80.120 93.510 80.460 94.430 ;
        RECT 81.360 93.820 82.280 94.160 ;
        RECT 83.000 93.190 83.380 110.130 ;
        RECT 83.700 97.870 84.080 110.130 ;
        RECT 83.700 96.570 84.040 97.490 ;
        RECT 83.700 93.190 84.080 96.270 ;
        RECT 84.400 93.190 84.780 110.130 ;
        RECT 85.100 97.870 85.480 110.130 ;
        RECT 85.100 96.570 85.440 97.490 ;
        RECT 85.100 93.190 85.480 96.270 ;
        RECT 85.800 93.190 86.180 110.130 ;
        RECT 86.500 97.870 86.880 110.130 ;
        RECT 86.500 96.570 86.840 97.490 ;
        RECT 86.500 93.190 86.880 96.270 ;
        RECT 87.200 93.190 87.580 110.130 ;
        RECT 87.900 97.870 88.280 110.130 ;
        RECT 87.900 96.570 88.240 97.490 ;
        RECT 87.900 93.190 88.280 96.270 ;
        RECT 88.600 93.190 88.980 110.130 ;
        RECT 89.300 103.990 89.680 110.130 ;
        RECT 89.300 102.690 89.640 103.610 ;
        RECT 89.300 93.190 89.680 102.390 ;
        RECT 90.000 93.190 90.380 110.130 ;
        RECT 90.700 103.990 91.080 110.130 ;
        RECT 90.700 102.690 91.040 103.610 ;
        RECT 90.700 93.190 91.080 102.390 ;
        RECT 91.400 93.190 91.780 110.130 ;
        RECT 92.100 107.050 92.480 110.130 ;
        RECT 92.100 105.750 92.440 106.670 ;
        RECT 92.100 93.190 92.480 105.450 ;
        RECT 92.800 93.190 93.180 110.130 ;
        RECT 93.500 94.810 93.880 110.130 ;
        RECT 93.500 93.510 93.840 94.430 ;
        RECT 94.200 93.190 94.580 110.130 ;
        RECT 94.900 100.930 95.280 110.130 ;
        RECT 94.900 99.630 95.240 100.550 ;
        RECT 94.900 93.190 95.280 99.330 ;
        RECT 95.600 93.190 95.980 110.130 ;
        RECT 96.300 107.050 96.680 110.130 ;
        RECT 96.300 105.750 96.640 106.670 ;
        RECT 96.300 93.190 96.680 105.450 ;
        RECT 97.000 93.190 97.380 110.130 ;
        RECT 97.700 103.990 98.080 110.130 ;
        RECT 97.700 102.690 98.040 103.610 ;
        RECT 97.700 93.190 98.080 102.390 ;
        RECT 98.400 93.190 98.780 110.130 ;
        RECT 99.100 103.990 99.480 110.130 ;
        RECT 99.100 102.690 99.440 103.610 ;
        RECT 99.100 93.190 99.480 102.390 ;
        RECT 99.800 93.190 100.180 110.130 ;
        RECT 100.500 97.870 100.880 110.130 ;
        RECT 100.500 96.570 100.840 97.490 ;
        RECT 100.500 93.190 100.880 96.270 ;
        RECT 101.200 93.190 101.580 110.130 ;
        RECT 101.900 97.870 102.280 110.130 ;
        RECT 101.900 96.570 102.240 97.490 ;
        RECT 101.900 93.190 102.280 96.270 ;
        RECT 102.600 93.190 102.980 110.130 ;
        RECT 103.300 97.870 103.680 110.130 ;
        RECT 103.300 96.570 103.640 97.490 ;
        RECT 103.300 93.190 103.680 96.270 ;
        RECT 104.000 93.190 104.380 110.130 ;
        RECT 104.700 97.870 105.080 110.130 ;
        RECT 104.700 96.570 105.040 97.490 ;
        RECT 104.700 93.190 105.080 96.270 ;
        RECT 105.400 93.190 105.780 110.130 ;
        RECT 106.100 97.870 106.480 110.130 ;
        RECT 106.100 96.570 106.440 97.490 ;
        RECT 106.100 93.190 106.480 96.270 ;
        RECT 106.800 93.190 107.180 110.130 ;
        RECT 107.500 97.870 107.880 110.130 ;
        RECT 107.500 96.570 107.840 97.490 ;
        RECT 107.500 93.190 107.880 96.270 ;
        RECT 108.200 93.190 108.580 110.130 ;
        RECT 108.900 97.870 109.280 110.130 ;
        RECT 108.900 96.570 109.240 97.490 ;
        RECT 108.900 93.190 109.280 96.270 ;
        RECT 109.600 93.190 109.980 110.130 ;
        RECT 110.300 97.870 110.680 110.130 ;
        RECT 110.300 96.570 110.640 97.490 ;
        RECT 110.300 93.190 110.680 96.270 ;
        RECT 111.000 93.190 111.380 110.130 ;
        RECT 111.700 103.990 112.080 110.130 ;
        RECT 111.700 102.690 112.040 103.610 ;
        RECT 111.700 93.190 112.080 102.390 ;
        RECT 112.400 93.190 112.780 110.130 ;
        RECT 113.100 103.990 113.480 110.130 ;
        RECT 113.100 102.690 113.440 103.610 ;
        RECT 113.100 93.190 113.480 102.390 ;
        RECT 113.800 93.190 114.180 110.130 ;
        RECT 114.500 107.050 114.880 110.130 ;
        RECT 114.500 105.750 114.840 106.670 ;
        RECT 114.500 93.190 114.880 105.450 ;
        RECT 115.200 93.190 115.580 110.130 ;
        RECT 115.900 100.930 116.280 110.130 ;
        RECT 115.900 99.630 116.240 100.550 ;
        RECT 115.900 93.190 116.280 99.330 ;
        RECT 116.600 93.190 116.980 110.130 ;
        RECT 117.300 108.810 117.640 109.730 ;
        RECT 117.300 93.190 117.680 108.510 ;
        RECT 118.000 93.190 118.380 110.130 ;
        RECT 118.700 107.050 119.080 110.130 ;
        RECT 118.700 105.750 119.040 106.670 ;
        RECT 118.700 93.190 119.080 105.450 ;
        RECT 119.400 93.190 119.780 110.130 ;
        RECT 120.100 103.990 120.480 110.130 ;
        RECT 120.100 102.690 120.440 103.610 ;
        RECT 120.100 93.190 120.480 102.390 ;
        RECT 120.800 93.190 121.180 110.130 ;
        RECT 121.500 103.990 121.880 110.130 ;
        RECT 121.500 102.690 121.840 103.610 ;
        RECT 121.500 93.190 121.880 102.390 ;
        RECT 122.200 93.190 122.580 110.130 ;
        RECT 122.900 97.870 123.280 110.130 ;
        RECT 122.900 96.570 123.240 97.490 ;
        RECT 122.900 93.190 123.280 96.270 ;
        RECT 123.600 93.190 123.980 110.130 ;
        RECT 124.300 97.870 124.680 110.130 ;
        RECT 124.300 96.570 124.640 97.490 ;
        RECT 124.300 93.190 124.680 96.270 ;
        RECT 125.000 93.190 125.380 110.130 ;
        RECT 125.700 97.870 126.080 110.130 ;
        RECT 125.700 96.570 126.040 97.490 ;
        RECT 125.700 93.190 126.080 96.270 ;
        RECT 126.400 93.190 126.780 110.130 ;
        RECT 127.100 97.870 127.480 110.130 ;
        RECT 127.100 96.570 127.440 97.490 ;
        RECT 127.100 93.190 127.480 96.270 ;
        RECT 127.800 93.190 128.180 110.130 ;
        RECT 128.500 93.190 128.880 110.130 ;
        RECT 140.920 100.490 141.220 116.030 ;
        RECT 143.680 115.590 144.600 115.930 ;
        RECT 143.680 115.010 144.600 115.050 ;
        RECT 145.060 115.010 145.360 119.990 ;
        RECT 149.020 118.090 149.320 121.750 ;
        RECT 149.800 118.090 150.720 118.130 ;
        RECT 149.020 117.790 150.720 118.090 ;
        RECT 147.640 117.350 148.560 117.690 ;
        RECT 147.640 116.470 148.560 116.810 ;
        RECT 143.680 114.710 145.360 115.010 ;
        RECT 149.800 114.570 150.720 114.610 ;
        RECT 149.800 114.270 151.480 114.570 ;
        RECT 149.800 112.810 150.720 112.850 ;
        RECT 149.020 112.510 150.720 112.810 ;
        RECT 143.680 112.070 144.600 112.410 ;
        RECT 147.640 112.070 148.560 112.410 ;
        RECT 147.640 111.490 148.560 111.530 ;
        RECT 149.020 111.490 149.320 112.510 ;
        RECT 147.640 111.190 149.320 111.490 ;
        RECT 141.520 111.050 142.440 111.090 ;
        RECT 141.520 110.750 143.200 111.050 ;
        RECT 142.900 109.730 143.200 110.750 ;
        RECT 143.680 110.310 144.600 110.650 ;
        RECT 147.640 110.310 148.560 110.650 ;
        RECT 143.680 109.730 144.600 109.770 ;
        RECT 142.900 109.430 144.600 109.730 ;
        RECT 149.020 107.530 149.320 111.190 ;
        RECT 149.800 109.290 150.720 109.330 ;
        RECT 151.180 109.290 151.480 114.270 ;
        RECT 149.800 108.990 151.480 109.290 ;
        RECT 149.800 107.530 150.720 107.570 ;
        RECT 149.020 107.230 150.720 107.530 ;
        RECT 143.680 106.790 144.600 107.130 ;
        RECT 147.640 106.790 148.560 107.130 ;
        RECT 141.520 105.770 142.440 105.810 ;
        RECT 141.520 105.470 142.600 105.770 ;
        RECT 142.300 105.170 143.200 105.470 ;
        RECT 142.900 100.930 143.200 105.170 ;
        RECT 143.680 103.270 144.600 103.610 ;
        RECT 147.640 103.270 148.560 103.610 ;
        RECT 143.680 101.510 144.600 101.850 ;
        RECT 147.640 101.510 148.560 101.850 ;
        RECT 143.680 100.930 144.600 100.970 ;
        RECT 142.900 100.630 144.600 100.930 ;
        RECT 147.640 100.630 148.560 100.970 ;
        RECT 141.520 100.490 142.440 100.530 ;
        RECT 140.920 100.190 142.440 100.490 ;
        RECT 147.640 99.170 148.560 99.210 ;
        RECT 151.180 99.170 151.480 108.990 ;
        RECT 147.640 98.870 151.480 99.170 ;
        RECT 143.680 97.990 144.600 98.330 ;
        RECT 147.640 97.990 148.560 98.330 ;
        RECT 147.640 97.410 148.560 97.450 ;
        RECT 147.640 97.110 149.320 97.410 ;
        RECT 143.680 96.230 144.600 96.570 ;
        RECT 147.640 96.230 148.560 96.570 ;
        RECT 143.680 95.650 144.600 95.690 ;
        RECT 143.680 95.350 145.360 95.650 ;
        RECT 141.520 94.910 142.440 95.250 ;
        RECT 83.000 93.110 128.880 93.190 ;
        RECT 131.580 93.110 131.920 93.730 ;
        RECT 83.000 92.810 131.920 93.110 ;
        RECT 83.000 92.730 128.880 92.810 ;
        RECT 81.360 91.720 82.280 92.060 ;
        RECT 81.360 88.660 82.280 89.000 ;
        RECT 81.360 85.600 82.280 85.940 ;
        RECT 81.360 82.540 82.280 82.880 ;
        RECT 81.360 79.480 82.280 79.820 ;
        RECT 81.360 76.420 82.280 76.760 ;
        RECT 83.000 75.790 83.380 92.730 ;
        RECT 83.700 80.470 84.080 92.730 ;
        RECT 83.700 79.170 84.040 80.090 ;
        RECT 83.700 75.790 84.080 78.870 ;
        RECT 84.400 75.790 84.780 92.730 ;
        RECT 85.100 80.470 85.480 92.730 ;
        RECT 85.100 79.170 85.440 80.090 ;
        RECT 85.100 75.790 85.480 78.870 ;
        RECT 85.800 75.790 86.180 92.730 ;
        RECT 86.500 80.470 86.880 92.730 ;
        RECT 86.500 79.170 86.840 80.090 ;
        RECT 86.500 75.790 86.880 78.870 ;
        RECT 87.200 75.790 87.580 92.730 ;
        RECT 87.900 80.470 88.280 92.730 ;
        RECT 87.900 79.170 88.240 80.090 ;
        RECT 87.900 75.790 88.280 78.870 ;
        RECT 88.600 75.790 88.980 92.730 ;
        RECT 89.300 86.590 89.680 92.730 ;
        RECT 89.300 85.290 89.640 86.210 ;
        RECT 89.300 75.790 89.680 84.990 ;
        RECT 90.000 75.790 90.380 92.730 ;
        RECT 90.700 86.590 91.080 92.730 ;
        RECT 90.700 85.290 91.040 86.210 ;
        RECT 90.700 75.790 91.080 84.990 ;
        RECT 91.400 75.790 91.780 92.730 ;
        RECT 92.100 89.650 92.480 92.730 ;
        RECT 92.100 88.350 92.440 89.270 ;
        RECT 92.100 75.790 92.480 88.050 ;
        RECT 92.800 75.790 93.180 92.730 ;
        RECT 93.500 77.410 93.880 92.730 ;
        RECT 93.500 76.110 93.840 77.030 ;
        RECT 94.200 75.790 94.580 92.730 ;
        RECT 94.900 83.530 95.280 92.730 ;
        RECT 94.900 82.230 95.240 83.150 ;
        RECT 94.900 75.790 95.280 81.930 ;
        RECT 95.600 75.790 95.980 92.730 ;
        RECT 96.300 89.650 96.680 92.730 ;
        RECT 96.300 88.350 96.640 89.270 ;
        RECT 96.300 75.790 96.680 88.050 ;
        RECT 97.000 75.790 97.380 92.730 ;
        RECT 97.700 86.590 98.080 92.730 ;
        RECT 97.700 85.290 98.040 86.210 ;
        RECT 97.700 75.790 98.080 84.990 ;
        RECT 98.400 75.790 98.780 92.730 ;
        RECT 99.100 86.590 99.480 92.730 ;
        RECT 99.100 85.290 99.440 86.210 ;
        RECT 99.100 75.790 99.480 84.990 ;
        RECT 99.800 75.790 100.180 92.730 ;
        RECT 100.500 80.470 100.880 92.730 ;
        RECT 100.500 79.170 100.840 80.090 ;
        RECT 100.500 75.790 100.880 78.870 ;
        RECT 101.200 75.790 101.580 92.730 ;
        RECT 101.900 80.470 102.280 92.730 ;
        RECT 101.900 79.170 102.240 80.090 ;
        RECT 101.900 75.790 102.280 78.870 ;
        RECT 102.600 75.790 102.980 92.730 ;
        RECT 103.300 80.470 103.680 92.730 ;
        RECT 103.300 79.170 103.640 80.090 ;
        RECT 103.300 75.790 103.680 78.870 ;
        RECT 104.000 75.790 104.380 92.730 ;
        RECT 104.700 80.470 105.080 92.730 ;
        RECT 104.700 79.170 105.040 80.090 ;
        RECT 104.700 75.790 105.080 78.870 ;
        RECT 105.400 75.790 105.780 92.730 ;
        RECT 106.100 80.470 106.480 92.730 ;
        RECT 106.100 79.170 106.440 80.090 ;
        RECT 106.100 75.790 106.480 78.870 ;
        RECT 106.800 75.790 107.180 92.730 ;
        RECT 107.500 80.470 107.880 92.730 ;
        RECT 107.500 79.170 107.840 80.090 ;
        RECT 107.500 75.790 107.880 78.870 ;
        RECT 108.200 75.790 108.580 92.730 ;
        RECT 108.900 80.470 109.280 92.730 ;
        RECT 108.900 79.170 109.240 80.090 ;
        RECT 108.900 75.790 109.280 78.870 ;
        RECT 109.600 75.790 109.980 92.730 ;
        RECT 110.300 80.470 110.680 92.730 ;
        RECT 110.300 79.170 110.640 80.090 ;
        RECT 110.300 75.790 110.680 78.870 ;
        RECT 111.000 75.790 111.380 92.730 ;
        RECT 111.700 86.590 112.080 92.730 ;
        RECT 111.700 85.290 112.040 86.210 ;
        RECT 111.700 75.790 112.080 84.990 ;
        RECT 112.400 75.790 112.780 92.730 ;
        RECT 113.100 86.590 113.480 92.730 ;
        RECT 113.100 85.290 113.440 86.210 ;
        RECT 113.100 75.790 113.480 84.990 ;
        RECT 113.800 75.790 114.180 92.730 ;
        RECT 114.500 89.650 114.880 92.730 ;
        RECT 114.500 88.350 114.840 89.270 ;
        RECT 114.500 75.790 114.880 88.050 ;
        RECT 115.200 75.790 115.580 92.730 ;
        RECT 115.900 83.530 116.280 92.730 ;
        RECT 115.900 82.230 116.240 83.150 ;
        RECT 115.900 75.790 116.280 81.930 ;
        RECT 116.600 75.790 116.980 92.730 ;
        RECT 117.300 91.410 117.640 92.330 ;
        RECT 117.300 75.790 117.680 91.110 ;
        RECT 118.000 75.790 118.380 92.730 ;
        RECT 118.700 89.650 119.080 92.730 ;
        RECT 118.700 88.350 119.040 89.270 ;
        RECT 118.700 75.790 119.080 88.050 ;
        RECT 119.400 75.790 119.780 92.730 ;
        RECT 120.100 86.590 120.480 92.730 ;
        RECT 120.100 85.290 120.440 86.210 ;
        RECT 120.100 75.790 120.480 84.990 ;
        RECT 120.800 75.790 121.180 92.730 ;
        RECT 121.500 86.590 121.880 92.730 ;
        RECT 121.500 85.290 121.840 86.210 ;
        RECT 121.500 75.790 121.880 84.990 ;
        RECT 122.200 75.790 122.580 92.730 ;
        RECT 122.900 80.470 123.280 92.730 ;
        RECT 122.900 79.170 123.240 80.090 ;
        RECT 122.900 75.790 123.280 78.870 ;
        RECT 123.600 75.790 123.980 92.730 ;
        RECT 124.300 80.470 124.680 92.730 ;
        RECT 124.300 79.170 124.640 80.090 ;
        RECT 124.300 75.790 124.680 78.870 ;
        RECT 125.000 75.790 125.380 92.730 ;
        RECT 125.700 80.470 126.080 92.730 ;
        RECT 125.700 79.170 126.040 80.090 ;
        RECT 125.700 75.790 126.080 78.870 ;
        RECT 126.400 75.790 126.780 92.730 ;
        RECT 127.100 80.470 127.480 92.730 ;
        RECT 127.100 79.170 127.440 80.090 ;
        RECT 127.100 75.790 127.480 78.870 ;
        RECT 127.800 75.790 128.180 92.730 ;
        RECT 128.500 75.790 128.880 92.730 ;
        RECT 141.520 91.690 142.440 91.730 ;
        RECT 140.920 91.390 142.440 91.690 ;
        RECT 83.000 75.710 128.880 75.790 ;
        RECT 131.580 75.710 131.920 76.330 ;
        RECT 83.000 75.410 131.920 75.710 ;
        RECT 140.920 75.850 141.220 91.390 ;
        RECT 143.680 90.950 144.600 91.290 ;
        RECT 143.680 90.370 144.600 90.410 ;
        RECT 145.060 90.370 145.360 95.350 ;
        RECT 149.020 93.450 149.320 97.110 ;
        RECT 149.800 93.450 150.720 93.490 ;
        RECT 149.020 93.150 150.720 93.450 ;
        RECT 147.640 92.710 148.560 93.050 ;
        RECT 147.640 91.830 148.560 92.170 ;
        RECT 143.680 90.070 145.360 90.370 ;
        RECT 149.800 89.930 150.720 89.970 ;
        RECT 149.800 89.630 151.480 89.930 ;
        RECT 149.800 88.170 150.720 88.210 ;
        RECT 149.020 87.870 150.720 88.170 ;
        RECT 143.680 87.430 144.600 87.770 ;
        RECT 147.640 87.430 148.560 87.770 ;
        RECT 147.640 86.850 148.560 86.890 ;
        RECT 149.020 86.850 149.320 87.870 ;
        RECT 147.640 86.550 149.320 86.850 ;
        RECT 141.520 86.410 142.440 86.450 ;
        RECT 141.520 86.110 143.200 86.410 ;
        RECT 142.900 85.090 143.200 86.110 ;
        RECT 143.680 85.670 144.600 86.010 ;
        RECT 147.640 85.670 148.560 86.010 ;
        RECT 143.680 85.090 144.600 85.130 ;
        RECT 142.900 84.790 144.600 85.090 ;
        RECT 149.020 82.890 149.320 86.550 ;
        RECT 149.800 84.650 150.720 84.690 ;
        RECT 151.180 84.650 151.480 89.630 ;
        RECT 149.800 84.350 151.480 84.650 ;
        RECT 149.800 82.890 150.720 82.930 ;
        RECT 149.020 82.590 150.720 82.890 ;
        RECT 143.680 82.150 144.600 82.490 ;
        RECT 147.640 82.150 148.560 82.490 ;
        RECT 141.520 81.130 142.440 81.170 ;
        RECT 141.520 80.830 142.600 81.130 ;
        RECT 142.300 80.530 143.200 80.830 ;
        RECT 142.900 76.290 143.200 80.530 ;
        RECT 143.680 78.630 144.600 78.970 ;
        RECT 147.640 78.630 148.560 78.970 ;
        RECT 143.680 76.870 144.600 77.210 ;
        RECT 147.640 76.870 148.560 77.210 ;
        RECT 143.680 76.290 144.600 76.330 ;
        RECT 142.900 75.990 144.600 76.290 ;
        RECT 147.640 75.990 148.560 76.330 ;
        RECT 141.520 75.850 142.440 75.890 ;
        RECT 140.920 75.550 142.440 75.850 ;
        RECT 83.000 75.330 128.880 75.410 ;
        RECT 81.360 74.320 82.280 74.660 ;
        RECT 81.360 71.260 82.280 71.600 ;
        RECT 81.360 68.200 82.280 68.540 ;
        RECT 81.360 65.140 82.280 65.480 ;
        RECT 81.360 62.080 82.280 62.420 ;
        RECT 81.360 59.360 81.700 59.670 ;
        RECT 83.000 59.360 83.380 75.330 ;
        RECT 83.700 63.070 84.080 75.330 ;
        RECT 83.700 61.770 84.040 62.690 ;
        RECT 81.360 59.020 83.380 59.360 ;
        RECT 81.360 58.750 81.700 59.020 ;
        RECT 58.840 56.920 59.760 57.260 ;
        RECT 61.560 56.610 61.900 57.530 ;
        RECT 79.220 56.610 79.560 57.530 ;
        RECT 83.000 58.390 83.380 59.020 ;
        RECT 83.700 58.390 84.080 61.470 ;
        RECT 84.400 58.390 84.780 75.330 ;
        RECT 85.100 63.070 85.480 75.330 ;
        RECT 85.100 61.770 85.440 62.690 ;
        RECT 85.100 58.390 85.480 61.470 ;
        RECT 85.800 58.390 86.180 75.330 ;
        RECT 86.500 63.070 86.880 75.330 ;
        RECT 86.500 61.770 86.840 62.690 ;
        RECT 86.500 58.390 86.880 61.470 ;
        RECT 87.200 58.390 87.580 75.330 ;
        RECT 87.900 63.070 88.280 75.330 ;
        RECT 87.900 61.770 88.240 62.690 ;
        RECT 87.900 58.390 88.280 61.470 ;
        RECT 88.600 58.390 88.980 75.330 ;
        RECT 89.300 69.190 89.680 75.330 ;
        RECT 89.300 67.890 89.640 68.810 ;
        RECT 89.300 58.390 89.680 67.590 ;
        RECT 90.000 58.390 90.380 75.330 ;
        RECT 90.700 69.190 91.080 75.330 ;
        RECT 90.700 67.890 91.040 68.810 ;
        RECT 90.700 58.390 91.080 67.590 ;
        RECT 91.400 58.390 91.780 75.330 ;
        RECT 92.100 72.250 92.480 75.330 ;
        RECT 92.100 70.950 92.440 71.870 ;
        RECT 92.100 58.390 92.480 70.650 ;
        RECT 92.800 58.390 93.180 75.330 ;
        RECT 93.500 60.010 93.880 75.330 ;
        RECT 93.500 58.710 93.840 59.630 ;
        RECT 94.200 58.390 94.580 75.330 ;
        RECT 94.900 66.130 95.280 75.330 ;
        RECT 94.900 64.830 95.240 65.750 ;
        RECT 94.900 58.390 95.280 64.530 ;
        RECT 95.600 58.390 95.980 75.330 ;
        RECT 96.300 72.250 96.680 75.330 ;
        RECT 96.300 70.950 96.640 71.870 ;
        RECT 96.300 58.390 96.680 70.650 ;
        RECT 97.000 58.390 97.380 75.330 ;
        RECT 97.700 69.190 98.080 75.330 ;
        RECT 97.700 67.890 98.040 68.810 ;
        RECT 97.700 58.390 98.080 67.590 ;
        RECT 98.400 58.390 98.780 75.330 ;
        RECT 99.100 69.190 99.480 75.330 ;
        RECT 99.100 67.890 99.440 68.810 ;
        RECT 99.100 58.390 99.480 67.590 ;
        RECT 99.800 58.390 100.180 75.330 ;
        RECT 100.500 63.070 100.880 75.330 ;
        RECT 100.500 61.770 100.840 62.690 ;
        RECT 100.500 58.390 100.880 61.470 ;
        RECT 101.200 58.390 101.580 75.330 ;
        RECT 101.900 63.070 102.280 75.330 ;
        RECT 101.900 61.770 102.240 62.690 ;
        RECT 101.900 58.390 102.280 61.470 ;
        RECT 102.600 58.390 102.980 75.330 ;
        RECT 103.300 63.070 103.680 75.330 ;
        RECT 103.300 61.770 103.640 62.690 ;
        RECT 103.300 58.390 103.680 61.470 ;
        RECT 104.000 58.390 104.380 75.330 ;
        RECT 104.700 63.070 105.080 75.330 ;
        RECT 104.700 61.770 105.040 62.690 ;
        RECT 104.700 58.390 105.080 61.470 ;
        RECT 105.400 58.390 105.780 75.330 ;
        RECT 106.100 63.070 106.480 75.330 ;
        RECT 106.100 61.770 106.440 62.690 ;
        RECT 106.100 58.390 106.480 61.470 ;
        RECT 106.800 58.390 107.180 75.330 ;
        RECT 107.500 63.070 107.880 75.330 ;
        RECT 107.500 61.770 107.840 62.690 ;
        RECT 107.500 58.390 107.880 61.470 ;
        RECT 108.200 58.390 108.580 75.330 ;
        RECT 108.900 63.070 109.280 75.330 ;
        RECT 108.900 61.770 109.240 62.690 ;
        RECT 108.900 58.390 109.280 61.470 ;
        RECT 109.600 58.390 109.980 75.330 ;
        RECT 110.300 63.070 110.680 75.330 ;
        RECT 110.300 61.770 110.640 62.690 ;
        RECT 110.300 58.390 110.680 61.470 ;
        RECT 111.000 58.390 111.380 75.330 ;
        RECT 111.700 69.190 112.080 75.330 ;
        RECT 111.700 67.890 112.040 68.810 ;
        RECT 111.700 58.390 112.080 67.590 ;
        RECT 112.400 58.390 112.780 75.330 ;
        RECT 113.100 69.190 113.480 75.330 ;
        RECT 113.100 67.890 113.440 68.810 ;
        RECT 113.100 58.390 113.480 67.590 ;
        RECT 113.800 58.390 114.180 75.330 ;
        RECT 114.500 72.250 114.880 75.330 ;
        RECT 114.500 70.950 114.840 71.870 ;
        RECT 114.500 58.390 114.880 70.650 ;
        RECT 115.200 58.390 115.580 75.330 ;
        RECT 115.900 66.130 116.280 75.330 ;
        RECT 115.900 64.830 116.240 65.750 ;
        RECT 115.900 58.390 116.280 64.530 ;
        RECT 116.600 58.390 116.980 75.330 ;
        RECT 117.300 74.010 117.640 74.930 ;
        RECT 117.300 58.390 117.680 73.710 ;
        RECT 118.000 58.390 118.380 75.330 ;
        RECT 118.700 72.250 119.080 75.330 ;
        RECT 118.700 70.950 119.040 71.870 ;
        RECT 118.700 58.390 119.080 70.650 ;
        RECT 119.400 58.390 119.780 75.330 ;
        RECT 120.100 69.190 120.480 75.330 ;
        RECT 120.100 67.890 120.440 68.810 ;
        RECT 120.100 58.390 120.480 67.590 ;
        RECT 120.800 58.390 121.180 75.330 ;
        RECT 121.500 69.190 121.880 75.330 ;
        RECT 121.500 67.890 121.840 68.810 ;
        RECT 121.500 58.390 121.880 67.590 ;
        RECT 122.200 58.390 122.580 75.330 ;
        RECT 122.900 63.070 123.280 75.330 ;
        RECT 122.900 61.770 123.240 62.690 ;
        RECT 122.900 58.390 123.280 61.470 ;
        RECT 123.600 58.390 123.980 75.330 ;
        RECT 124.300 63.070 124.680 75.330 ;
        RECT 124.300 61.770 124.640 62.690 ;
        RECT 124.300 58.390 124.680 61.470 ;
        RECT 125.000 58.390 125.380 75.330 ;
        RECT 125.700 63.070 126.080 75.330 ;
        RECT 125.700 61.770 126.040 62.690 ;
        RECT 125.700 58.390 126.080 61.470 ;
        RECT 126.400 58.390 126.780 75.330 ;
        RECT 127.100 63.070 127.480 75.330 ;
        RECT 127.100 61.770 127.440 62.690 ;
        RECT 127.100 58.390 127.480 61.470 ;
        RECT 127.800 58.390 128.180 75.330 ;
        RECT 128.500 58.390 128.880 75.330 ;
        RECT 147.640 74.530 148.560 74.570 ;
        RECT 151.180 74.530 151.480 84.350 ;
        RECT 147.640 74.230 151.480 74.530 ;
        RECT 143.680 73.350 144.600 73.690 ;
        RECT 147.640 73.350 148.560 73.690 ;
        RECT 147.640 72.770 148.560 72.810 ;
        RECT 147.640 72.470 149.320 72.770 ;
        RECT 143.680 71.590 144.600 71.930 ;
        RECT 147.640 71.590 148.560 71.930 ;
        RECT 143.680 71.010 144.600 71.050 ;
        RECT 143.680 70.710 145.360 71.010 ;
        RECT 141.520 70.270 142.440 70.610 ;
        RECT 141.520 67.050 142.440 67.090 ;
        RECT 140.920 66.750 142.440 67.050 ;
        RECT 83.000 58.310 128.880 58.390 ;
        RECT 131.580 58.310 131.920 58.930 ;
        RECT 83.000 58.010 131.920 58.310 ;
        RECT 83.000 57.930 128.880 58.010 ;
        RECT 81.360 56.920 82.280 57.260 ;
        RECT 61.560 54.470 61.860 56.610 ;
        RECT 79.260 54.470 79.560 56.610 ;
        RECT 58.840 53.860 59.760 54.200 ;
        RECT 61.560 53.550 61.900 54.470 ;
        RECT 79.220 53.550 79.560 54.470 ;
        RECT 81.360 53.860 82.280 54.200 ;
        RECT 61.560 51.410 61.860 53.550 ;
        RECT 79.260 51.410 79.560 53.550 ;
        RECT 58.840 50.800 59.760 51.140 ;
        RECT 61.560 50.490 61.900 51.410 ;
        RECT 79.220 50.490 79.560 51.410 ;
        RECT 81.360 50.800 82.280 51.140 ;
        RECT 61.560 48.350 61.860 50.490 ;
        RECT 79.260 48.350 79.560 50.490 ;
        RECT 58.840 47.740 59.760 48.080 ;
        RECT 61.560 47.430 61.900 48.350 ;
        RECT 79.220 47.430 79.560 48.350 ;
        RECT 81.360 47.740 82.280 48.080 ;
        RECT 61.560 45.290 61.860 47.430 ;
        RECT 79.260 45.290 79.560 47.430 ;
        RECT 58.840 44.680 59.760 45.020 ;
        RECT 61.560 44.370 61.900 45.290 ;
        RECT 79.220 44.370 79.560 45.290 ;
        RECT 81.360 44.680 82.280 45.020 ;
        RECT 61.560 42.230 61.860 44.370 ;
        RECT 79.260 42.230 79.560 44.370 ;
        RECT 58.840 41.620 59.760 41.960 ;
        RECT 61.560 41.310 61.900 42.230 ;
        RECT 79.220 41.310 79.560 42.230 ;
        RECT 81.360 41.620 82.280 41.960 ;
        RECT 12.240 40.910 58.120 40.990 ;
        RECT 8.640 40.610 58.120 40.910 ;
        RECT 83.000 40.990 83.380 57.930 ;
        RECT 83.700 45.670 84.080 57.930 ;
        RECT 83.700 44.370 84.040 45.290 ;
        RECT 83.700 40.990 84.080 44.070 ;
        RECT 84.400 40.990 84.780 57.930 ;
        RECT 85.100 45.670 85.480 57.930 ;
        RECT 85.100 44.370 85.440 45.290 ;
        RECT 85.100 40.990 85.480 44.070 ;
        RECT 85.800 40.990 86.180 57.930 ;
        RECT 86.500 45.670 86.880 57.930 ;
        RECT 86.500 44.370 86.840 45.290 ;
        RECT 86.500 40.990 86.880 44.070 ;
        RECT 87.200 40.990 87.580 57.930 ;
        RECT 87.900 45.670 88.280 57.930 ;
        RECT 87.900 44.370 88.240 45.290 ;
        RECT 87.900 40.990 88.280 44.070 ;
        RECT 88.600 40.990 88.980 57.930 ;
        RECT 89.300 51.790 89.680 57.930 ;
        RECT 89.300 50.490 89.640 51.410 ;
        RECT 89.300 40.990 89.680 50.190 ;
        RECT 90.000 40.990 90.380 57.930 ;
        RECT 90.700 51.790 91.080 57.930 ;
        RECT 90.700 50.490 91.040 51.410 ;
        RECT 90.700 40.990 91.080 50.190 ;
        RECT 91.400 40.990 91.780 57.930 ;
        RECT 92.100 54.850 92.480 57.930 ;
        RECT 92.100 53.550 92.440 54.470 ;
        RECT 92.100 40.990 92.480 53.250 ;
        RECT 92.800 40.990 93.180 57.930 ;
        RECT 93.500 42.610 93.880 57.930 ;
        RECT 93.500 41.310 93.840 42.230 ;
        RECT 94.200 40.990 94.580 57.930 ;
        RECT 94.900 48.730 95.280 57.930 ;
        RECT 94.900 47.430 95.240 48.350 ;
        RECT 94.900 40.990 95.280 47.130 ;
        RECT 95.600 40.990 95.980 57.930 ;
        RECT 96.300 54.850 96.680 57.930 ;
        RECT 96.300 53.550 96.640 54.470 ;
        RECT 96.300 40.990 96.680 53.250 ;
        RECT 97.000 40.990 97.380 57.930 ;
        RECT 97.700 51.790 98.080 57.930 ;
        RECT 97.700 50.490 98.040 51.410 ;
        RECT 97.700 40.990 98.080 50.190 ;
        RECT 98.400 40.990 98.780 57.930 ;
        RECT 99.100 51.790 99.480 57.930 ;
        RECT 99.100 50.490 99.440 51.410 ;
        RECT 99.100 40.990 99.480 50.190 ;
        RECT 99.800 40.990 100.180 57.930 ;
        RECT 100.500 45.670 100.880 57.930 ;
        RECT 100.500 44.370 100.840 45.290 ;
        RECT 100.500 40.990 100.880 44.070 ;
        RECT 101.200 40.990 101.580 57.930 ;
        RECT 101.900 45.670 102.280 57.930 ;
        RECT 101.900 44.370 102.240 45.290 ;
        RECT 101.900 40.990 102.280 44.070 ;
        RECT 102.600 40.990 102.980 57.930 ;
        RECT 103.300 45.670 103.680 57.930 ;
        RECT 103.300 44.370 103.640 45.290 ;
        RECT 103.300 40.990 103.680 44.070 ;
        RECT 104.000 40.990 104.380 57.930 ;
        RECT 104.700 45.670 105.080 57.930 ;
        RECT 104.700 44.370 105.040 45.290 ;
        RECT 104.700 40.990 105.080 44.070 ;
        RECT 105.400 40.990 105.780 57.930 ;
        RECT 106.100 45.670 106.480 57.930 ;
        RECT 106.100 44.370 106.440 45.290 ;
        RECT 106.100 40.990 106.480 44.070 ;
        RECT 106.800 40.990 107.180 57.930 ;
        RECT 107.500 45.670 107.880 57.930 ;
        RECT 107.500 44.370 107.840 45.290 ;
        RECT 107.500 40.990 107.880 44.070 ;
        RECT 108.200 40.990 108.580 57.930 ;
        RECT 108.900 45.670 109.280 57.930 ;
        RECT 108.900 44.370 109.240 45.290 ;
        RECT 108.900 40.990 109.280 44.070 ;
        RECT 109.600 40.990 109.980 57.930 ;
        RECT 110.300 45.670 110.680 57.930 ;
        RECT 110.300 44.370 110.640 45.290 ;
        RECT 110.300 40.990 110.680 44.070 ;
        RECT 111.000 40.990 111.380 57.930 ;
        RECT 111.700 51.790 112.080 57.930 ;
        RECT 111.700 50.490 112.040 51.410 ;
        RECT 111.700 40.990 112.080 50.190 ;
        RECT 112.400 40.990 112.780 57.930 ;
        RECT 113.100 51.790 113.480 57.930 ;
        RECT 113.100 50.490 113.440 51.410 ;
        RECT 113.100 40.990 113.480 50.190 ;
        RECT 113.800 40.990 114.180 57.930 ;
        RECT 114.500 54.850 114.880 57.930 ;
        RECT 114.500 53.550 114.840 54.470 ;
        RECT 114.500 40.990 114.880 53.250 ;
        RECT 115.200 40.990 115.580 57.930 ;
        RECT 115.900 48.730 116.280 57.930 ;
        RECT 115.900 47.430 116.240 48.350 ;
        RECT 115.900 40.990 116.280 47.130 ;
        RECT 116.600 40.990 116.980 57.930 ;
        RECT 117.300 56.610 117.640 57.530 ;
        RECT 117.300 40.990 117.680 56.310 ;
        RECT 118.000 40.990 118.380 57.930 ;
        RECT 118.700 54.850 119.080 57.930 ;
        RECT 118.700 53.550 119.040 54.470 ;
        RECT 118.700 40.990 119.080 53.250 ;
        RECT 119.400 40.990 119.780 57.930 ;
        RECT 120.100 51.790 120.480 57.930 ;
        RECT 120.100 50.490 120.440 51.410 ;
        RECT 120.100 40.990 120.480 50.190 ;
        RECT 120.800 40.990 121.180 57.930 ;
        RECT 121.500 51.790 121.880 57.930 ;
        RECT 121.500 50.490 121.840 51.410 ;
        RECT 121.500 40.990 121.880 50.190 ;
        RECT 122.200 40.990 122.580 57.930 ;
        RECT 122.900 45.670 123.280 57.930 ;
        RECT 122.900 44.370 123.240 45.290 ;
        RECT 122.900 40.990 123.280 44.070 ;
        RECT 123.600 40.990 123.980 57.930 ;
        RECT 124.300 45.670 124.680 57.930 ;
        RECT 124.300 44.370 124.640 45.290 ;
        RECT 124.300 40.990 124.680 44.070 ;
        RECT 125.000 40.990 125.380 57.930 ;
        RECT 125.700 45.670 126.080 57.930 ;
        RECT 125.700 44.370 126.040 45.290 ;
        RECT 125.700 40.990 126.080 44.070 ;
        RECT 126.400 40.990 126.780 57.930 ;
        RECT 127.100 45.670 127.480 57.930 ;
        RECT 127.100 44.370 127.440 45.290 ;
        RECT 127.100 40.990 127.480 44.070 ;
        RECT 127.800 40.990 128.180 57.930 ;
        RECT 128.500 40.990 128.880 57.930 ;
        RECT 140.920 51.210 141.220 66.750 ;
        RECT 143.680 66.310 144.600 66.650 ;
        RECT 143.680 65.730 144.600 65.770 ;
        RECT 145.060 65.730 145.360 70.710 ;
        RECT 149.020 68.810 149.320 72.470 ;
        RECT 149.800 68.810 150.720 68.850 ;
        RECT 149.020 68.510 150.720 68.810 ;
        RECT 147.640 68.070 148.560 68.410 ;
        RECT 147.640 67.190 148.560 67.530 ;
        RECT 143.680 65.430 145.360 65.730 ;
        RECT 149.800 65.290 150.720 65.330 ;
        RECT 149.800 64.990 151.480 65.290 ;
        RECT 149.800 63.530 150.720 63.570 ;
        RECT 149.020 63.230 150.720 63.530 ;
        RECT 143.680 62.790 144.600 63.130 ;
        RECT 147.640 62.790 148.560 63.130 ;
        RECT 147.640 62.210 148.560 62.250 ;
        RECT 149.020 62.210 149.320 63.230 ;
        RECT 147.640 61.910 149.320 62.210 ;
        RECT 141.520 61.770 142.440 61.810 ;
        RECT 141.520 61.470 143.200 61.770 ;
        RECT 142.900 60.450 143.200 61.470 ;
        RECT 143.680 61.030 144.600 61.370 ;
        RECT 147.640 61.030 148.560 61.370 ;
        RECT 143.680 60.450 144.600 60.490 ;
        RECT 142.900 60.150 144.600 60.450 ;
        RECT 149.020 58.250 149.320 61.910 ;
        RECT 149.800 60.010 150.720 60.050 ;
        RECT 151.180 60.010 151.480 64.990 ;
        RECT 149.800 59.710 151.480 60.010 ;
        RECT 149.800 58.250 150.720 58.290 ;
        RECT 149.020 57.950 150.720 58.250 ;
        RECT 143.680 57.510 144.600 57.850 ;
        RECT 147.640 57.510 148.560 57.850 ;
        RECT 141.520 56.490 142.440 56.530 ;
        RECT 141.520 56.190 142.600 56.490 ;
        RECT 142.300 55.890 143.200 56.190 ;
        RECT 142.900 51.650 143.200 55.890 ;
        RECT 143.680 53.990 144.600 54.330 ;
        RECT 147.640 53.990 148.560 54.330 ;
        RECT 143.680 52.230 144.600 52.570 ;
        RECT 147.640 52.230 148.560 52.570 ;
        RECT 143.680 51.650 144.600 51.690 ;
        RECT 142.900 51.350 144.600 51.650 ;
        RECT 147.640 51.350 148.560 51.690 ;
        RECT 141.520 51.210 142.440 51.250 ;
        RECT 140.920 50.910 142.440 51.210 ;
        RECT 147.640 49.890 148.560 49.930 ;
        RECT 151.180 49.890 151.480 59.710 ;
        RECT 147.640 49.590 151.480 49.890 ;
        RECT 143.680 48.710 144.600 49.050 ;
        RECT 147.640 48.710 148.560 49.050 ;
        RECT 147.640 48.130 148.560 48.170 ;
        RECT 147.640 47.830 149.320 48.130 ;
        RECT 143.680 46.950 144.600 47.290 ;
        RECT 147.640 46.950 148.560 47.290 ;
        RECT 143.680 46.370 144.600 46.410 ;
        RECT 143.680 46.070 145.360 46.370 ;
        RECT 141.520 45.630 142.440 45.970 ;
        RECT 141.520 42.410 142.440 42.450 ;
        RECT 140.920 42.110 142.440 42.410 ;
        RECT 83.000 40.910 128.880 40.990 ;
        RECT 131.580 40.910 131.920 41.530 ;
        RECT 83.000 40.610 131.920 40.910 ;
        RECT 13.600 38.540 49.240 38.980 ;
        RECT 13.600 37.660 48.520 38.100 ;
        RECT 13.600 36.340 13.960 37.660 ;
        RECT 48.880 37.220 49.240 38.540 ;
        RECT 14.320 36.780 49.240 37.220 ;
        RECT 13.600 35.900 48.520 36.340 ;
        RECT 13.600 34.580 13.960 35.900 ;
        RECT 48.880 35.460 49.240 36.780 ;
        RECT 14.320 35.020 49.240 35.460 ;
        RECT 92.080 38.540 127.720 38.980 ;
        RECT 92.080 37.220 92.440 38.540 ;
        RECT 92.800 37.660 127.720 38.100 ;
        RECT 92.080 36.780 127.000 37.220 ;
        RECT 92.080 35.460 92.440 36.780 ;
        RECT 127.360 36.340 127.720 37.660 ;
        RECT 92.800 35.900 127.720 36.340 ;
        RECT 92.080 35.020 127.000 35.460 ;
        RECT 127.360 34.580 127.720 35.900 ;
        RECT 13.600 34.140 49.240 34.580 ;
        RECT 92.080 34.140 127.720 34.580 ;
        RECT 13.600 33.260 49.240 33.700 ;
        RECT 13.600 32.380 48.520 32.820 ;
        RECT 13.600 31.060 13.960 32.380 ;
        RECT 48.880 31.940 49.240 33.260 ;
        RECT 92.080 33.260 127.720 33.700 ;
        RECT 54.800 32.010 55.720 32.350 ;
        RECT 58.760 32.010 59.680 32.350 ;
        RECT 81.640 32.010 82.560 32.350 ;
        RECT 85.600 32.010 86.520 32.350 ;
        RECT 14.320 31.500 49.240 31.940 ;
        RECT 13.600 30.620 48.520 31.060 ;
        RECT 13.600 29.300 13.960 30.620 ;
        RECT 48.880 30.180 49.240 31.500 ;
        RECT 92.080 31.940 92.440 33.260 ;
        RECT 92.800 32.380 127.720 32.820 ;
        RECT 92.080 31.500 127.000 31.940 ;
        RECT 54.800 31.130 55.720 31.470 ;
        RECT 58.760 31.130 59.680 31.470 ;
        RECT 81.640 31.130 82.560 31.470 ;
        RECT 85.600 31.130 86.520 31.470 ;
        RECT 58.760 30.550 59.680 30.590 ;
        RECT 81.640 30.550 82.560 30.590 ;
        RECT 58.760 30.250 67.660 30.550 ;
        RECT 61.680 30.210 62.600 30.250 ;
        RECT 14.320 29.740 49.240 30.180 ;
        RECT 54.800 29.370 55.720 29.710 ;
        RECT 58.760 29.370 59.680 29.710 ;
        RECT 13.600 28.860 49.240 29.300 ;
        RECT 54.800 28.490 55.720 28.830 ;
        RECT 58.760 28.490 59.680 28.830 ;
        RECT 13.600 27.980 49.240 28.420 ;
        RECT 13.600 27.100 48.520 27.540 ;
        RECT 13.600 25.780 13.960 27.100 ;
        RECT 48.880 26.660 49.240 27.980 ;
        RECT 54.800 27.610 55.720 27.950 ;
        RECT 58.760 27.610 59.680 27.950 ;
        RECT 54.800 27.180 55.720 27.240 ;
        RECT 54.800 26.900 60.460 27.180 ;
        RECT 55.180 26.880 60.460 26.900 ;
        RECT 14.320 26.220 49.240 26.660 ;
        RECT 13.600 25.340 48.520 25.780 ;
        RECT 13.600 24.020 13.960 25.340 ;
        RECT 48.880 24.900 49.240 26.220 ;
        RECT 54.800 25.850 55.720 26.190 ;
        RECT 58.760 25.850 59.680 26.190 ;
        RECT 54.800 24.970 55.720 25.310 ;
        RECT 58.680 24.970 59.600 25.310 ;
        RECT 14.320 24.460 49.240 24.900 ;
        RECT 60.160 24.830 60.460 26.880 ;
        RECT 67.360 26.590 67.660 30.250 ;
        RECT 73.660 30.250 82.560 30.550 ;
        RECT 68.120 26.590 69.040 26.630 ;
        RECT 67.360 26.290 69.040 26.590 ;
        RECT 72.280 26.590 73.200 26.630 ;
        RECT 73.660 26.590 73.960 30.250 ;
        RECT 78.720 30.210 79.640 30.250 ;
        RECT 92.080 30.180 92.440 31.500 ;
        RECT 127.360 31.060 127.720 32.380 ;
        RECT 92.800 30.620 127.720 31.060 ;
        RECT 92.080 29.740 127.000 30.180 ;
        RECT 81.640 29.370 82.560 29.710 ;
        RECT 85.600 29.370 86.520 29.710 ;
        RECT 127.360 29.300 127.720 30.620 ;
        RECT 92.080 28.860 127.720 29.300 ;
        RECT 81.640 28.490 82.560 28.830 ;
        RECT 85.600 28.490 86.520 28.830 ;
        RECT 92.080 27.980 127.720 28.420 ;
        RECT 81.640 27.610 82.560 27.950 ;
        RECT 85.600 27.610 86.520 27.950 ;
        RECT 85.600 27.180 86.520 27.240 ;
        RECT 72.280 26.290 73.960 26.590 ;
        RECT 80.860 26.900 86.520 27.180 ;
        RECT 80.860 26.880 86.140 26.900 ;
        RECT 65.800 25.850 66.720 26.190 ;
        RECT 74.440 25.850 75.360 26.190 ;
        RECT 60.920 24.830 61.840 24.870 ;
        RECT 60.160 24.530 61.840 24.830 ;
        RECT 79.480 24.830 80.400 24.870 ;
        RECT 80.860 24.830 81.160 26.880 ;
        RECT 92.080 26.660 92.440 27.980 ;
        RECT 92.800 27.100 127.720 27.540 ;
        RECT 92.080 26.220 127.000 26.660 ;
        RECT 81.640 25.850 82.560 26.190 ;
        RECT 85.600 25.850 86.520 26.190 ;
        RECT 81.720 24.970 82.640 25.310 ;
        RECT 85.600 24.970 86.520 25.310 ;
        RECT 79.480 24.530 81.160 24.830 ;
        RECT 92.080 24.900 92.440 26.220 ;
        RECT 127.360 25.780 127.720 27.100 ;
        RECT 140.920 26.570 141.220 42.110 ;
        RECT 143.680 41.670 144.600 42.010 ;
        RECT 143.680 41.090 144.600 41.130 ;
        RECT 145.060 41.090 145.360 46.070 ;
        RECT 149.020 44.170 149.320 47.830 ;
        RECT 149.800 44.170 150.720 44.210 ;
        RECT 149.020 43.870 150.720 44.170 ;
        RECT 147.640 43.430 148.560 43.770 ;
        RECT 147.640 42.550 148.560 42.890 ;
        RECT 143.680 40.790 145.360 41.090 ;
        RECT 149.800 40.650 150.720 40.690 ;
        RECT 149.800 40.350 151.480 40.650 ;
        RECT 149.800 38.890 150.720 38.930 ;
        RECT 149.020 38.590 150.720 38.890 ;
        RECT 143.680 38.150 144.600 38.490 ;
        RECT 147.640 38.150 148.560 38.490 ;
        RECT 147.640 37.570 148.560 37.610 ;
        RECT 149.020 37.570 149.320 38.590 ;
        RECT 147.640 37.270 149.320 37.570 ;
        RECT 141.520 37.130 142.440 37.170 ;
        RECT 141.520 36.830 143.200 37.130 ;
        RECT 142.900 35.810 143.200 36.830 ;
        RECT 143.680 36.390 144.600 36.730 ;
        RECT 147.640 36.390 148.560 36.730 ;
        RECT 143.680 35.810 144.600 35.850 ;
        RECT 142.900 35.510 144.600 35.810 ;
        RECT 149.020 33.610 149.320 37.270 ;
        RECT 149.800 35.370 150.720 35.410 ;
        RECT 151.180 35.370 151.480 40.350 ;
        RECT 149.800 35.070 151.480 35.370 ;
        RECT 149.800 33.610 150.720 33.650 ;
        RECT 149.020 33.310 150.720 33.610 ;
        RECT 143.680 32.870 144.600 33.210 ;
        RECT 147.640 32.870 148.560 33.210 ;
        RECT 141.520 31.850 142.440 31.890 ;
        RECT 141.520 31.550 142.600 31.850 ;
        RECT 142.300 31.250 143.200 31.550 ;
        RECT 142.900 27.010 143.200 31.250 ;
        RECT 143.680 29.350 144.600 29.690 ;
        RECT 147.640 29.350 148.560 29.690 ;
        RECT 143.680 27.590 144.600 27.930 ;
        RECT 147.640 27.590 148.560 27.930 ;
        RECT 143.680 27.010 144.600 27.050 ;
        RECT 142.900 26.710 144.600 27.010 ;
        RECT 147.640 26.710 148.560 27.050 ;
        RECT 141.520 26.570 142.440 26.610 ;
        RECT 140.920 26.270 142.440 26.570 ;
        RECT 92.800 25.340 127.720 25.780 ;
        RECT 92.080 24.460 127.000 24.900 ;
        RECT 127.360 24.020 127.720 25.340 ;
        RECT 147.640 25.250 148.560 25.290 ;
        RECT 151.180 25.250 151.480 35.070 ;
        RECT 147.640 24.950 151.480 25.250 ;
        RECT 143.680 24.070 144.600 24.410 ;
        RECT 147.640 24.070 148.560 24.410 ;
        RECT 13.600 23.580 49.240 24.020 ;
        RECT 92.080 23.580 127.720 24.020 ;
        RECT 52.640 23.510 53.560 23.550 ;
        RECT 54.800 23.510 55.720 23.550 ;
        RECT 52.640 23.210 55.720 23.510 ;
        RECT 85.600 23.510 86.520 23.550 ;
        RECT 87.760 23.510 88.680 23.550 ;
        RECT 85.600 23.210 88.680 23.510 ;
        RECT 13.600 22.700 49.240 23.140 ;
        RECT 60.920 22.770 61.840 23.110 ;
        RECT 79.480 22.770 80.400 23.110 ;
        RECT 13.600 21.820 48.520 22.260 ;
        RECT 13.600 20.500 13.960 21.820 ;
        RECT 48.880 21.380 49.240 22.700 ;
        RECT 92.080 22.700 127.720 23.140 ;
        RECT 58.760 22.330 59.680 22.670 ;
        RECT 81.640 22.330 82.560 22.670 ;
        RECT 58.760 21.750 59.680 21.790 ;
        RECT 81.640 21.750 82.560 21.790 ;
        RECT 58.760 21.450 65.500 21.750 ;
        RECT 14.320 20.940 49.240 21.380 ;
        RECT 13.600 20.060 48.520 20.500 ;
        RECT 13.600 18.740 13.960 20.060 ;
        RECT 48.880 19.620 49.240 20.940 ;
        RECT 54.800 20.570 55.720 20.910 ;
        RECT 14.320 19.180 49.240 19.620 ;
        RECT 52.640 19.250 53.560 19.590 ;
        RECT 54.800 18.810 55.720 19.150 ;
        RECT 58.760 18.810 59.680 19.150 ;
        RECT 13.600 18.300 49.240 18.740 ;
        RECT 54.800 17.930 55.720 18.270 ;
        RECT 58.760 17.930 59.680 18.270 ;
        RECT 65.200 18.230 65.500 21.450 ;
        RECT 75.820 21.450 82.560 21.750 ;
        RECT 65.800 18.810 66.720 19.150 ;
        RECT 74.440 18.810 75.360 19.150 ;
        RECT 65.960 18.230 66.880 18.270 ;
        RECT 65.200 17.930 66.880 18.230 ;
        RECT 74.440 18.230 75.360 18.270 ;
        RECT 75.820 18.230 76.120 21.450 ;
        RECT 92.080 21.380 92.440 22.700 ;
        RECT 143.680 22.310 144.600 22.650 ;
        RECT 147.640 22.310 148.560 22.650 ;
        RECT 92.800 21.820 127.720 22.260 ;
        RECT 92.080 20.940 127.000 21.380 ;
        RECT 85.600 20.570 86.520 20.910 ;
        RECT 92.080 19.620 92.440 20.940 ;
        RECT 127.360 20.500 127.720 21.820 ;
        RECT 147.640 21.430 148.560 21.770 ;
        RECT 92.800 20.060 127.720 20.500 ;
        RECT 87.760 19.250 88.680 19.590 ;
        RECT 92.080 19.180 127.000 19.620 ;
        RECT 81.640 18.810 82.560 19.150 ;
        RECT 85.600 18.810 86.520 19.150 ;
        RECT 127.360 18.740 127.720 20.060 ;
        RECT 143.680 18.790 144.600 19.130 ;
        RECT 147.640 18.790 148.560 19.130 ;
        RECT 92.080 18.300 127.720 18.740 ;
        RECT 74.440 17.930 76.120 18.230 ;
        RECT 81.640 17.930 82.560 18.270 ;
        RECT 85.600 17.930 86.520 18.270 ;
        RECT 13.600 17.420 49.240 17.860 ;
        RECT 52.640 17.790 53.560 17.830 ;
        RECT 52.640 17.490 54.340 17.790 ;
        RECT 68.040 17.490 68.960 17.830 ;
        RECT 72.360 17.490 73.280 17.830 ;
        RECT 87.760 17.790 88.680 17.830 ;
        RECT 86.980 17.490 88.680 17.790 ;
        RECT 13.600 16.540 48.520 16.980 ;
        RECT 13.600 15.220 13.960 16.540 ;
        RECT 48.880 16.100 49.240 17.420 ;
        RECT 54.040 16.470 54.340 17.490 ;
        RECT 54.800 16.470 55.720 16.510 ;
        RECT 54.040 16.170 55.720 16.470 ;
        RECT 58.760 16.360 59.680 16.700 ;
        RECT 81.640 16.360 82.560 16.700 ;
        RECT 85.600 16.470 86.520 16.510 ;
        RECT 86.980 16.470 87.280 17.490 ;
        RECT 85.600 16.170 87.280 16.470 ;
        RECT 92.080 17.420 127.720 17.860 ;
        RECT 14.320 15.660 49.240 16.100 ;
        RECT 92.080 16.100 92.440 17.420 ;
        RECT 143.680 17.030 144.600 17.370 ;
        RECT 147.640 17.030 148.560 17.370 ;
        RECT 92.800 16.540 127.720 16.980 ;
        RECT 60.840 15.730 61.760 16.070 ;
        RECT 79.560 15.730 80.480 16.070 ;
        RECT 13.600 14.780 48.520 15.220 ;
        RECT 13.600 13.460 13.960 14.780 ;
        RECT 48.880 14.340 49.240 15.660 ;
        RECT 54.800 15.290 55.720 15.630 ;
        RECT 58.760 15.290 59.680 15.630 ;
        RECT 54.800 14.410 55.720 14.750 ;
        RECT 58.760 14.410 59.680 14.750 ;
        RECT 14.320 13.900 49.240 14.340 ;
        RECT 54.800 13.530 55.720 13.870 ;
        RECT 58.760 13.530 59.680 13.870 ;
        RECT 13.600 13.020 49.240 13.460 ;
        RECT 58.680 9.640 59.600 10.560 ;
        RECT 54.720 6.040 55.640 6.960 ;
        RECT 61.150 5.360 61.450 15.730 ;
        RECT 65.880 14.370 66.800 14.710 ;
        RECT 74.520 14.370 75.440 14.710 ;
        RECT 79.870 5.360 80.170 15.730 ;
        RECT 92.080 15.660 127.000 16.100 ;
        RECT 81.640 15.290 82.560 15.630 ;
        RECT 85.600 15.290 86.520 15.630 ;
        RECT 81.640 14.410 82.560 14.750 ;
        RECT 85.600 14.410 86.520 14.750 ;
        RECT 92.080 14.340 92.440 15.660 ;
        RECT 127.360 15.220 127.720 16.540 ;
        RECT 143.680 15.270 144.600 15.610 ;
        RECT 147.640 15.270 148.560 15.610 ;
        RECT 92.800 14.780 127.720 15.220 ;
        RECT 92.080 13.900 127.000 14.340 ;
        RECT 81.640 13.530 82.560 13.870 ;
        RECT 85.600 13.530 86.520 13.870 ;
        RECT 127.360 13.460 127.720 14.780 ;
        RECT 143.680 14.390 144.600 14.730 ;
        RECT 92.080 13.020 127.720 13.460 ;
        RECT 143.680 11.750 144.600 12.090 ;
        RECT 147.640 11.750 148.560 12.090 ;
        RECT 81.640 9.640 82.560 10.560 ;
        RECT 143.680 9.990 144.600 10.330 ;
        RECT 147.640 9.990 148.560 10.330 ;
        RECT 143.680 9.110 144.600 9.450 ;
        RECT 147.640 9.110 148.560 9.450 ;
        RECT 85.600 6.040 86.520 6.960 ;
        RECT 143.680 6.470 144.600 6.810 ;
        RECT 147.640 6.470 148.560 6.810 ;
        RECT 60.840 5.020 61.760 5.360 ;
        RECT 79.560 5.020 80.480 5.360 ;
        RECT 143.680 4.710 144.600 5.050 ;
        RECT 147.640 4.710 148.560 5.050 ;
        RECT 61.600 4.000 62.520 4.340 ;
        RECT 78.720 4.000 79.640 4.340 ;
        RECT 143.680 3.830 144.600 4.170 ;
        RECT 147.640 3.830 148.560 4.170 ;
        RECT 143.680 2.950 144.600 3.290 ;
        RECT 147.640 2.950 148.560 3.290 ;
      LAYER via ;
        RECT 24.640 221.770 24.920 222.050 ;
        RECT 25.160 221.770 25.440 222.050 ;
        RECT 24.640 221.250 24.920 221.530 ;
        RECT 25.160 221.250 25.440 221.530 ;
        RECT 27.600 221.770 27.880 222.050 ;
        RECT 28.120 221.770 28.400 222.050 ;
        RECT 27.600 221.250 27.880 221.530 ;
        RECT 28.120 221.250 28.400 221.530 ;
        RECT 49.840 221.770 50.120 222.050 ;
        RECT 50.360 221.770 50.640 222.050 ;
        RECT 49.840 221.250 50.120 221.530 ;
        RECT 50.360 221.250 50.640 221.530 ;
        RECT 52.800 221.770 53.080 222.050 ;
        RECT 53.320 221.770 53.600 222.050 ;
        RECT 52.800 221.250 53.080 221.530 ;
        RECT 53.320 221.250 53.600 221.530 ;
        RECT 75.040 221.770 75.320 222.050 ;
        RECT 75.560 221.770 75.840 222.050 ;
        RECT 75.040 221.250 75.320 221.530 ;
        RECT 75.560 221.250 75.840 221.530 ;
        RECT 78.000 221.770 78.280 222.050 ;
        RECT 78.520 221.770 78.800 222.050 ;
        RECT 78.000 221.250 78.280 221.530 ;
        RECT 78.520 221.250 78.800 221.530 ;
        RECT 100.240 221.770 100.520 222.050 ;
        RECT 100.760 221.770 101.040 222.050 ;
        RECT 100.240 221.250 100.520 221.530 ;
        RECT 100.760 221.250 101.040 221.530 ;
        RECT 143.740 222.100 144.020 222.380 ;
        RECT 144.260 222.100 144.540 222.380 ;
        RECT 147.700 222.100 147.980 222.380 ;
        RECT 148.220 222.100 148.500 222.380 ;
        RECT 103.200 221.770 103.480 222.050 ;
        RECT 103.720 221.770 104.000 222.050 ;
        RECT 103.200 221.250 103.480 221.530 ;
        RECT 103.720 221.250 104.000 221.530 ;
        RECT 143.740 221.220 144.020 221.500 ;
        RECT 144.260 221.220 144.540 221.500 ;
        RECT 147.700 221.220 147.980 221.500 ;
        RECT 148.220 221.220 148.500 221.500 ;
        RECT 143.740 219.460 144.020 219.740 ;
        RECT 144.260 219.460 144.540 219.740 ;
        RECT 147.700 219.460 147.980 219.740 ;
        RECT 148.220 219.460 148.500 219.740 ;
        RECT 21.760 218.170 22.040 218.450 ;
        RECT 22.280 218.170 22.560 218.450 ;
        RECT 21.760 217.650 22.040 217.930 ;
        RECT 22.280 217.650 22.560 217.930 ;
        RECT 30.480 218.170 30.760 218.450 ;
        RECT 31.000 218.170 31.280 218.450 ;
        RECT 30.480 217.650 30.760 217.930 ;
        RECT 31.000 217.650 31.280 217.930 ;
        RECT 46.960 218.170 47.240 218.450 ;
        RECT 47.480 218.170 47.760 218.450 ;
        RECT 46.960 217.650 47.240 217.930 ;
        RECT 47.480 217.650 47.760 217.930 ;
        RECT 55.680 218.170 55.960 218.450 ;
        RECT 56.200 218.170 56.480 218.450 ;
        RECT 55.680 217.650 55.960 217.930 ;
        RECT 56.200 217.650 56.480 217.930 ;
        RECT 72.160 218.170 72.440 218.450 ;
        RECT 72.680 218.170 72.960 218.450 ;
        RECT 72.160 217.650 72.440 217.930 ;
        RECT 72.680 217.650 72.960 217.930 ;
        RECT 80.880 218.170 81.160 218.450 ;
        RECT 81.400 218.170 81.680 218.450 ;
        RECT 80.880 217.650 81.160 217.930 ;
        RECT 81.400 217.650 81.680 217.930 ;
        RECT 97.360 218.170 97.640 218.450 ;
        RECT 97.880 218.170 98.160 218.450 ;
        RECT 97.360 217.650 97.640 217.930 ;
        RECT 97.880 217.650 98.160 217.930 ;
        RECT 106.080 218.170 106.360 218.450 ;
        RECT 106.600 218.170 106.880 218.450 ;
        RECT 106.080 217.650 106.360 217.930 ;
        RECT 106.600 217.650 106.880 217.930 ;
        RECT 122.560 218.170 122.840 218.450 ;
        RECT 123.080 218.170 123.360 218.450 ;
        RECT 141.580 218.140 141.860 218.420 ;
        RECT 142.100 218.140 142.380 218.420 ;
        RECT 122.560 217.650 122.840 217.930 ;
        RECT 123.080 217.650 123.360 217.930 ;
        RECT 17.800 214.570 18.080 214.850 ;
        RECT 18.320 214.570 18.600 214.850 ;
        RECT 17.800 214.050 18.080 214.330 ;
        RECT 18.320 214.050 18.600 214.330 ;
        RECT 34.440 214.570 34.720 214.850 ;
        RECT 34.960 214.570 35.240 214.850 ;
        RECT 34.440 214.050 34.720 214.330 ;
        RECT 34.960 214.050 35.240 214.330 ;
        RECT 43.000 214.570 43.280 214.850 ;
        RECT 43.520 214.570 43.800 214.850 ;
        RECT 43.000 214.050 43.280 214.330 ;
        RECT 43.520 214.050 43.800 214.330 ;
        RECT 59.640 214.570 59.920 214.850 ;
        RECT 60.160 214.570 60.440 214.850 ;
        RECT 59.640 214.050 59.920 214.330 ;
        RECT 60.160 214.050 60.440 214.330 ;
        RECT 68.200 214.570 68.480 214.850 ;
        RECT 68.720 214.570 69.000 214.850 ;
        RECT 68.200 214.050 68.480 214.330 ;
        RECT 68.720 214.050 69.000 214.330 ;
        RECT 84.840 214.570 85.120 214.850 ;
        RECT 85.360 214.570 85.640 214.850 ;
        RECT 84.840 214.050 85.120 214.330 ;
        RECT 85.360 214.050 85.640 214.330 ;
        RECT 93.400 214.570 93.680 214.850 ;
        RECT 93.920 214.570 94.200 214.850 ;
        RECT 93.400 214.050 93.680 214.330 ;
        RECT 93.920 214.050 94.200 214.330 ;
        RECT 110.040 214.570 110.320 214.850 ;
        RECT 110.560 214.570 110.840 214.850 ;
        RECT 110.040 214.050 110.320 214.330 ;
        RECT 110.560 214.050 110.840 214.330 ;
        RECT 118.600 214.570 118.880 214.850 ;
        RECT 119.120 214.570 119.400 214.850 ;
        RECT 118.600 214.050 118.880 214.330 ;
        RECT 119.120 214.050 119.400 214.330 ;
        RECT 17.800 210.830 18.080 211.110 ;
        RECT 18.320 210.830 18.600 211.110 ;
        RECT 21.760 210.830 22.040 211.110 ;
        RECT 22.280 210.830 22.560 211.110 ;
        RECT 30.560 210.830 30.840 211.110 ;
        RECT 31.080 210.830 31.360 211.110 ;
        RECT 34.520 210.830 34.800 211.110 ;
        RECT 35.040 210.830 35.320 211.110 ;
        RECT 43.000 210.830 43.280 211.110 ;
        RECT 43.520 210.830 43.800 211.110 ;
        RECT 46.960 210.830 47.240 211.110 ;
        RECT 47.480 210.830 47.760 211.110 ;
        RECT 55.760 210.830 56.040 211.110 ;
        RECT 56.280 210.830 56.560 211.110 ;
        RECT 59.720 210.830 60.000 211.110 ;
        RECT 60.240 210.830 60.520 211.110 ;
        RECT 68.200 210.830 68.480 211.110 ;
        RECT 68.720 210.830 69.000 211.110 ;
        RECT 72.160 210.830 72.440 211.110 ;
        RECT 72.680 210.830 72.960 211.110 ;
        RECT 80.960 210.830 81.240 211.110 ;
        RECT 81.480 210.830 81.760 211.110 ;
        RECT 84.920 210.830 85.200 211.110 ;
        RECT 85.440 210.830 85.720 211.110 ;
        RECT 93.400 210.830 93.680 211.110 ;
        RECT 93.920 210.830 94.200 211.110 ;
        RECT 97.360 210.830 97.640 211.110 ;
        RECT 97.880 210.830 98.160 211.110 ;
        RECT 106.160 210.830 106.440 211.110 ;
        RECT 106.680 210.830 106.960 211.110 ;
        RECT 110.120 210.830 110.400 211.110 ;
        RECT 110.640 210.830 110.920 211.110 ;
        RECT 17.800 209.950 18.080 210.230 ;
        RECT 18.320 209.950 18.600 210.230 ;
        RECT 21.760 209.950 22.040 210.230 ;
        RECT 22.280 209.950 22.560 210.230 ;
        RECT 30.560 209.950 30.840 210.230 ;
        RECT 31.080 209.950 31.360 210.230 ;
        RECT 34.520 209.950 34.800 210.230 ;
        RECT 35.040 209.950 35.320 210.230 ;
        RECT 43.000 209.950 43.280 210.230 ;
        RECT 43.520 209.950 43.800 210.230 ;
        RECT 46.960 209.950 47.240 210.230 ;
        RECT 47.480 209.950 47.760 210.230 ;
        RECT 55.760 209.950 56.040 210.230 ;
        RECT 56.280 209.950 56.560 210.230 ;
        RECT 59.720 209.950 60.000 210.230 ;
        RECT 60.240 209.950 60.520 210.230 ;
        RECT 68.200 209.950 68.480 210.230 ;
        RECT 68.720 209.950 69.000 210.230 ;
        RECT 72.160 209.950 72.440 210.230 ;
        RECT 72.680 209.950 72.960 210.230 ;
        RECT 80.960 209.950 81.240 210.230 ;
        RECT 81.480 209.950 81.760 210.230 ;
        RECT 84.920 209.950 85.200 210.230 ;
        RECT 85.440 209.950 85.720 210.230 ;
        RECT 93.400 209.950 93.680 210.230 ;
        RECT 93.920 209.950 94.200 210.230 ;
        RECT 97.360 209.950 97.640 210.230 ;
        RECT 97.880 209.950 98.160 210.230 ;
        RECT 106.160 209.950 106.440 210.230 ;
        RECT 106.680 209.950 106.960 210.230 ;
        RECT 110.120 209.950 110.400 210.230 ;
        RECT 110.640 209.950 110.920 210.230 ;
        RECT 21.760 209.260 22.040 209.540 ;
        RECT 22.280 209.260 22.560 209.540 ;
        RECT 46.960 209.260 47.240 209.540 ;
        RECT 47.480 209.260 47.760 209.540 ;
        RECT 72.160 209.260 72.440 209.540 ;
        RECT 72.680 209.260 72.960 209.540 ;
        RECT 97.360 209.260 97.640 209.540 ;
        RECT 97.880 209.260 98.160 209.540 ;
        RECT 106.000 209.070 106.280 209.350 ;
        RECT 106.520 209.070 106.800 209.350 ;
        RECT 118.600 209.070 118.880 209.350 ;
        RECT 119.120 209.070 119.400 209.350 ;
        RECT 122.560 209.070 122.840 209.350 ;
        RECT 123.080 209.070 123.360 209.350 ;
        RECT 17.800 208.190 18.080 208.470 ;
        RECT 18.320 208.190 18.600 208.470 ;
        RECT 21.760 208.190 22.040 208.470 ;
        RECT 22.280 208.190 22.560 208.470 ;
        RECT 30.560 208.190 30.840 208.470 ;
        RECT 31.080 208.190 31.360 208.470 ;
        RECT 17.800 207.310 18.080 207.590 ;
        RECT 18.320 207.310 18.600 207.590 ;
        RECT 34.520 208.190 34.800 208.470 ;
        RECT 35.040 208.190 35.320 208.470 ;
        RECT 43.000 208.190 43.280 208.470 ;
        RECT 43.520 208.190 43.800 208.470 ;
        RECT 46.960 208.190 47.240 208.470 ;
        RECT 47.480 208.190 47.760 208.470 ;
        RECT 55.760 208.190 56.040 208.470 ;
        RECT 56.280 208.190 56.560 208.470 ;
        RECT 34.520 207.310 34.800 207.590 ;
        RECT 35.040 207.310 35.320 207.590 ;
        RECT 43.000 207.310 43.280 207.590 ;
        RECT 43.520 207.310 43.800 207.590 ;
        RECT 36.520 206.870 36.800 207.150 ;
        RECT 37.040 206.870 37.320 207.150 ;
        RECT 59.720 208.190 60.000 208.470 ;
        RECT 60.240 208.190 60.520 208.470 ;
        RECT 68.200 208.190 68.480 208.470 ;
        RECT 68.720 208.190 69.000 208.470 ;
        RECT 72.160 208.190 72.440 208.470 ;
        RECT 72.680 208.190 72.960 208.470 ;
        RECT 80.960 208.190 81.240 208.470 ;
        RECT 81.480 208.190 81.760 208.470 ;
        RECT 59.720 207.310 60.000 207.590 ;
        RECT 60.240 207.310 60.520 207.590 ;
        RECT 68.200 207.310 68.480 207.590 ;
        RECT 68.720 207.310 69.000 207.590 ;
        RECT 61.720 206.870 62.000 207.150 ;
        RECT 62.240 206.870 62.520 207.150 ;
        RECT 84.920 208.190 85.200 208.470 ;
        RECT 85.440 208.190 85.720 208.470 ;
        RECT 93.400 208.190 93.680 208.470 ;
        RECT 93.920 208.190 94.200 208.470 ;
        RECT 97.360 208.190 97.640 208.470 ;
        RECT 97.880 208.190 98.160 208.470 ;
        RECT 106.160 208.190 106.440 208.470 ;
        RECT 106.680 208.190 106.960 208.470 ;
        RECT 110.120 208.190 110.400 208.470 ;
        RECT 110.640 208.190 110.920 208.470 ;
        RECT 118.600 208.190 118.880 208.470 ;
        RECT 119.120 208.190 119.400 208.470 ;
        RECT 122.560 208.190 122.840 208.470 ;
        RECT 123.080 208.190 123.360 208.470 ;
        RECT 84.920 207.310 85.200 207.590 ;
        RECT 85.440 207.310 85.720 207.590 ;
        RECT 93.400 207.310 93.680 207.590 ;
        RECT 93.920 207.310 94.200 207.590 ;
        RECT 110.120 207.310 110.400 207.590 ;
        RECT 110.640 207.310 110.920 207.590 ;
        RECT 86.920 206.870 87.200 207.150 ;
        RECT 87.440 206.870 87.720 207.150 ;
        RECT 112.120 206.870 112.400 207.150 ;
        RECT 112.640 206.870 112.920 207.150 ;
        RECT 116.440 207.060 116.720 207.340 ;
        RECT 116.960 207.060 117.240 207.340 ;
        RECT 118.600 206.430 118.880 206.710 ;
        RECT 119.120 206.430 119.400 206.710 ;
        RECT 122.560 206.430 122.840 206.710 ;
        RECT 123.080 206.430 123.360 206.710 ;
        RECT 118.600 205.550 118.880 205.830 ;
        RECT 119.120 205.550 119.400 205.830 ;
        RECT 124.800 205.110 125.080 205.390 ;
        RECT 125.320 205.110 125.600 205.390 ;
        RECT 17.800 204.670 18.080 204.950 ;
        RECT 18.320 204.670 18.600 204.950 ;
        RECT 21.760 204.670 22.040 204.950 ;
        RECT 22.280 204.670 22.560 204.950 ;
        RECT 30.560 204.670 30.840 204.950 ;
        RECT 31.080 204.670 31.360 204.950 ;
        RECT 34.520 204.670 34.800 204.950 ;
        RECT 35.040 204.670 35.320 204.950 ;
        RECT 43.000 204.670 43.280 204.950 ;
        RECT 43.520 204.670 43.800 204.950 ;
        RECT 46.960 204.670 47.240 204.950 ;
        RECT 47.480 204.670 47.760 204.950 ;
        RECT 55.760 204.670 56.040 204.950 ;
        RECT 56.280 204.670 56.560 204.950 ;
        RECT 59.720 204.670 60.000 204.950 ;
        RECT 60.240 204.670 60.520 204.950 ;
        RECT 68.200 204.670 68.480 204.950 ;
        RECT 68.720 204.670 69.000 204.950 ;
        RECT 72.160 204.670 72.440 204.950 ;
        RECT 72.680 204.670 72.960 204.950 ;
        RECT 80.960 204.670 81.240 204.950 ;
        RECT 81.480 204.670 81.760 204.950 ;
        RECT 84.920 204.670 85.200 204.950 ;
        RECT 85.440 204.670 85.720 204.950 ;
        RECT 93.400 204.670 93.680 204.950 ;
        RECT 93.920 204.670 94.200 204.950 ;
        RECT 97.360 204.670 97.640 204.950 ;
        RECT 97.880 204.670 98.160 204.950 ;
        RECT 106.160 204.670 106.440 204.950 ;
        RECT 106.680 204.670 106.960 204.950 ;
        RECT 110.120 204.670 110.400 204.950 ;
        RECT 110.640 204.670 110.920 204.950 ;
        RECT 124.720 203.350 125.000 203.630 ;
        RECT 125.240 203.350 125.520 203.630 ;
        RECT 17.800 202.910 18.080 203.190 ;
        RECT 18.320 202.910 18.600 203.190 ;
        RECT 21.760 202.910 22.040 203.190 ;
        RECT 22.280 202.910 22.560 203.190 ;
        RECT 30.560 202.910 30.840 203.190 ;
        RECT 31.080 202.910 31.360 203.190 ;
        RECT 34.520 202.910 34.800 203.190 ;
        RECT 35.040 202.910 35.320 203.190 ;
        RECT 43.000 202.910 43.280 203.190 ;
        RECT 43.520 202.910 43.800 203.190 ;
        RECT 46.960 202.910 47.240 203.190 ;
        RECT 47.480 202.910 47.760 203.190 ;
        RECT 55.760 202.910 56.040 203.190 ;
        RECT 56.280 202.910 56.560 203.190 ;
        RECT 59.720 202.910 60.000 203.190 ;
        RECT 60.240 202.910 60.520 203.190 ;
        RECT 68.200 202.910 68.480 203.190 ;
        RECT 68.720 202.910 69.000 203.190 ;
        RECT 72.160 202.910 72.440 203.190 ;
        RECT 72.680 202.910 72.960 203.190 ;
        RECT 80.960 202.910 81.240 203.190 ;
        RECT 81.480 202.910 81.760 203.190 ;
        RECT 84.920 202.910 85.200 203.190 ;
        RECT 85.440 202.910 85.720 203.190 ;
        RECT 93.400 202.910 93.680 203.190 ;
        RECT 93.920 202.910 94.200 203.190 ;
        RECT 97.360 202.910 97.640 203.190 ;
        RECT 97.880 202.910 98.160 203.190 ;
        RECT 106.160 202.910 106.440 203.190 ;
        RECT 106.680 202.910 106.960 203.190 ;
        RECT 110.120 202.910 110.400 203.190 ;
        RECT 110.640 202.910 110.920 203.190 ;
        RECT 118.600 202.910 118.880 203.190 ;
        RECT 119.120 202.910 119.400 203.190 ;
        RECT 122.560 202.910 122.840 203.190 ;
        RECT 123.080 202.910 123.360 203.190 ;
        RECT 21.760 202.030 22.040 202.310 ;
        RECT 22.280 202.030 22.560 202.310 ;
        RECT 30.560 202.030 30.840 202.310 ;
        RECT 31.080 202.030 31.360 202.310 ;
        RECT 46.960 202.030 47.240 202.310 ;
        RECT 47.480 202.030 47.760 202.310 ;
        RECT 55.760 202.030 56.040 202.310 ;
        RECT 56.280 202.030 56.560 202.310 ;
        RECT 72.160 202.030 72.440 202.310 ;
        RECT 72.680 202.030 72.960 202.310 ;
        RECT 80.960 202.030 81.240 202.310 ;
        RECT 81.480 202.030 81.760 202.310 ;
        RECT 97.360 202.030 97.640 202.310 ;
        RECT 97.880 202.030 98.160 202.310 ;
        RECT 106.160 202.030 106.440 202.310 ;
        RECT 106.680 202.030 106.960 202.310 ;
        RECT 122.560 202.030 122.840 202.310 ;
        RECT 123.080 202.030 123.360 202.310 ;
        RECT 17.800 199.390 18.080 199.670 ;
        RECT 18.320 199.390 18.600 199.670 ;
        RECT 21.760 199.390 22.040 199.670 ;
        RECT 22.280 199.390 22.560 199.670 ;
        RECT 30.560 199.390 30.840 199.670 ;
        RECT 31.080 199.390 31.360 199.670 ;
        RECT 34.520 199.390 34.800 199.670 ;
        RECT 35.040 199.390 35.320 199.670 ;
        RECT 17.800 197.630 18.080 197.910 ;
        RECT 18.320 197.630 18.600 197.910 ;
        RECT 21.760 197.630 22.040 197.910 ;
        RECT 22.280 197.630 22.560 197.910 ;
        RECT 30.560 197.630 30.840 197.910 ;
        RECT 31.080 197.630 31.360 197.910 ;
        RECT 34.520 197.630 34.800 197.910 ;
        RECT 35.040 197.630 35.320 197.910 ;
        RECT 17.800 195.870 18.080 196.150 ;
        RECT 18.320 195.870 18.600 196.150 ;
        RECT 21.760 195.870 22.040 196.150 ;
        RECT 22.280 195.870 22.560 196.150 ;
        RECT 17.800 192.350 18.080 192.630 ;
        RECT 18.320 192.350 18.600 192.630 ;
        RECT 21.760 192.350 22.040 192.630 ;
        RECT 22.280 192.350 22.560 192.630 ;
        RECT 17.800 191.470 18.080 191.750 ;
        RECT 18.320 191.470 18.600 191.750 ;
        RECT 21.760 191.470 22.040 191.750 ;
        RECT 22.280 191.470 22.560 191.750 ;
        RECT 15.640 191.030 15.920 191.310 ;
        RECT 16.160 191.030 16.440 191.310 ;
        RECT 17.800 188.830 18.080 189.110 ;
        RECT 18.320 188.830 18.600 189.110 ;
        RECT 17.800 187.950 18.080 188.230 ;
        RECT 18.320 187.950 18.600 188.230 ;
        RECT 21.760 187.950 22.040 188.230 ;
        RECT 22.280 187.950 22.560 188.230 ;
        RECT 17.800 185.310 18.080 185.590 ;
        RECT 18.320 185.310 18.600 185.590 ;
        RECT 17.800 184.430 18.080 184.710 ;
        RECT 18.320 184.430 18.600 184.710 ;
        RECT 21.760 184.430 22.040 184.710 ;
        RECT 22.280 184.430 22.560 184.710 ;
        RECT 20.940 182.870 21.220 183.150 ;
        RECT 20.940 182.350 21.220 182.630 ;
        RECT 17.800 181.790 18.080 182.070 ;
        RECT 18.320 181.790 18.600 182.070 ;
        RECT 21.760 181.790 22.040 182.070 ;
        RECT 22.280 181.790 22.560 182.070 ;
        RECT 17.800 180.910 18.080 181.190 ;
        RECT 18.320 180.910 18.600 181.190 ;
        RECT 21.760 180.910 22.040 181.190 ;
        RECT 22.280 180.910 22.560 181.190 ;
        RECT 17.800 178.270 18.080 178.550 ;
        RECT 18.320 178.270 18.600 178.550 ;
        RECT 17.800 177.390 18.080 177.670 ;
        RECT 18.320 177.390 18.600 177.670 ;
        RECT 21.760 177.390 22.040 177.670 ;
        RECT 22.280 177.390 22.560 177.670 ;
        RECT 20.065 175.830 20.345 176.110 ;
        RECT 20.065 175.310 20.345 175.590 ;
        RECT 15.720 168.110 16.000 168.390 ;
        RECT 16.240 168.110 16.520 168.390 ;
        RECT 15.640 159.350 15.920 159.630 ;
        RECT 16.160 159.350 16.440 159.630 ;
        RECT 15.640 155.830 15.920 156.110 ;
        RECT 16.160 155.830 16.440 156.110 ;
        RECT 17.800 174.750 18.080 175.030 ;
        RECT 18.320 174.750 18.600 175.030 ;
        RECT 21.760 174.750 22.040 175.030 ;
        RECT 22.280 174.750 22.560 175.030 ;
        RECT 17.800 173.870 18.080 174.150 ;
        RECT 18.320 173.870 18.600 174.150 ;
        RECT 21.760 173.870 22.040 174.150 ;
        RECT 22.280 173.870 22.560 174.150 ;
        RECT 17.800 171.230 18.080 171.510 ;
        RECT 18.320 171.230 18.600 171.510 ;
        RECT 17.800 170.350 18.080 170.630 ;
        RECT 18.320 170.350 18.600 170.630 ;
        RECT 21.760 170.350 22.040 170.630 ;
        RECT 22.280 170.350 22.560 170.630 ;
        RECT 19.265 168.790 19.545 169.070 ;
        RECT 19.265 168.270 19.545 168.550 ;
        RECT 17.800 167.710 18.080 167.990 ;
        RECT 18.320 167.710 18.600 167.990 ;
        RECT 21.760 167.710 22.040 167.990 ;
        RECT 22.280 167.710 22.560 167.990 ;
        RECT 17.800 166.830 18.080 167.110 ;
        RECT 18.320 166.830 18.600 167.110 ;
        RECT 21.760 166.830 22.040 167.110 ;
        RECT 22.280 166.830 22.560 167.110 ;
        RECT 17.800 164.190 18.080 164.470 ;
        RECT 18.320 164.190 18.600 164.470 ;
        RECT 17.800 163.310 18.080 163.590 ;
        RECT 18.320 163.310 18.600 163.590 ;
        RECT 21.760 163.310 22.040 163.590 ;
        RECT 22.280 163.310 22.560 163.590 ;
        RECT 17.800 160.670 18.080 160.950 ;
        RECT 18.320 160.670 18.600 160.950 ;
        RECT 21.760 160.670 22.040 160.950 ;
        RECT 22.280 160.670 22.560 160.950 ;
        RECT 23.920 159.350 24.200 159.630 ;
        RECT 24.440 159.350 24.720 159.630 ;
        RECT 17.800 155.390 18.080 155.670 ;
        RECT 18.320 155.390 18.600 155.670 ;
        RECT 21.760 155.390 22.040 155.670 ;
        RECT 22.280 155.390 22.560 155.670 ;
        RECT 15.720 150.510 16.000 150.790 ;
        RECT 16.240 150.510 16.520 150.790 ;
        RECT 17.800 150.110 18.080 150.390 ;
        RECT 18.320 150.110 18.600 150.390 ;
        RECT 21.760 150.110 22.040 150.390 ;
        RECT 22.280 150.110 22.560 150.390 ;
        RECT 17.800 148.350 18.080 148.630 ;
        RECT 18.320 148.350 18.600 148.630 ;
        RECT 21.760 148.350 22.040 148.630 ;
        RECT 22.280 148.350 22.560 148.630 ;
        RECT 21.760 147.470 22.040 147.750 ;
        RECT 22.280 147.470 22.560 147.750 ;
        RECT 17.800 146.590 18.080 146.870 ;
        RECT 18.320 146.590 18.600 146.870 ;
        RECT 17.800 145.710 18.080 145.990 ;
        RECT 18.320 145.710 18.600 145.990 ;
        RECT 17.800 143.070 18.080 143.350 ;
        RECT 18.320 143.070 18.600 143.350 ;
        RECT 21.840 143.030 22.120 143.310 ;
        RECT 22.360 143.030 22.640 143.310 ;
        RECT 30.560 195.870 30.840 196.150 ;
        RECT 31.080 195.870 31.360 196.150 ;
        RECT 34.520 195.870 34.800 196.150 ;
        RECT 35.040 195.870 35.320 196.150 ;
        RECT 43.000 199.390 43.280 199.670 ;
        RECT 43.520 199.390 43.800 199.670 ;
        RECT 46.960 199.390 47.240 199.670 ;
        RECT 47.480 199.390 47.760 199.670 ;
        RECT 55.760 199.390 56.040 199.670 ;
        RECT 56.280 199.390 56.560 199.670 ;
        RECT 59.720 199.390 60.000 199.670 ;
        RECT 60.240 199.390 60.520 199.670 ;
        RECT 43.000 197.630 43.280 197.910 ;
        RECT 43.520 197.630 43.800 197.910 ;
        RECT 46.960 197.630 47.240 197.910 ;
        RECT 47.480 197.630 47.760 197.910 ;
        RECT 55.760 197.630 56.040 197.910 ;
        RECT 56.280 197.630 56.560 197.910 ;
        RECT 59.720 197.630 60.000 197.910 ;
        RECT 60.240 197.630 60.520 197.910 ;
        RECT 43.000 195.870 43.280 196.150 ;
        RECT 43.520 195.870 43.800 196.150 ;
        RECT 46.960 195.870 47.240 196.150 ;
        RECT 47.480 195.870 47.760 196.150 ;
        RECT 30.560 192.350 30.840 192.630 ;
        RECT 31.080 192.350 31.360 192.630 ;
        RECT 34.520 192.350 34.800 192.630 ;
        RECT 35.040 192.350 35.320 192.630 ;
        RECT 43.000 192.350 43.280 192.630 ;
        RECT 43.520 192.350 43.800 192.630 ;
        RECT 46.960 192.350 47.240 192.630 ;
        RECT 47.480 192.350 47.760 192.630 ;
        RECT 30.560 191.470 30.840 191.750 ;
        RECT 31.080 191.470 31.360 191.750 ;
        RECT 34.520 191.470 34.800 191.750 ;
        RECT 35.040 191.470 35.320 191.750 ;
        RECT 43.000 191.470 43.280 191.750 ;
        RECT 43.520 191.470 43.800 191.750 ;
        RECT 46.960 191.470 47.240 191.750 ;
        RECT 47.480 191.470 47.760 191.750 ;
        RECT 36.520 191.030 36.800 191.310 ;
        RECT 37.040 191.030 37.320 191.310 ;
        RECT 40.840 191.030 41.120 191.310 ;
        RECT 41.360 191.030 41.640 191.310 ;
        RECT 34.520 188.830 34.800 189.110 ;
        RECT 35.040 188.830 35.320 189.110 ;
        RECT 43.000 188.830 43.280 189.110 ;
        RECT 43.520 188.830 43.800 189.110 ;
        RECT 30.560 187.950 30.840 188.230 ;
        RECT 31.080 187.950 31.360 188.230 ;
        RECT 34.520 187.950 34.800 188.230 ;
        RECT 35.040 187.950 35.320 188.230 ;
        RECT 43.000 187.950 43.280 188.230 ;
        RECT 43.520 187.950 43.800 188.230 ;
        RECT 46.960 187.950 47.240 188.230 ;
        RECT 47.480 187.950 47.760 188.230 ;
        RECT 34.520 185.310 34.800 185.590 ;
        RECT 35.040 185.310 35.320 185.590 ;
        RECT 43.000 185.310 43.280 185.590 ;
        RECT 43.520 185.310 43.800 185.590 ;
        RECT 30.560 184.430 30.840 184.710 ;
        RECT 31.080 184.430 31.360 184.710 ;
        RECT 34.520 184.430 34.800 184.710 ;
        RECT 35.040 184.430 35.320 184.710 ;
        RECT 43.000 184.430 43.280 184.710 ;
        RECT 43.520 184.430 43.800 184.710 ;
        RECT 46.960 184.430 47.240 184.710 ;
        RECT 47.480 184.430 47.760 184.710 ;
        RECT 31.900 182.870 32.180 183.150 ;
        RECT 31.900 182.350 32.180 182.630 ;
        RECT 46.140 182.870 46.420 183.150 ;
        RECT 46.140 182.350 46.420 182.630 ;
        RECT 30.560 181.790 30.840 182.070 ;
        RECT 31.080 181.790 31.360 182.070 ;
        RECT 34.520 181.790 34.800 182.070 ;
        RECT 35.040 181.790 35.320 182.070 ;
        RECT 43.000 181.790 43.280 182.070 ;
        RECT 43.520 181.790 43.800 182.070 ;
        RECT 46.960 181.790 47.240 182.070 ;
        RECT 47.480 181.790 47.760 182.070 ;
        RECT 30.560 180.910 30.840 181.190 ;
        RECT 31.080 180.910 31.360 181.190 ;
        RECT 34.520 180.910 34.800 181.190 ;
        RECT 35.040 180.910 35.320 181.190 ;
        RECT 43.000 180.910 43.280 181.190 ;
        RECT 43.520 180.910 43.800 181.190 ;
        RECT 46.960 180.910 47.240 181.190 ;
        RECT 47.480 180.910 47.760 181.190 ;
        RECT 34.520 178.270 34.800 178.550 ;
        RECT 35.040 178.270 35.320 178.550 ;
        RECT 43.000 178.270 43.280 178.550 ;
        RECT 43.520 178.270 43.800 178.550 ;
        RECT 30.560 177.390 30.840 177.670 ;
        RECT 31.080 177.390 31.360 177.670 ;
        RECT 34.520 177.390 34.800 177.670 ;
        RECT 35.040 177.390 35.320 177.670 ;
        RECT 43.000 177.390 43.280 177.670 ;
        RECT 43.520 177.390 43.800 177.670 ;
        RECT 46.960 177.390 47.240 177.670 ;
        RECT 47.480 177.390 47.760 177.670 ;
        RECT 32.775 175.830 33.055 176.110 ;
        RECT 32.775 175.310 33.055 175.590 ;
        RECT 45.265 175.830 45.545 176.110 ;
        RECT 45.265 175.310 45.545 175.590 ;
        RECT 30.560 174.750 30.840 175.030 ;
        RECT 31.080 174.750 31.360 175.030 ;
        RECT 34.520 174.750 34.800 175.030 ;
        RECT 35.040 174.750 35.320 175.030 ;
        RECT 30.560 173.870 30.840 174.150 ;
        RECT 31.080 173.870 31.360 174.150 ;
        RECT 34.520 173.870 34.800 174.150 ;
        RECT 35.040 173.870 35.320 174.150 ;
        RECT 34.520 171.230 34.800 171.510 ;
        RECT 35.040 171.230 35.320 171.510 ;
        RECT 30.560 170.350 30.840 170.630 ;
        RECT 31.080 170.350 31.360 170.630 ;
        RECT 34.520 170.350 34.800 170.630 ;
        RECT 35.040 170.350 35.320 170.630 ;
        RECT 33.575 168.790 33.855 169.070 ;
        RECT 33.575 168.270 33.855 168.550 ;
        RECT 30.560 167.710 30.840 167.990 ;
        RECT 31.080 167.710 31.360 167.990 ;
        RECT 34.520 167.710 34.800 167.990 ;
        RECT 35.040 167.710 35.320 167.990 ;
        RECT 30.560 166.830 30.840 167.110 ;
        RECT 31.080 166.830 31.360 167.110 ;
        RECT 34.520 166.830 34.800 167.110 ;
        RECT 35.040 166.830 35.320 167.110 ;
        RECT 34.520 164.190 34.800 164.470 ;
        RECT 35.040 164.190 35.320 164.470 ;
        RECT 30.560 163.310 30.840 163.590 ;
        RECT 31.080 163.310 31.360 163.590 ;
        RECT 34.520 163.310 34.800 163.590 ;
        RECT 35.040 163.310 35.320 163.590 ;
        RECT 30.560 160.670 30.840 160.950 ;
        RECT 31.080 160.670 31.360 160.950 ;
        RECT 34.520 160.670 34.800 160.950 ;
        RECT 35.040 160.670 35.320 160.950 ;
        RECT 28.240 159.350 28.520 159.630 ;
        RECT 28.760 159.350 29.040 159.630 ;
        RECT 30.560 155.390 30.840 155.670 ;
        RECT 31.080 155.390 31.360 155.670 ;
        RECT 34.520 155.390 34.800 155.670 ;
        RECT 35.040 155.390 35.320 155.670 ;
        RECT 36.600 168.110 36.880 168.390 ;
        RECT 37.120 168.110 37.400 168.390 ;
        RECT 40.920 168.110 41.200 168.390 ;
        RECT 41.440 168.110 41.720 168.390 ;
        RECT 36.520 155.830 36.800 156.110 ;
        RECT 37.040 155.830 37.320 156.110 ;
        RECT 30.560 150.110 30.840 150.390 ;
        RECT 31.080 150.110 31.360 150.390 ;
        RECT 34.520 150.110 34.800 150.390 ;
        RECT 35.040 150.110 35.320 150.390 ;
        RECT 30.560 148.350 30.840 148.630 ;
        RECT 31.080 148.350 31.360 148.630 ;
        RECT 34.520 148.350 34.800 148.630 ;
        RECT 35.040 148.350 35.320 148.630 ;
        RECT 30.560 147.470 30.840 147.750 ;
        RECT 31.080 147.470 31.360 147.750 ;
        RECT 34.520 146.590 34.800 146.870 ;
        RECT 35.040 146.590 35.320 146.870 ;
        RECT 34.520 145.710 34.800 145.990 ;
        RECT 35.040 145.710 35.320 145.990 ;
        RECT 36.600 150.510 36.880 150.790 ;
        RECT 37.120 150.510 37.400 150.790 ;
        RECT 30.480 143.030 30.760 143.310 ;
        RECT 31.000 143.030 31.280 143.310 ;
        RECT 34.520 143.070 34.800 143.350 ;
        RECT 35.040 143.070 35.320 143.350 ;
        RECT 21.760 142.190 22.040 142.470 ;
        RECT 22.280 142.190 22.560 142.470 ;
        RECT 30.560 142.190 30.840 142.470 ;
        RECT 31.080 142.190 31.360 142.470 ;
        RECT 15.720 141.710 16.000 141.990 ;
        RECT 16.240 141.710 16.520 141.990 ;
        RECT 36.600 141.710 36.880 141.990 ;
        RECT 37.120 141.710 37.400 141.990 ;
        RECT 40.840 155.830 41.120 156.110 ;
        RECT 41.360 155.830 41.640 156.110 ;
        RECT 43.000 174.750 43.280 175.030 ;
        RECT 43.520 174.750 43.800 175.030 ;
        RECT 46.960 174.750 47.240 175.030 ;
        RECT 47.480 174.750 47.760 175.030 ;
        RECT 43.000 173.870 43.280 174.150 ;
        RECT 43.520 173.870 43.800 174.150 ;
        RECT 46.960 173.870 47.240 174.150 ;
        RECT 47.480 173.870 47.760 174.150 ;
        RECT 43.000 171.230 43.280 171.510 ;
        RECT 43.520 171.230 43.800 171.510 ;
        RECT 43.000 170.350 43.280 170.630 ;
        RECT 43.520 170.350 43.800 170.630 ;
        RECT 46.960 170.350 47.240 170.630 ;
        RECT 47.480 170.350 47.760 170.630 ;
        RECT 44.465 168.790 44.745 169.070 ;
        RECT 44.465 168.270 44.745 168.550 ;
        RECT 43.000 167.710 43.280 167.990 ;
        RECT 43.520 167.710 43.800 167.990 ;
        RECT 46.960 167.710 47.240 167.990 ;
        RECT 47.480 167.710 47.760 167.990 ;
        RECT 43.000 166.830 43.280 167.110 ;
        RECT 43.520 166.830 43.800 167.110 ;
        RECT 46.960 166.830 47.240 167.110 ;
        RECT 47.480 166.830 47.760 167.110 ;
        RECT 43.000 164.190 43.280 164.470 ;
        RECT 43.520 164.190 43.800 164.470 ;
        RECT 43.000 163.310 43.280 163.590 ;
        RECT 43.520 163.310 43.800 163.590 ;
        RECT 46.960 163.310 47.240 163.590 ;
        RECT 47.480 163.310 47.760 163.590 ;
        RECT 43.000 160.670 43.280 160.950 ;
        RECT 43.520 160.670 43.800 160.950 ;
        RECT 46.960 160.670 47.240 160.950 ;
        RECT 47.480 160.670 47.760 160.950 ;
        RECT 49.120 159.350 49.400 159.630 ;
        RECT 49.640 159.350 49.920 159.630 ;
        RECT 43.000 155.390 43.280 155.670 ;
        RECT 43.520 155.390 43.800 155.670 ;
        RECT 46.960 155.390 47.240 155.670 ;
        RECT 47.480 155.390 47.760 155.670 ;
        RECT 40.920 150.510 41.200 150.790 ;
        RECT 41.440 150.510 41.720 150.790 ;
        RECT 43.000 150.110 43.280 150.390 ;
        RECT 43.520 150.110 43.800 150.390 ;
        RECT 46.960 150.110 47.240 150.390 ;
        RECT 47.480 150.110 47.760 150.390 ;
        RECT 43.000 148.350 43.280 148.630 ;
        RECT 43.520 148.350 43.800 148.630 ;
        RECT 46.960 148.350 47.240 148.630 ;
        RECT 47.480 148.350 47.760 148.630 ;
        RECT 46.960 147.470 47.240 147.750 ;
        RECT 47.480 147.470 47.760 147.750 ;
        RECT 43.000 146.590 43.280 146.870 ;
        RECT 43.520 146.590 43.800 146.870 ;
        RECT 43.000 145.710 43.280 145.990 ;
        RECT 43.520 145.710 43.800 145.990 ;
        RECT 43.000 143.070 43.280 143.350 ;
        RECT 43.520 143.070 43.800 143.350 ;
        RECT 47.040 143.030 47.320 143.310 ;
        RECT 47.560 143.030 47.840 143.310 ;
        RECT 55.760 195.870 56.040 196.150 ;
        RECT 56.280 195.870 56.560 196.150 ;
        RECT 59.720 195.870 60.000 196.150 ;
        RECT 60.240 195.870 60.520 196.150 ;
        RECT 68.200 199.390 68.480 199.670 ;
        RECT 68.720 199.390 69.000 199.670 ;
        RECT 72.160 199.390 72.440 199.670 ;
        RECT 72.680 199.390 72.960 199.670 ;
        RECT 80.960 199.390 81.240 199.670 ;
        RECT 81.480 199.390 81.760 199.670 ;
        RECT 84.920 199.390 85.200 199.670 ;
        RECT 85.440 199.390 85.720 199.670 ;
        RECT 68.200 197.630 68.480 197.910 ;
        RECT 68.720 197.630 69.000 197.910 ;
        RECT 72.160 197.630 72.440 197.910 ;
        RECT 72.680 197.630 72.960 197.910 ;
        RECT 80.960 197.630 81.240 197.910 ;
        RECT 81.480 197.630 81.760 197.910 ;
        RECT 84.920 197.630 85.200 197.910 ;
        RECT 85.440 197.630 85.720 197.910 ;
        RECT 68.200 195.870 68.480 196.150 ;
        RECT 68.720 195.870 69.000 196.150 ;
        RECT 72.160 195.870 72.440 196.150 ;
        RECT 72.680 195.870 72.960 196.150 ;
        RECT 55.760 192.350 56.040 192.630 ;
        RECT 56.280 192.350 56.560 192.630 ;
        RECT 59.720 192.350 60.000 192.630 ;
        RECT 60.240 192.350 60.520 192.630 ;
        RECT 68.200 192.350 68.480 192.630 ;
        RECT 68.720 192.350 69.000 192.630 ;
        RECT 72.160 192.350 72.440 192.630 ;
        RECT 72.680 192.350 72.960 192.630 ;
        RECT 55.760 191.470 56.040 191.750 ;
        RECT 56.280 191.470 56.560 191.750 ;
        RECT 59.720 191.470 60.000 191.750 ;
        RECT 60.240 191.470 60.520 191.750 ;
        RECT 68.200 191.470 68.480 191.750 ;
        RECT 68.720 191.470 69.000 191.750 ;
        RECT 72.160 191.470 72.440 191.750 ;
        RECT 72.680 191.470 72.960 191.750 ;
        RECT 61.720 191.030 62.000 191.310 ;
        RECT 62.240 191.030 62.520 191.310 ;
        RECT 66.040 191.030 66.320 191.310 ;
        RECT 66.560 191.030 66.840 191.310 ;
        RECT 59.720 188.830 60.000 189.110 ;
        RECT 60.240 188.830 60.520 189.110 ;
        RECT 68.200 188.830 68.480 189.110 ;
        RECT 68.720 188.830 69.000 189.110 ;
        RECT 55.760 187.950 56.040 188.230 ;
        RECT 56.280 187.950 56.560 188.230 ;
        RECT 59.720 187.950 60.000 188.230 ;
        RECT 60.240 187.950 60.520 188.230 ;
        RECT 68.200 187.950 68.480 188.230 ;
        RECT 68.720 187.950 69.000 188.230 ;
        RECT 72.160 187.950 72.440 188.230 ;
        RECT 72.680 187.950 72.960 188.230 ;
        RECT 59.720 185.310 60.000 185.590 ;
        RECT 60.240 185.310 60.520 185.590 ;
        RECT 68.200 185.310 68.480 185.590 ;
        RECT 68.720 185.310 69.000 185.590 ;
        RECT 55.760 184.430 56.040 184.710 ;
        RECT 56.280 184.430 56.560 184.710 ;
        RECT 59.720 184.430 60.000 184.710 ;
        RECT 60.240 184.430 60.520 184.710 ;
        RECT 68.200 184.430 68.480 184.710 ;
        RECT 68.720 184.430 69.000 184.710 ;
        RECT 72.160 184.430 72.440 184.710 ;
        RECT 72.680 184.430 72.960 184.710 ;
        RECT 57.100 182.870 57.380 183.150 ;
        RECT 57.100 182.350 57.380 182.630 ;
        RECT 71.340 182.870 71.620 183.150 ;
        RECT 71.340 182.350 71.620 182.630 ;
        RECT 55.760 181.790 56.040 182.070 ;
        RECT 56.280 181.790 56.560 182.070 ;
        RECT 59.720 181.790 60.000 182.070 ;
        RECT 60.240 181.790 60.520 182.070 ;
        RECT 68.200 181.790 68.480 182.070 ;
        RECT 68.720 181.790 69.000 182.070 ;
        RECT 72.160 181.790 72.440 182.070 ;
        RECT 72.680 181.790 72.960 182.070 ;
        RECT 55.760 180.910 56.040 181.190 ;
        RECT 56.280 180.910 56.560 181.190 ;
        RECT 59.720 180.910 60.000 181.190 ;
        RECT 60.240 180.910 60.520 181.190 ;
        RECT 68.200 180.910 68.480 181.190 ;
        RECT 68.720 180.910 69.000 181.190 ;
        RECT 72.160 180.910 72.440 181.190 ;
        RECT 72.680 180.910 72.960 181.190 ;
        RECT 59.720 178.270 60.000 178.550 ;
        RECT 60.240 178.270 60.520 178.550 ;
        RECT 68.200 178.270 68.480 178.550 ;
        RECT 68.720 178.270 69.000 178.550 ;
        RECT 55.760 177.390 56.040 177.670 ;
        RECT 56.280 177.390 56.560 177.670 ;
        RECT 59.720 177.390 60.000 177.670 ;
        RECT 60.240 177.390 60.520 177.670 ;
        RECT 68.200 177.390 68.480 177.670 ;
        RECT 68.720 177.390 69.000 177.670 ;
        RECT 72.160 177.390 72.440 177.670 ;
        RECT 72.680 177.390 72.960 177.670 ;
        RECT 57.975 175.830 58.255 176.110 ;
        RECT 57.975 175.310 58.255 175.590 ;
        RECT 70.465 175.830 70.745 176.110 ;
        RECT 70.465 175.310 70.745 175.590 ;
        RECT 55.760 174.750 56.040 175.030 ;
        RECT 56.280 174.750 56.560 175.030 ;
        RECT 59.720 174.750 60.000 175.030 ;
        RECT 60.240 174.750 60.520 175.030 ;
        RECT 55.760 173.870 56.040 174.150 ;
        RECT 56.280 173.870 56.560 174.150 ;
        RECT 59.720 173.870 60.000 174.150 ;
        RECT 60.240 173.870 60.520 174.150 ;
        RECT 59.720 171.230 60.000 171.510 ;
        RECT 60.240 171.230 60.520 171.510 ;
        RECT 55.760 170.350 56.040 170.630 ;
        RECT 56.280 170.350 56.560 170.630 ;
        RECT 59.720 170.350 60.000 170.630 ;
        RECT 60.240 170.350 60.520 170.630 ;
        RECT 58.775 168.790 59.055 169.070 ;
        RECT 58.775 168.270 59.055 168.550 ;
        RECT 55.760 167.710 56.040 167.990 ;
        RECT 56.280 167.710 56.560 167.990 ;
        RECT 59.720 167.710 60.000 167.990 ;
        RECT 60.240 167.710 60.520 167.990 ;
        RECT 55.760 166.830 56.040 167.110 ;
        RECT 56.280 166.830 56.560 167.110 ;
        RECT 59.720 166.830 60.000 167.110 ;
        RECT 60.240 166.830 60.520 167.110 ;
        RECT 59.720 164.190 60.000 164.470 ;
        RECT 60.240 164.190 60.520 164.470 ;
        RECT 55.760 163.310 56.040 163.590 ;
        RECT 56.280 163.310 56.560 163.590 ;
        RECT 59.720 163.310 60.000 163.590 ;
        RECT 60.240 163.310 60.520 163.590 ;
        RECT 55.760 160.670 56.040 160.950 ;
        RECT 56.280 160.670 56.560 160.950 ;
        RECT 59.720 160.670 60.000 160.950 ;
        RECT 60.240 160.670 60.520 160.950 ;
        RECT 53.440 159.350 53.720 159.630 ;
        RECT 53.960 159.350 54.240 159.630 ;
        RECT 55.760 155.390 56.040 155.670 ;
        RECT 56.280 155.390 56.560 155.670 ;
        RECT 59.720 155.390 60.000 155.670 ;
        RECT 60.240 155.390 60.520 155.670 ;
        RECT 61.800 168.110 62.080 168.390 ;
        RECT 62.320 168.110 62.600 168.390 ;
        RECT 66.120 168.110 66.400 168.390 ;
        RECT 66.640 168.110 66.920 168.390 ;
        RECT 61.720 155.830 62.000 156.110 ;
        RECT 62.240 155.830 62.520 156.110 ;
        RECT 55.760 150.110 56.040 150.390 ;
        RECT 56.280 150.110 56.560 150.390 ;
        RECT 59.720 150.110 60.000 150.390 ;
        RECT 60.240 150.110 60.520 150.390 ;
        RECT 55.760 148.350 56.040 148.630 ;
        RECT 56.280 148.350 56.560 148.630 ;
        RECT 59.720 148.350 60.000 148.630 ;
        RECT 60.240 148.350 60.520 148.630 ;
        RECT 55.760 147.470 56.040 147.750 ;
        RECT 56.280 147.470 56.560 147.750 ;
        RECT 59.720 146.590 60.000 146.870 ;
        RECT 60.240 146.590 60.520 146.870 ;
        RECT 59.720 145.710 60.000 145.990 ;
        RECT 60.240 145.710 60.520 145.990 ;
        RECT 61.800 150.510 62.080 150.790 ;
        RECT 62.320 150.510 62.600 150.790 ;
        RECT 55.680 143.030 55.960 143.310 ;
        RECT 56.200 143.030 56.480 143.310 ;
        RECT 59.720 143.070 60.000 143.350 ;
        RECT 60.240 143.070 60.520 143.350 ;
        RECT 46.960 142.190 47.240 142.470 ;
        RECT 47.480 142.190 47.760 142.470 ;
        RECT 55.760 142.190 56.040 142.470 ;
        RECT 56.280 142.190 56.560 142.470 ;
        RECT 40.920 141.710 41.200 141.990 ;
        RECT 41.440 141.710 41.720 141.990 ;
        RECT 61.800 141.710 62.080 141.990 ;
        RECT 62.320 141.710 62.600 141.990 ;
        RECT 66.040 155.830 66.320 156.110 ;
        RECT 66.560 155.830 66.840 156.110 ;
        RECT 68.200 174.750 68.480 175.030 ;
        RECT 68.720 174.750 69.000 175.030 ;
        RECT 72.160 174.750 72.440 175.030 ;
        RECT 72.680 174.750 72.960 175.030 ;
        RECT 68.200 173.870 68.480 174.150 ;
        RECT 68.720 173.870 69.000 174.150 ;
        RECT 72.160 173.870 72.440 174.150 ;
        RECT 72.680 173.870 72.960 174.150 ;
        RECT 68.200 171.230 68.480 171.510 ;
        RECT 68.720 171.230 69.000 171.510 ;
        RECT 68.200 170.350 68.480 170.630 ;
        RECT 68.720 170.350 69.000 170.630 ;
        RECT 72.160 170.350 72.440 170.630 ;
        RECT 72.680 170.350 72.960 170.630 ;
        RECT 69.665 168.790 69.945 169.070 ;
        RECT 69.665 168.270 69.945 168.550 ;
        RECT 68.200 167.710 68.480 167.990 ;
        RECT 68.720 167.710 69.000 167.990 ;
        RECT 72.160 167.710 72.440 167.990 ;
        RECT 72.680 167.710 72.960 167.990 ;
        RECT 68.200 166.830 68.480 167.110 ;
        RECT 68.720 166.830 69.000 167.110 ;
        RECT 72.160 166.830 72.440 167.110 ;
        RECT 72.680 166.830 72.960 167.110 ;
        RECT 68.200 164.190 68.480 164.470 ;
        RECT 68.720 164.190 69.000 164.470 ;
        RECT 68.200 163.310 68.480 163.590 ;
        RECT 68.720 163.310 69.000 163.590 ;
        RECT 72.160 163.310 72.440 163.590 ;
        RECT 72.680 163.310 72.960 163.590 ;
        RECT 68.200 160.670 68.480 160.950 ;
        RECT 68.720 160.670 69.000 160.950 ;
        RECT 72.160 160.670 72.440 160.950 ;
        RECT 72.680 160.670 72.960 160.950 ;
        RECT 74.320 159.350 74.600 159.630 ;
        RECT 74.840 159.350 75.120 159.630 ;
        RECT 68.200 155.390 68.480 155.670 ;
        RECT 68.720 155.390 69.000 155.670 ;
        RECT 72.160 155.390 72.440 155.670 ;
        RECT 72.680 155.390 72.960 155.670 ;
        RECT 66.120 150.510 66.400 150.790 ;
        RECT 66.640 150.510 66.920 150.790 ;
        RECT 68.200 150.110 68.480 150.390 ;
        RECT 68.720 150.110 69.000 150.390 ;
        RECT 72.160 150.110 72.440 150.390 ;
        RECT 72.680 150.110 72.960 150.390 ;
        RECT 68.200 148.350 68.480 148.630 ;
        RECT 68.720 148.350 69.000 148.630 ;
        RECT 72.160 148.350 72.440 148.630 ;
        RECT 72.680 148.350 72.960 148.630 ;
        RECT 72.160 147.470 72.440 147.750 ;
        RECT 72.680 147.470 72.960 147.750 ;
        RECT 68.200 146.590 68.480 146.870 ;
        RECT 68.720 146.590 69.000 146.870 ;
        RECT 68.200 145.710 68.480 145.990 ;
        RECT 68.720 145.710 69.000 145.990 ;
        RECT 68.200 143.070 68.480 143.350 ;
        RECT 68.720 143.070 69.000 143.350 ;
        RECT 72.240 143.030 72.520 143.310 ;
        RECT 72.760 143.030 73.040 143.310 ;
        RECT 80.960 195.870 81.240 196.150 ;
        RECT 81.480 195.870 81.760 196.150 ;
        RECT 84.920 195.870 85.200 196.150 ;
        RECT 85.440 195.870 85.720 196.150 ;
        RECT 93.400 199.390 93.680 199.670 ;
        RECT 93.920 199.390 94.200 199.670 ;
        RECT 97.360 199.390 97.640 199.670 ;
        RECT 97.880 199.390 98.160 199.670 ;
        RECT 106.160 199.390 106.440 199.670 ;
        RECT 106.680 199.390 106.960 199.670 ;
        RECT 110.120 199.390 110.400 199.670 ;
        RECT 110.640 199.390 110.920 199.670 ;
        RECT 110.040 198.510 110.320 198.790 ;
        RECT 110.560 198.510 110.840 198.790 ;
        RECT 93.400 197.630 93.680 197.910 ;
        RECT 93.920 197.630 94.200 197.910 ;
        RECT 97.360 197.630 97.640 197.910 ;
        RECT 97.880 197.630 98.160 197.910 ;
        RECT 106.160 197.630 106.440 197.910 ;
        RECT 106.680 197.630 106.960 197.910 ;
        RECT 110.120 197.630 110.400 197.910 ;
        RECT 110.640 197.630 110.920 197.910 ;
        RECT 93.400 195.870 93.680 196.150 ;
        RECT 93.920 195.870 94.200 196.150 ;
        RECT 97.360 195.870 97.640 196.150 ;
        RECT 97.880 195.870 98.160 196.150 ;
        RECT 80.960 192.350 81.240 192.630 ;
        RECT 81.480 192.350 81.760 192.630 ;
        RECT 84.920 192.350 85.200 192.630 ;
        RECT 85.440 192.350 85.720 192.630 ;
        RECT 93.400 192.350 93.680 192.630 ;
        RECT 93.920 192.350 94.200 192.630 ;
        RECT 97.360 192.350 97.640 192.630 ;
        RECT 97.880 192.350 98.160 192.630 ;
        RECT 80.960 191.470 81.240 191.750 ;
        RECT 81.480 191.470 81.760 191.750 ;
        RECT 84.920 191.470 85.200 191.750 ;
        RECT 85.440 191.470 85.720 191.750 ;
        RECT 93.400 191.470 93.680 191.750 ;
        RECT 93.920 191.470 94.200 191.750 ;
        RECT 97.360 191.470 97.640 191.750 ;
        RECT 97.880 191.470 98.160 191.750 ;
        RECT 86.920 191.030 87.200 191.310 ;
        RECT 87.440 191.030 87.720 191.310 ;
        RECT 91.240 191.030 91.520 191.310 ;
        RECT 91.760 191.030 92.040 191.310 ;
        RECT 84.920 188.830 85.200 189.110 ;
        RECT 85.440 188.830 85.720 189.110 ;
        RECT 93.400 188.830 93.680 189.110 ;
        RECT 93.920 188.830 94.200 189.110 ;
        RECT 80.960 187.950 81.240 188.230 ;
        RECT 81.480 187.950 81.760 188.230 ;
        RECT 84.920 187.950 85.200 188.230 ;
        RECT 85.440 187.950 85.720 188.230 ;
        RECT 93.400 187.950 93.680 188.230 ;
        RECT 93.920 187.950 94.200 188.230 ;
        RECT 97.360 187.950 97.640 188.230 ;
        RECT 97.880 187.950 98.160 188.230 ;
        RECT 84.920 185.310 85.200 185.590 ;
        RECT 85.440 185.310 85.720 185.590 ;
        RECT 93.400 185.310 93.680 185.590 ;
        RECT 93.920 185.310 94.200 185.590 ;
        RECT 80.960 184.430 81.240 184.710 ;
        RECT 81.480 184.430 81.760 184.710 ;
        RECT 84.920 184.430 85.200 184.710 ;
        RECT 85.440 184.430 85.720 184.710 ;
        RECT 93.400 184.430 93.680 184.710 ;
        RECT 93.920 184.430 94.200 184.710 ;
        RECT 97.360 184.430 97.640 184.710 ;
        RECT 97.880 184.430 98.160 184.710 ;
        RECT 82.300 182.870 82.580 183.150 ;
        RECT 82.300 182.350 82.580 182.630 ;
        RECT 96.540 182.870 96.820 183.150 ;
        RECT 96.540 182.350 96.820 182.630 ;
        RECT 80.960 181.790 81.240 182.070 ;
        RECT 81.480 181.790 81.760 182.070 ;
        RECT 84.920 181.790 85.200 182.070 ;
        RECT 85.440 181.790 85.720 182.070 ;
        RECT 93.400 181.790 93.680 182.070 ;
        RECT 93.920 181.790 94.200 182.070 ;
        RECT 97.360 181.790 97.640 182.070 ;
        RECT 97.880 181.790 98.160 182.070 ;
        RECT 80.960 180.910 81.240 181.190 ;
        RECT 81.480 180.910 81.760 181.190 ;
        RECT 84.920 180.910 85.200 181.190 ;
        RECT 85.440 180.910 85.720 181.190 ;
        RECT 93.400 180.910 93.680 181.190 ;
        RECT 93.920 180.910 94.200 181.190 ;
        RECT 97.360 180.910 97.640 181.190 ;
        RECT 97.880 180.910 98.160 181.190 ;
        RECT 84.920 178.270 85.200 178.550 ;
        RECT 85.440 178.270 85.720 178.550 ;
        RECT 93.400 178.270 93.680 178.550 ;
        RECT 93.920 178.270 94.200 178.550 ;
        RECT 80.960 177.390 81.240 177.670 ;
        RECT 81.480 177.390 81.760 177.670 ;
        RECT 84.920 177.390 85.200 177.670 ;
        RECT 85.440 177.390 85.720 177.670 ;
        RECT 93.400 177.390 93.680 177.670 ;
        RECT 93.920 177.390 94.200 177.670 ;
        RECT 97.360 177.390 97.640 177.670 ;
        RECT 97.880 177.390 98.160 177.670 ;
        RECT 83.175 175.830 83.455 176.110 ;
        RECT 83.175 175.310 83.455 175.590 ;
        RECT 95.665 175.830 95.945 176.110 ;
        RECT 95.665 175.310 95.945 175.590 ;
        RECT 80.960 174.750 81.240 175.030 ;
        RECT 81.480 174.750 81.760 175.030 ;
        RECT 84.920 174.750 85.200 175.030 ;
        RECT 85.440 174.750 85.720 175.030 ;
        RECT 80.960 173.870 81.240 174.150 ;
        RECT 81.480 173.870 81.760 174.150 ;
        RECT 84.920 173.870 85.200 174.150 ;
        RECT 85.440 173.870 85.720 174.150 ;
        RECT 84.920 171.230 85.200 171.510 ;
        RECT 85.440 171.230 85.720 171.510 ;
        RECT 80.960 170.350 81.240 170.630 ;
        RECT 81.480 170.350 81.760 170.630 ;
        RECT 84.920 170.350 85.200 170.630 ;
        RECT 85.440 170.350 85.720 170.630 ;
        RECT 83.975 168.790 84.255 169.070 ;
        RECT 83.975 168.270 84.255 168.550 ;
        RECT 80.960 167.710 81.240 167.990 ;
        RECT 81.480 167.710 81.760 167.990 ;
        RECT 84.920 167.710 85.200 167.990 ;
        RECT 85.440 167.710 85.720 167.990 ;
        RECT 80.960 166.830 81.240 167.110 ;
        RECT 81.480 166.830 81.760 167.110 ;
        RECT 84.920 166.830 85.200 167.110 ;
        RECT 85.440 166.830 85.720 167.110 ;
        RECT 84.920 164.190 85.200 164.470 ;
        RECT 85.440 164.190 85.720 164.470 ;
        RECT 80.960 163.310 81.240 163.590 ;
        RECT 81.480 163.310 81.760 163.590 ;
        RECT 84.920 163.310 85.200 163.590 ;
        RECT 85.440 163.310 85.720 163.590 ;
        RECT 80.960 160.670 81.240 160.950 ;
        RECT 81.480 160.670 81.760 160.950 ;
        RECT 84.920 160.670 85.200 160.950 ;
        RECT 85.440 160.670 85.720 160.950 ;
        RECT 78.640 159.350 78.920 159.630 ;
        RECT 79.160 159.350 79.440 159.630 ;
        RECT 80.960 155.390 81.240 155.670 ;
        RECT 81.480 155.390 81.760 155.670 ;
        RECT 84.920 155.390 85.200 155.670 ;
        RECT 85.440 155.390 85.720 155.670 ;
        RECT 87.000 168.110 87.280 168.390 ;
        RECT 87.520 168.110 87.800 168.390 ;
        RECT 91.320 168.110 91.600 168.390 ;
        RECT 91.840 168.110 92.120 168.390 ;
        RECT 86.920 155.830 87.200 156.110 ;
        RECT 87.440 155.830 87.720 156.110 ;
        RECT 80.960 150.110 81.240 150.390 ;
        RECT 81.480 150.110 81.760 150.390 ;
        RECT 84.920 150.110 85.200 150.390 ;
        RECT 85.440 150.110 85.720 150.390 ;
        RECT 80.960 148.350 81.240 148.630 ;
        RECT 81.480 148.350 81.760 148.630 ;
        RECT 84.920 148.350 85.200 148.630 ;
        RECT 85.440 148.350 85.720 148.630 ;
        RECT 80.960 147.470 81.240 147.750 ;
        RECT 81.480 147.470 81.760 147.750 ;
        RECT 84.920 146.590 85.200 146.870 ;
        RECT 85.440 146.590 85.720 146.870 ;
        RECT 84.920 145.710 85.200 145.990 ;
        RECT 85.440 145.710 85.720 145.990 ;
        RECT 87.000 150.510 87.280 150.790 ;
        RECT 87.520 150.510 87.800 150.790 ;
        RECT 80.880 143.030 81.160 143.310 ;
        RECT 81.400 143.030 81.680 143.310 ;
        RECT 84.920 143.070 85.200 143.350 ;
        RECT 85.440 143.070 85.720 143.350 ;
        RECT 72.160 142.190 72.440 142.470 ;
        RECT 72.680 142.190 72.960 142.470 ;
        RECT 80.960 142.190 81.240 142.470 ;
        RECT 81.480 142.190 81.760 142.470 ;
        RECT 66.120 141.710 66.400 141.990 ;
        RECT 66.640 141.710 66.920 141.990 ;
        RECT 87.000 141.710 87.280 141.990 ;
        RECT 87.520 141.710 87.800 141.990 ;
        RECT 91.240 155.830 91.520 156.110 ;
        RECT 91.760 155.830 92.040 156.110 ;
        RECT 93.400 174.750 93.680 175.030 ;
        RECT 93.920 174.750 94.200 175.030 ;
        RECT 97.360 174.750 97.640 175.030 ;
        RECT 97.880 174.750 98.160 175.030 ;
        RECT 93.400 173.870 93.680 174.150 ;
        RECT 93.920 173.870 94.200 174.150 ;
        RECT 97.360 173.870 97.640 174.150 ;
        RECT 97.880 173.870 98.160 174.150 ;
        RECT 93.400 171.230 93.680 171.510 ;
        RECT 93.920 171.230 94.200 171.510 ;
        RECT 93.400 170.350 93.680 170.630 ;
        RECT 93.920 170.350 94.200 170.630 ;
        RECT 97.360 170.350 97.640 170.630 ;
        RECT 97.880 170.350 98.160 170.630 ;
        RECT 94.865 168.790 95.145 169.070 ;
        RECT 94.865 168.270 95.145 168.550 ;
        RECT 93.400 167.710 93.680 167.990 ;
        RECT 93.920 167.710 94.200 167.990 ;
        RECT 97.360 167.710 97.640 167.990 ;
        RECT 97.880 167.710 98.160 167.990 ;
        RECT 93.400 166.830 93.680 167.110 ;
        RECT 93.920 166.830 94.200 167.110 ;
        RECT 97.360 166.830 97.640 167.110 ;
        RECT 97.880 166.830 98.160 167.110 ;
        RECT 93.400 164.190 93.680 164.470 ;
        RECT 93.920 164.190 94.200 164.470 ;
        RECT 93.400 163.310 93.680 163.590 ;
        RECT 93.920 163.310 94.200 163.590 ;
        RECT 97.360 163.310 97.640 163.590 ;
        RECT 97.880 163.310 98.160 163.590 ;
        RECT 93.400 160.670 93.680 160.950 ;
        RECT 93.920 160.670 94.200 160.950 ;
        RECT 97.360 160.670 97.640 160.950 ;
        RECT 97.880 160.670 98.160 160.950 ;
        RECT 99.520 159.350 99.800 159.630 ;
        RECT 100.040 159.350 100.320 159.630 ;
        RECT 93.400 155.390 93.680 155.670 ;
        RECT 93.920 155.390 94.200 155.670 ;
        RECT 97.360 155.390 97.640 155.670 ;
        RECT 97.880 155.390 98.160 155.670 ;
        RECT 91.320 150.510 91.600 150.790 ;
        RECT 91.840 150.510 92.120 150.790 ;
        RECT 93.400 150.110 93.680 150.390 ;
        RECT 93.920 150.110 94.200 150.390 ;
        RECT 97.360 150.110 97.640 150.390 ;
        RECT 97.880 150.110 98.160 150.390 ;
        RECT 93.400 148.350 93.680 148.630 ;
        RECT 93.920 148.350 94.200 148.630 ;
        RECT 97.360 148.350 97.640 148.630 ;
        RECT 97.880 148.350 98.160 148.630 ;
        RECT 97.360 147.470 97.640 147.750 ;
        RECT 97.880 147.470 98.160 147.750 ;
        RECT 93.400 146.590 93.680 146.870 ;
        RECT 93.920 146.590 94.200 146.870 ;
        RECT 93.400 145.710 93.680 145.990 ;
        RECT 93.920 145.710 94.200 145.990 ;
        RECT 93.400 143.070 93.680 143.350 ;
        RECT 93.920 143.070 94.200 143.350 ;
        RECT 97.440 143.030 97.720 143.310 ;
        RECT 97.960 143.030 98.240 143.310 ;
        RECT 106.160 195.870 106.440 196.150 ;
        RECT 106.680 195.870 106.960 196.150 ;
        RECT 110.120 195.870 110.400 196.150 ;
        RECT 110.640 195.870 110.920 196.150 ;
        RECT 118.600 199.390 118.880 199.670 ;
        RECT 119.120 199.390 119.400 199.670 ;
        RECT 122.560 199.390 122.840 199.670 ;
        RECT 123.080 199.390 123.360 199.670 ;
        RECT 143.740 214.180 144.020 214.460 ;
        RECT 144.260 214.180 144.540 214.460 ;
        RECT 147.700 215.940 147.980 216.220 ;
        RECT 148.220 215.940 148.500 216.220 ;
        RECT 147.700 215.060 147.980 215.340 ;
        RECT 148.220 215.060 148.500 215.340 ;
        RECT 149.860 212.860 150.140 213.140 ;
        RECT 150.380 212.860 150.660 213.140 ;
        RECT 143.740 210.660 144.020 210.940 ;
        RECT 144.260 210.660 144.540 210.940 ;
        RECT 147.700 210.660 147.980 210.940 ;
        RECT 148.220 210.660 148.500 210.940 ;
        RECT 143.740 208.900 144.020 209.180 ;
        RECT 144.260 208.900 144.540 209.180 ;
        RECT 147.700 208.900 147.980 209.180 ;
        RECT 148.220 208.900 148.500 209.180 ;
        RECT 143.740 205.380 144.020 205.660 ;
        RECT 144.260 205.380 144.540 205.660 ;
        RECT 147.700 205.380 147.980 205.660 ;
        RECT 148.220 205.380 148.500 205.660 ;
        RECT 143.740 201.860 144.020 202.140 ;
        RECT 144.260 201.860 144.540 202.140 ;
        RECT 147.700 201.860 147.980 202.140 ;
        RECT 148.220 201.860 148.500 202.140 ;
        RECT 143.740 200.100 144.020 200.380 ;
        RECT 144.260 200.100 144.540 200.380 ;
        RECT 147.700 200.100 147.980 200.380 ;
        RECT 148.220 200.100 148.500 200.380 ;
        RECT 147.700 199.220 147.980 199.500 ;
        RECT 148.220 199.220 148.500 199.500 ;
        RECT 112.120 194.550 112.400 194.830 ;
        RECT 112.640 194.550 112.920 194.830 ;
        RECT 106.160 192.350 106.440 192.630 ;
        RECT 106.680 192.350 106.960 192.630 ;
        RECT 110.120 192.350 110.400 192.630 ;
        RECT 110.640 192.350 110.920 192.630 ;
        RECT 106.160 191.470 106.440 191.750 ;
        RECT 106.680 191.470 106.960 191.750 ;
        RECT 110.120 191.470 110.400 191.750 ;
        RECT 110.640 191.470 110.920 191.750 ;
        RECT 112.120 191.030 112.400 191.310 ;
        RECT 112.640 191.030 112.920 191.310 ;
        RECT 110.120 188.830 110.400 189.110 ;
        RECT 110.640 188.830 110.920 189.110 ;
        RECT 106.160 187.950 106.440 188.230 ;
        RECT 106.680 187.950 106.960 188.230 ;
        RECT 110.120 187.950 110.400 188.230 ;
        RECT 110.640 187.950 110.920 188.230 ;
        RECT 118.600 197.630 118.880 197.910 ;
        RECT 119.120 197.630 119.400 197.910 ;
        RECT 122.560 197.630 122.840 197.910 ;
        RECT 123.080 197.630 123.360 197.910 ;
        RECT 143.740 196.580 144.020 196.860 ;
        RECT 144.260 196.580 144.540 196.860 ;
        RECT 147.700 196.580 147.980 196.860 ;
        RECT 148.220 196.580 148.500 196.860 ;
        RECT 143.740 194.820 144.020 195.100 ;
        RECT 144.260 194.820 144.540 195.100 ;
        RECT 147.700 194.820 147.980 195.100 ;
        RECT 148.220 194.820 148.500 195.100 ;
        RECT 141.580 193.500 141.860 193.780 ;
        RECT 142.100 193.500 142.380 193.780 ;
        RECT 110.120 185.310 110.400 185.590 ;
        RECT 110.640 185.310 110.920 185.590 ;
        RECT 106.160 184.430 106.440 184.710 ;
        RECT 106.680 184.430 106.960 184.710 ;
        RECT 110.120 184.430 110.400 184.710 ;
        RECT 110.640 184.430 110.920 184.710 ;
        RECT 107.500 182.870 107.780 183.150 ;
        RECT 107.500 182.350 107.780 182.630 ;
        RECT 106.160 181.790 106.440 182.070 ;
        RECT 106.680 181.790 106.960 182.070 ;
        RECT 110.120 181.790 110.400 182.070 ;
        RECT 110.640 181.790 110.920 182.070 ;
        RECT 106.160 180.910 106.440 181.190 ;
        RECT 106.680 180.910 106.960 181.190 ;
        RECT 110.120 180.910 110.400 181.190 ;
        RECT 110.640 180.910 110.920 181.190 ;
        RECT 110.120 178.270 110.400 178.550 ;
        RECT 110.640 178.270 110.920 178.550 ;
        RECT 106.160 177.390 106.440 177.670 ;
        RECT 106.680 177.390 106.960 177.670 ;
        RECT 110.120 177.390 110.400 177.670 ;
        RECT 110.640 177.390 110.920 177.670 ;
        RECT 108.375 175.830 108.655 176.110 ;
        RECT 108.375 175.310 108.655 175.590 ;
        RECT 106.160 174.750 106.440 175.030 ;
        RECT 106.680 174.750 106.960 175.030 ;
        RECT 110.120 174.750 110.400 175.030 ;
        RECT 110.640 174.750 110.920 175.030 ;
        RECT 106.160 173.870 106.440 174.150 ;
        RECT 106.680 173.870 106.960 174.150 ;
        RECT 110.120 173.870 110.400 174.150 ;
        RECT 110.640 173.870 110.920 174.150 ;
        RECT 110.120 171.230 110.400 171.510 ;
        RECT 110.640 171.230 110.920 171.510 ;
        RECT 106.160 170.350 106.440 170.630 ;
        RECT 106.680 170.350 106.960 170.630 ;
        RECT 110.120 170.350 110.400 170.630 ;
        RECT 110.640 170.350 110.920 170.630 ;
        RECT 109.175 168.790 109.455 169.070 ;
        RECT 109.175 168.270 109.455 168.550 ;
        RECT 106.160 167.710 106.440 167.990 ;
        RECT 106.680 167.710 106.960 167.990 ;
        RECT 110.120 167.710 110.400 167.990 ;
        RECT 110.640 167.710 110.920 167.990 ;
        RECT 106.160 166.830 106.440 167.110 ;
        RECT 106.680 166.830 106.960 167.110 ;
        RECT 110.120 166.830 110.400 167.110 ;
        RECT 110.640 166.830 110.920 167.110 ;
        RECT 110.120 164.190 110.400 164.470 ;
        RECT 110.640 164.190 110.920 164.470 ;
        RECT 106.160 163.310 106.440 163.590 ;
        RECT 106.680 163.310 106.960 163.590 ;
        RECT 110.120 163.310 110.400 163.590 ;
        RECT 110.640 163.310 110.920 163.590 ;
        RECT 106.160 160.670 106.440 160.950 ;
        RECT 106.680 160.670 106.960 160.950 ;
        RECT 110.120 160.670 110.400 160.950 ;
        RECT 110.640 160.670 110.920 160.950 ;
        RECT 103.840 159.350 104.120 159.630 ;
        RECT 104.360 159.350 104.640 159.630 ;
        RECT 106.160 155.390 106.440 155.670 ;
        RECT 106.680 155.390 106.960 155.670 ;
        RECT 110.120 155.390 110.400 155.670 ;
        RECT 110.640 155.390 110.920 155.670 ;
        RECT 112.200 168.110 112.480 168.390 ;
        RECT 112.720 168.110 113.000 168.390 ;
        RECT 112.120 155.830 112.400 156.110 ;
        RECT 112.640 155.830 112.920 156.110 ;
        RECT 106.160 150.110 106.440 150.390 ;
        RECT 106.680 150.110 106.960 150.390 ;
        RECT 110.120 150.110 110.400 150.390 ;
        RECT 110.640 150.110 110.920 150.390 ;
        RECT 106.160 148.350 106.440 148.630 ;
        RECT 106.680 148.350 106.960 148.630 ;
        RECT 110.120 148.350 110.400 148.630 ;
        RECT 110.640 148.350 110.920 148.630 ;
        RECT 106.160 147.470 106.440 147.750 ;
        RECT 106.680 147.470 106.960 147.750 ;
        RECT 110.120 146.590 110.400 146.870 ;
        RECT 110.640 146.590 110.920 146.870 ;
        RECT 110.120 145.710 110.400 145.990 ;
        RECT 110.640 145.710 110.920 145.990 ;
        RECT 112.200 150.510 112.480 150.790 ;
        RECT 112.720 150.510 113.000 150.790 ;
        RECT 106.080 143.030 106.360 143.310 ;
        RECT 106.600 143.030 106.880 143.310 ;
        RECT 110.120 143.070 110.400 143.350 ;
        RECT 110.640 143.070 110.920 143.350 ;
        RECT 97.360 142.190 97.640 142.470 ;
        RECT 97.880 142.190 98.160 142.470 ;
        RECT 106.160 142.190 106.440 142.470 ;
        RECT 106.680 142.190 106.960 142.470 ;
        RECT 91.320 141.710 91.600 141.990 ;
        RECT 91.840 141.710 92.120 141.990 ;
        RECT 112.200 141.710 112.480 141.990 ;
        RECT 112.720 141.710 113.000 141.990 ;
        RECT 116.440 182.230 116.720 182.510 ;
        RECT 116.960 182.230 117.240 182.510 ;
        RECT 122.560 186.190 122.840 186.470 ;
        RECT 123.080 186.190 123.360 186.470 ;
        RECT 118.600 185.310 118.880 185.590 ;
        RECT 119.120 185.310 119.400 185.590 ;
        RECT 122.560 184.430 122.840 184.710 ;
        RECT 123.080 184.430 123.360 184.710 ;
        RECT 122.560 181.790 122.840 182.070 ;
        RECT 123.080 181.790 123.360 182.070 ;
        RECT 122.560 180.910 122.840 181.190 ;
        RECT 123.080 180.910 123.360 181.190 ;
        RECT 122.560 178.270 122.840 178.550 ;
        RECT 123.080 178.270 123.360 178.550 ;
        RECT 122.560 177.390 122.840 177.670 ;
        RECT 123.080 177.390 123.360 177.670 ;
        RECT 122.560 174.750 122.840 175.030 ;
        RECT 123.080 174.750 123.360 175.030 ;
        RECT 122.560 173.870 122.840 174.150 ;
        RECT 123.080 173.870 123.360 174.150 ;
        RECT 118.600 172.990 118.880 173.270 ;
        RECT 119.120 172.990 119.400 173.270 ;
        RECT 118.600 172.110 118.880 172.390 ;
        RECT 119.120 172.110 119.400 172.390 ;
        RECT 122.560 172.110 122.840 172.390 ;
        RECT 123.080 172.110 123.360 172.390 ;
        RECT 122.560 170.350 122.840 170.630 ;
        RECT 123.080 170.350 123.360 170.630 ;
        RECT 118.600 169.470 118.880 169.750 ;
        RECT 119.120 169.470 119.400 169.750 ;
        RECT 122.560 169.470 122.840 169.750 ;
        RECT 123.080 169.470 123.360 169.750 ;
        RECT 118.600 168.590 118.880 168.870 ;
        RECT 119.120 168.590 119.400 168.870 ;
        RECT 122.560 168.590 122.840 168.870 ;
        RECT 123.080 168.590 123.360 168.870 ;
        RECT 118.680 167.020 118.960 167.300 ;
        RECT 119.200 167.020 119.480 167.300 ;
        RECT 124.720 176.950 125.000 177.230 ;
        RECT 125.240 176.950 125.520 177.230 ;
        RECT 143.740 189.540 144.020 189.820 ;
        RECT 144.260 189.540 144.540 189.820 ;
        RECT 147.700 191.300 147.980 191.580 ;
        RECT 148.220 191.300 148.500 191.580 ;
        RECT 147.700 190.420 147.980 190.700 ;
        RECT 148.220 190.420 148.500 190.700 ;
        RECT 149.860 188.220 150.140 188.500 ;
        RECT 150.380 188.220 150.660 188.500 ;
        RECT 143.740 186.020 144.020 186.300 ;
        RECT 144.260 186.020 144.540 186.300 ;
        RECT 147.700 186.020 147.980 186.300 ;
        RECT 148.220 186.020 148.500 186.300 ;
        RECT 143.740 184.260 144.020 184.540 ;
        RECT 144.260 184.260 144.540 184.540 ;
        RECT 147.700 184.260 147.980 184.540 ;
        RECT 148.220 184.260 148.500 184.540 ;
        RECT 143.740 180.740 144.020 181.020 ;
        RECT 144.260 180.740 144.540 181.020 ;
        RECT 147.700 180.740 147.980 181.020 ;
        RECT 148.220 180.740 148.500 181.020 ;
        RECT 143.740 177.220 144.020 177.500 ;
        RECT 144.260 177.220 144.540 177.500 ;
        RECT 147.700 177.220 147.980 177.500 ;
        RECT 148.220 177.220 148.500 177.500 ;
        RECT 143.740 175.460 144.020 175.740 ;
        RECT 144.260 175.460 144.540 175.740 ;
        RECT 147.700 175.460 147.980 175.740 ;
        RECT 148.220 175.460 148.500 175.740 ;
        RECT 147.700 174.580 147.980 174.860 ;
        RECT 148.220 174.580 148.500 174.860 ;
        RECT 143.740 171.940 144.020 172.220 ;
        RECT 144.260 171.940 144.540 172.220 ;
        RECT 147.700 171.940 147.980 172.220 ;
        RECT 148.220 171.940 148.500 172.220 ;
        RECT 143.740 170.180 144.020 170.460 ;
        RECT 144.260 170.180 144.540 170.460 ;
        RECT 147.700 170.180 147.980 170.460 ;
        RECT 148.220 170.180 148.500 170.460 ;
        RECT 141.580 168.860 141.860 169.140 ;
        RECT 142.100 168.860 142.380 169.140 ;
        RECT 118.600 165.950 118.880 166.230 ;
        RECT 119.120 165.950 119.400 166.230 ;
        RECT 122.560 165.950 122.840 166.230 ;
        RECT 123.080 165.950 123.360 166.230 ;
        RECT 122.560 165.070 122.840 165.350 ;
        RECT 123.080 165.070 123.360 165.350 ;
        RECT 122.560 162.430 122.840 162.710 ;
        RECT 123.080 162.430 123.360 162.710 ;
        RECT 122.560 161.550 122.840 161.830 ;
        RECT 123.080 161.550 123.360 161.830 ;
        RECT 122.560 158.910 122.840 159.190 ;
        RECT 123.080 158.910 123.360 159.190 ;
        RECT 122.560 158.030 122.840 158.310 ;
        RECT 123.080 158.030 123.360 158.310 ;
        RECT 124.720 157.590 125.000 157.870 ;
        RECT 125.240 157.590 125.520 157.870 ;
        RECT 116.440 150.550 116.720 150.830 ;
        RECT 116.960 150.550 117.240 150.830 ;
        RECT 122.560 155.390 122.840 155.670 ;
        RECT 123.080 155.390 123.360 155.670 ;
        RECT 122.560 154.510 122.840 154.790 ;
        RECT 123.080 154.510 123.360 154.790 ;
        RECT 118.600 153.630 118.880 153.910 ;
        RECT 119.120 153.630 119.400 153.910 ;
        RECT 143.740 164.900 144.020 165.180 ;
        RECT 144.260 164.900 144.540 165.180 ;
        RECT 147.700 166.660 147.980 166.940 ;
        RECT 148.220 166.660 148.500 166.940 ;
        RECT 147.700 165.780 147.980 166.060 ;
        RECT 148.220 165.780 148.500 166.060 ;
        RECT 149.860 163.580 150.140 163.860 ;
        RECT 150.380 163.580 150.660 163.860 ;
        RECT 143.740 161.380 144.020 161.660 ;
        RECT 144.260 161.380 144.540 161.660 ;
        RECT 147.700 161.380 147.980 161.660 ;
        RECT 148.220 161.380 148.500 161.660 ;
        RECT 143.740 159.620 144.020 159.900 ;
        RECT 144.260 159.620 144.540 159.900 ;
        RECT 147.700 159.620 147.980 159.900 ;
        RECT 148.220 159.620 148.500 159.900 ;
        RECT 143.740 156.100 144.020 156.380 ;
        RECT 144.260 156.100 144.540 156.380 ;
        RECT 147.700 156.100 147.980 156.380 ;
        RECT 148.220 156.100 148.500 156.380 ;
        RECT 143.740 152.580 144.020 152.860 ;
        RECT 144.260 152.580 144.540 152.860 ;
        RECT 147.700 152.580 147.980 152.860 ;
        RECT 148.220 152.580 148.500 152.860 ;
        RECT 143.740 150.820 144.020 151.100 ;
        RECT 144.260 150.820 144.540 151.100 ;
        RECT 147.700 150.820 147.980 151.100 ;
        RECT 148.220 150.820 148.500 151.100 ;
        RECT 147.700 149.940 147.980 150.220 ;
        RECT 148.220 149.940 148.500 150.220 ;
        RECT 143.740 147.300 144.020 147.580 ;
        RECT 144.260 147.300 144.540 147.580 ;
        RECT 147.700 147.300 147.980 147.580 ;
        RECT 148.220 147.300 148.500 147.580 ;
        RECT 143.740 145.540 144.020 145.820 ;
        RECT 144.260 145.540 144.540 145.820 ;
        RECT 147.700 145.540 147.980 145.820 ;
        RECT 148.220 145.540 148.500 145.820 ;
        RECT 141.580 144.220 141.860 144.500 ;
        RECT 142.100 144.220 142.380 144.500 ;
        RECT 122.560 142.190 122.840 142.470 ;
        RECT 123.080 142.190 123.360 142.470 ;
        RECT 118.600 141.310 118.880 141.590 ;
        RECT 119.120 141.310 119.400 141.590 ;
        RECT 17.800 140.430 18.080 140.710 ;
        RECT 18.320 140.430 18.600 140.710 ;
        RECT 21.760 140.430 22.040 140.710 ;
        RECT 22.280 140.430 22.560 140.710 ;
        RECT 30.560 140.430 30.840 140.710 ;
        RECT 31.080 140.430 31.360 140.710 ;
        RECT 34.520 140.430 34.800 140.710 ;
        RECT 35.040 140.430 35.320 140.710 ;
        RECT 43.000 140.430 43.280 140.710 ;
        RECT 43.520 140.430 43.800 140.710 ;
        RECT 46.960 140.430 47.240 140.710 ;
        RECT 47.480 140.430 47.760 140.710 ;
        RECT 55.760 140.430 56.040 140.710 ;
        RECT 56.280 140.430 56.560 140.710 ;
        RECT 59.720 140.430 60.000 140.710 ;
        RECT 60.240 140.430 60.520 140.710 ;
        RECT 68.200 140.430 68.480 140.710 ;
        RECT 68.720 140.430 69.000 140.710 ;
        RECT 72.160 140.430 72.440 140.710 ;
        RECT 72.680 140.430 72.960 140.710 ;
        RECT 80.960 140.430 81.240 140.710 ;
        RECT 81.480 140.430 81.760 140.710 ;
        RECT 84.920 140.430 85.200 140.710 ;
        RECT 85.440 140.430 85.720 140.710 ;
        RECT 93.400 140.430 93.680 140.710 ;
        RECT 93.920 140.430 94.200 140.710 ;
        RECT 97.360 140.430 97.640 140.710 ;
        RECT 97.880 140.430 98.160 140.710 ;
        RECT 106.160 140.430 106.440 140.710 ;
        RECT 106.680 140.430 106.960 140.710 ;
        RECT 110.120 140.430 110.400 140.710 ;
        RECT 110.640 140.430 110.920 140.710 ;
        RECT 118.600 140.430 118.880 140.710 ;
        RECT 119.120 140.430 119.400 140.710 ;
        RECT 122.560 140.430 122.840 140.710 ;
        RECT 123.080 140.430 123.360 140.710 ;
        RECT 17.800 139.550 18.080 139.830 ;
        RECT 18.320 139.550 18.600 139.830 ;
        RECT 21.760 139.550 22.040 139.830 ;
        RECT 22.280 139.550 22.560 139.830 ;
        RECT 30.560 139.550 30.840 139.830 ;
        RECT 31.080 139.550 31.360 139.830 ;
        RECT 34.520 139.550 34.800 139.830 ;
        RECT 35.040 139.550 35.320 139.830 ;
        RECT 43.000 139.550 43.280 139.830 ;
        RECT 43.520 139.550 43.800 139.830 ;
        RECT 46.960 139.550 47.240 139.830 ;
        RECT 47.480 139.550 47.760 139.830 ;
        RECT 55.760 139.550 56.040 139.830 ;
        RECT 56.280 139.550 56.560 139.830 ;
        RECT 59.720 139.550 60.000 139.830 ;
        RECT 60.240 139.550 60.520 139.830 ;
        RECT 68.200 139.550 68.480 139.830 ;
        RECT 68.720 139.550 69.000 139.830 ;
        RECT 72.160 139.550 72.440 139.830 ;
        RECT 72.680 139.550 72.960 139.830 ;
        RECT 80.960 139.550 81.240 139.830 ;
        RECT 81.480 139.550 81.760 139.830 ;
        RECT 84.920 139.550 85.200 139.830 ;
        RECT 85.440 139.550 85.720 139.830 ;
        RECT 93.400 139.550 93.680 139.830 ;
        RECT 93.920 139.550 94.200 139.830 ;
        RECT 97.360 139.550 97.640 139.830 ;
        RECT 97.880 139.550 98.160 139.830 ;
        RECT 106.160 139.550 106.440 139.830 ;
        RECT 106.680 139.550 106.960 139.830 ;
        RECT 110.120 139.550 110.400 139.830 ;
        RECT 110.640 139.550 110.920 139.830 ;
        RECT 118.600 139.550 118.880 139.830 ;
        RECT 119.120 139.550 119.400 139.830 ;
        RECT 122.560 139.550 122.840 139.830 ;
        RECT 123.080 139.550 123.360 139.830 ;
        RECT 72.050 135.620 72.330 135.900 ;
        RECT 72.050 135.100 72.330 135.380 ;
        RECT 65.150 128.830 65.430 129.110 ;
        RECT 65.150 128.310 65.430 128.590 ;
        RECT 63.350 127.860 63.630 128.140 ;
        RECT 63.350 127.340 63.630 127.620 ;
        RECT 61.550 126.890 61.830 127.170 ;
        RECT 61.550 126.370 61.830 126.650 ;
        RECT 60.650 120.100 60.930 120.380 ;
        RECT 60.650 119.580 60.930 119.860 ;
        RECT 12.310 101.240 12.590 101.520 ;
        RECT 12.310 100.720 12.590 101.000 ;
        RECT 13.710 97.150 13.990 97.430 ;
        RECT 13.710 96.630 13.990 96.910 ;
        RECT 15.110 97.150 15.390 97.430 ;
        RECT 15.110 96.630 15.390 96.910 ;
        RECT 16.510 97.150 16.790 97.430 ;
        RECT 16.510 96.630 16.790 96.910 ;
        RECT 17.910 97.150 18.190 97.430 ;
        RECT 17.910 96.630 18.190 96.910 ;
        RECT 19.310 103.270 19.590 103.550 ;
        RECT 19.310 102.750 19.590 103.030 ;
        RECT 20.710 103.270 20.990 103.550 ;
        RECT 20.710 102.750 20.990 103.030 ;
        RECT 22.110 106.330 22.390 106.610 ;
        RECT 22.110 105.810 22.390 106.090 ;
        RECT 23.510 109.390 23.790 109.670 ;
        RECT 23.510 108.870 23.790 109.150 ;
        RECT 24.910 100.210 25.190 100.490 ;
        RECT 24.910 99.690 25.190 99.970 ;
        RECT 26.310 106.330 26.590 106.610 ;
        RECT 26.310 105.810 26.590 106.090 ;
        RECT 27.710 103.270 27.990 103.550 ;
        RECT 27.710 102.750 27.990 103.030 ;
        RECT 29.110 103.270 29.390 103.550 ;
        RECT 29.110 102.750 29.390 103.030 ;
        RECT 30.510 97.150 30.790 97.430 ;
        RECT 30.510 96.630 30.790 96.910 ;
        RECT 31.910 97.150 32.190 97.430 ;
        RECT 31.910 96.630 32.190 96.910 ;
        RECT 33.310 97.150 33.590 97.430 ;
        RECT 33.310 96.630 33.590 96.910 ;
        RECT 34.710 97.150 34.990 97.430 ;
        RECT 34.710 96.630 34.990 96.910 ;
        RECT 36.110 97.150 36.390 97.430 ;
        RECT 36.110 96.630 36.390 96.910 ;
        RECT 37.510 97.150 37.790 97.430 ;
        RECT 37.510 96.630 37.790 96.910 ;
        RECT 38.910 97.150 39.190 97.430 ;
        RECT 38.910 96.630 39.190 96.910 ;
        RECT 40.310 97.150 40.590 97.430 ;
        RECT 40.310 96.630 40.590 96.910 ;
        RECT 41.710 103.270 41.990 103.550 ;
        RECT 41.710 102.750 41.990 103.030 ;
        RECT 43.110 103.270 43.390 103.550 ;
        RECT 43.110 102.750 43.390 103.030 ;
        RECT 44.510 106.330 44.790 106.610 ;
        RECT 44.510 105.810 44.790 106.090 ;
        RECT 45.910 100.210 46.190 100.490 ;
        RECT 45.910 99.690 46.190 99.970 ;
        RECT 47.310 94.090 47.590 94.370 ;
        RECT 47.310 93.570 47.590 93.850 ;
        RECT 48.710 106.330 48.990 106.610 ;
        RECT 48.710 105.810 48.990 106.090 ;
        RECT 50.110 103.270 50.390 103.550 ;
        RECT 50.110 102.750 50.390 103.030 ;
        RECT 51.510 103.270 51.790 103.550 ;
        RECT 51.510 102.750 51.790 103.030 ;
        RECT 52.910 97.150 53.190 97.430 ;
        RECT 52.910 96.630 53.190 96.910 ;
        RECT 54.310 97.150 54.590 97.430 ;
        RECT 54.310 96.630 54.590 96.910 ;
        RECT 55.710 97.150 55.990 97.430 ;
        RECT 55.710 96.630 55.990 96.910 ;
        RECT 57.110 97.150 57.390 97.430 ;
        RECT 57.110 96.630 57.390 96.910 ;
        RECT 62.450 121.070 62.730 121.350 ;
        RECT 62.450 120.550 62.730 120.830 ;
        RECT 64.250 122.040 64.530 122.320 ;
        RECT 64.250 121.520 64.530 121.800 ;
        RECT 68.750 125.920 69.030 126.200 ;
        RECT 68.750 125.400 69.030 125.680 ;
        RECT 67.850 124.950 68.130 125.230 ;
        RECT 67.850 124.430 68.130 124.710 ;
        RECT 66.950 123.980 67.230 124.260 ;
        RECT 66.950 123.460 67.230 123.740 ;
        RECT 66.050 123.010 66.330 123.290 ;
        RECT 66.050 122.490 66.330 122.770 ;
        RECT 72.950 134.650 73.230 134.930 ;
        RECT 72.950 134.130 73.230 134.410 ;
        RECT 73.850 133.680 74.130 133.960 ;
        RECT 73.850 133.160 74.130 133.440 ;
        RECT 74.750 132.710 75.030 132.990 ;
        RECT 74.750 132.190 75.030 132.470 ;
        RECT 75.650 131.740 75.930 132.020 ;
        RECT 75.650 131.220 75.930 131.500 ;
        RECT 77.450 130.770 77.730 131.050 ;
        RECT 77.450 130.250 77.730 130.530 ;
        RECT 76.550 119.130 76.830 119.410 ;
        RECT 76.550 118.610 76.830 118.890 ;
        RECT 79.250 129.800 79.530 130.080 ;
        RECT 79.250 129.280 79.530 129.560 ;
        RECT 78.350 118.160 78.630 118.440 ;
        RECT 78.350 117.640 78.630 117.920 ;
        RECT 143.740 140.260 144.020 140.540 ;
        RECT 144.260 140.260 144.540 140.540 ;
        RECT 147.700 142.020 147.980 142.300 ;
        RECT 148.220 142.020 148.500 142.300 ;
        RECT 147.700 141.140 147.980 141.420 ;
        RECT 148.220 141.140 148.500 141.420 ;
        RECT 149.860 138.940 150.140 139.220 ;
        RECT 150.380 138.940 150.660 139.220 ;
        RECT 143.740 136.740 144.020 137.020 ;
        RECT 144.260 136.740 144.540 137.020 ;
        RECT 147.700 136.740 147.980 137.020 ;
        RECT 148.220 136.740 148.500 137.020 ;
        RECT 143.740 134.980 144.020 135.260 ;
        RECT 144.260 134.980 144.540 135.260 ;
        RECT 147.700 134.980 147.980 135.260 ;
        RECT 148.220 134.980 148.500 135.260 ;
        RECT 143.740 131.460 144.020 131.740 ;
        RECT 144.260 131.460 144.540 131.740 ;
        RECT 147.700 131.460 147.980 131.740 ;
        RECT 148.220 131.460 148.500 131.740 ;
        RECT 143.740 127.940 144.020 128.220 ;
        RECT 144.260 127.940 144.540 128.220 ;
        RECT 147.700 127.940 147.980 128.220 ;
        RECT 148.220 127.940 148.500 128.220 ;
        RECT 143.740 126.180 144.020 126.460 ;
        RECT 144.260 126.180 144.540 126.460 ;
        RECT 147.700 126.180 147.980 126.460 ;
        RECT 148.220 126.180 148.500 126.460 ;
        RECT 147.700 125.300 147.980 125.580 ;
        RECT 148.220 125.300 148.500 125.580 ;
        RECT 143.740 122.660 144.020 122.940 ;
        RECT 144.260 122.660 144.540 122.940 ;
        RECT 147.700 122.660 147.980 122.940 ;
        RECT 148.220 122.660 148.500 122.940 ;
        RECT 143.740 120.900 144.020 121.180 ;
        RECT 144.260 120.900 144.540 121.180 ;
        RECT 147.700 120.900 147.980 121.180 ;
        RECT 148.220 120.900 148.500 121.180 ;
        RECT 141.580 119.580 141.860 119.860 ;
        RECT 142.100 119.580 142.380 119.860 ;
        RECT 80.150 117.190 80.430 117.470 ;
        RECT 80.150 116.670 80.430 116.950 ;
        RECT 58.900 109.150 59.180 109.430 ;
        RECT 59.420 109.150 59.700 109.430 ;
        RECT 60.690 109.390 60.970 109.670 ;
        RECT 60.690 108.870 60.970 109.150 ;
        RECT 58.900 106.090 59.180 106.370 ;
        RECT 59.420 106.090 59.700 106.370 ;
        RECT 60.690 106.330 60.970 106.610 ;
        RECT 60.690 105.810 60.970 106.090 ;
        RECT 58.900 103.030 59.180 103.310 ;
        RECT 59.420 103.030 59.700 103.310 ;
        RECT 60.690 103.270 60.970 103.550 ;
        RECT 60.690 102.750 60.970 103.030 ;
        RECT 58.900 99.970 59.180 100.250 ;
        RECT 59.420 99.970 59.700 100.250 ;
        RECT 60.690 100.210 60.970 100.490 ;
        RECT 60.690 99.690 60.970 99.970 ;
        RECT 58.900 96.910 59.180 97.190 ;
        RECT 59.420 96.910 59.700 97.190 ;
        RECT 60.690 97.150 60.970 97.430 ;
        RECT 60.690 96.630 60.970 96.910 ;
        RECT 58.900 93.850 59.180 94.130 ;
        RECT 59.420 93.850 59.700 94.130 ;
        RECT 60.690 94.090 60.970 94.370 ;
        RECT 60.690 93.570 60.970 93.850 ;
        RECT 12.310 83.840 12.590 84.120 ;
        RECT 12.310 83.320 12.590 83.600 ;
        RECT 13.710 79.750 13.990 80.030 ;
        RECT 13.710 79.230 13.990 79.510 ;
        RECT 15.110 79.750 15.390 80.030 ;
        RECT 15.110 79.230 15.390 79.510 ;
        RECT 16.510 79.750 16.790 80.030 ;
        RECT 16.510 79.230 16.790 79.510 ;
        RECT 17.910 79.750 18.190 80.030 ;
        RECT 17.910 79.230 18.190 79.510 ;
        RECT 19.310 85.870 19.590 86.150 ;
        RECT 19.310 85.350 19.590 85.630 ;
        RECT 20.710 85.870 20.990 86.150 ;
        RECT 20.710 85.350 20.990 85.630 ;
        RECT 22.110 88.930 22.390 89.210 ;
        RECT 22.110 88.410 22.390 88.690 ;
        RECT 23.510 91.990 23.790 92.270 ;
        RECT 23.510 91.470 23.790 91.750 ;
        RECT 24.910 82.810 25.190 83.090 ;
        RECT 24.910 82.290 25.190 82.570 ;
        RECT 26.310 88.930 26.590 89.210 ;
        RECT 26.310 88.410 26.590 88.690 ;
        RECT 27.710 85.870 27.990 86.150 ;
        RECT 27.710 85.350 27.990 85.630 ;
        RECT 29.110 85.870 29.390 86.150 ;
        RECT 29.110 85.350 29.390 85.630 ;
        RECT 30.510 79.750 30.790 80.030 ;
        RECT 30.510 79.230 30.790 79.510 ;
        RECT 31.910 79.750 32.190 80.030 ;
        RECT 31.910 79.230 32.190 79.510 ;
        RECT 33.310 79.750 33.590 80.030 ;
        RECT 33.310 79.230 33.590 79.510 ;
        RECT 34.710 79.750 34.990 80.030 ;
        RECT 34.710 79.230 34.990 79.510 ;
        RECT 36.110 79.750 36.390 80.030 ;
        RECT 36.110 79.230 36.390 79.510 ;
        RECT 37.510 79.750 37.790 80.030 ;
        RECT 37.510 79.230 37.790 79.510 ;
        RECT 38.910 79.750 39.190 80.030 ;
        RECT 38.910 79.230 39.190 79.510 ;
        RECT 40.310 79.750 40.590 80.030 ;
        RECT 40.310 79.230 40.590 79.510 ;
        RECT 41.710 85.870 41.990 86.150 ;
        RECT 41.710 85.350 41.990 85.630 ;
        RECT 43.110 85.870 43.390 86.150 ;
        RECT 43.110 85.350 43.390 85.630 ;
        RECT 44.510 88.930 44.790 89.210 ;
        RECT 44.510 88.410 44.790 88.690 ;
        RECT 45.910 82.810 46.190 83.090 ;
        RECT 45.910 82.290 46.190 82.570 ;
        RECT 47.310 76.690 47.590 76.970 ;
        RECT 47.310 76.170 47.590 76.450 ;
        RECT 48.710 88.930 48.990 89.210 ;
        RECT 48.710 88.410 48.990 88.690 ;
        RECT 50.110 85.870 50.390 86.150 ;
        RECT 50.110 85.350 50.390 85.630 ;
        RECT 51.510 85.870 51.790 86.150 ;
        RECT 51.510 85.350 51.790 85.630 ;
        RECT 52.910 79.750 53.190 80.030 ;
        RECT 52.910 79.230 53.190 79.510 ;
        RECT 54.310 79.750 54.590 80.030 ;
        RECT 54.310 79.230 54.590 79.510 ;
        RECT 55.710 79.750 55.990 80.030 ;
        RECT 55.710 79.230 55.990 79.510 ;
        RECT 57.110 79.750 57.390 80.030 ;
        RECT 57.110 79.230 57.390 79.510 ;
        RECT 58.900 91.750 59.180 92.030 ;
        RECT 59.420 91.750 59.700 92.030 ;
        RECT 58.900 88.690 59.180 88.970 ;
        RECT 59.420 88.690 59.700 88.970 ;
        RECT 58.900 85.630 59.180 85.910 ;
        RECT 59.420 85.630 59.700 85.910 ;
        RECT 58.900 82.570 59.180 82.850 ;
        RECT 59.420 82.570 59.700 82.850 ;
        RECT 58.900 79.510 59.180 79.790 ;
        RECT 59.420 79.510 59.700 79.790 ;
        RECT 58.900 76.450 59.180 76.730 ;
        RECT 59.420 76.450 59.700 76.730 ;
        RECT 12.310 66.440 12.590 66.720 ;
        RECT 12.310 65.920 12.590 66.200 ;
        RECT 13.710 62.350 13.990 62.630 ;
        RECT 13.710 61.830 13.990 62.110 ;
        RECT 15.110 62.350 15.390 62.630 ;
        RECT 15.110 61.830 15.390 62.110 ;
        RECT 16.510 62.350 16.790 62.630 ;
        RECT 16.510 61.830 16.790 62.110 ;
        RECT 17.910 62.350 18.190 62.630 ;
        RECT 17.910 61.830 18.190 62.110 ;
        RECT 19.310 68.470 19.590 68.750 ;
        RECT 19.310 67.950 19.590 68.230 ;
        RECT 20.710 68.470 20.990 68.750 ;
        RECT 20.710 67.950 20.990 68.230 ;
        RECT 22.110 71.530 22.390 71.810 ;
        RECT 22.110 71.010 22.390 71.290 ;
        RECT 23.510 74.590 23.790 74.870 ;
        RECT 23.510 74.070 23.790 74.350 ;
        RECT 24.910 65.410 25.190 65.690 ;
        RECT 24.910 64.890 25.190 65.170 ;
        RECT 26.310 71.530 26.590 71.810 ;
        RECT 26.310 71.010 26.590 71.290 ;
        RECT 27.710 68.470 27.990 68.750 ;
        RECT 27.710 67.950 27.990 68.230 ;
        RECT 29.110 68.470 29.390 68.750 ;
        RECT 29.110 67.950 29.390 68.230 ;
        RECT 30.510 62.350 30.790 62.630 ;
        RECT 30.510 61.830 30.790 62.110 ;
        RECT 31.910 62.350 32.190 62.630 ;
        RECT 31.910 61.830 32.190 62.110 ;
        RECT 33.310 62.350 33.590 62.630 ;
        RECT 33.310 61.830 33.590 62.110 ;
        RECT 34.710 62.350 34.990 62.630 ;
        RECT 34.710 61.830 34.990 62.110 ;
        RECT 36.110 62.350 36.390 62.630 ;
        RECT 36.110 61.830 36.390 62.110 ;
        RECT 37.510 62.350 37.790 62.630 ;
        RECT 37.510 61.830 37.790 62.110 ;
        RECT 38.910 62.350 39.190 62.630 ;
        RECT 38.910 61.830 39.190 62.110 ;
        RECT 40.310 62.350 40.590 62.630 ;
        RECT 40.310 61.830 40.590 62.110 ;
        RECT 41.710 68.470 41.990 68.750 ;
        RECT 41.710 67.950 41.990 68.230 ;
        RECT 43.110 68.470 43.390 68.750 ;
        RECT 43.110 67.950 43.390 68.230 ;
        RECT 44.510 71.530 44.790 71.810 ;
        RECT 44.510 71.010 44.790 71.290 ;
        RECT 45.910 65.410 46.190 65.690 ;
        RECT 45.910 64.890 46.190 65.170 ;
        RECT 47.310 59.290 47.590 59.570 ;
        RECT 47.310 58.770 47.590 59.050 ;
        RECT 48.710 71.530 48.990 71.810 ;
        RECT 48.710 71.010 48.990 71.290 ;
        RECT 50.110 68.470 50.390 68.750 ;
        RECT 50.110 67.950 50.390 68.230 ;
        RECT 51.510 68.470 51.790 68.750 ;
        RECT 51.510 67.950 51.790 68.230 ;
        RECT 52.910 62.350 53.190 62.630 ;
        RECT 52.910 61.830 53.190 62.110 ;
        RECT 54.310 62.350 54.590 62.630 ;
        RECT 54.310 61.830 54.590 62.110 ;
        RECT 55.710 62.350 55.990 62.630 ;
        RECT 55.710 61.830 55.990 62.110 ;
        RECT 57.110 62.350 57.390 62.630 ;
        RECT 57.110 61.830 57.390 62.110 ;
        RECT 58.900 74.350 59.180 74.630 ;
        RECT 59.420 74.350 59.700 74.630 ;
        RECT 58.900 71.290 59.180 71.570 ;
        RECT 59.420 71.290 59.700 71.570 ;
        RECT 58.900 68.230 59.180 68.510 ;
        RECT 59.420 68.230 59.700 68.510 ;
        RECT 58.900 65.170 59.180 65.450 ;
        RECT 59.420 65.170 59.700 65.450 ;
        RECT 58.900 62.110 59.180 62.390 ;
        RECT 59.420 62.110 59.700 62.390 ;
        RECT 12.310 49.040 12.590 49.320 ;
        RECT 12.310 48.520 12.590 48.800 ;
        RECT 13.710 44.950 13.990 45.230 ;
        RECT 13.710 44.430 13.990 44.710 ;
        RECT 15.110 44.950 15.390 45.230 ;
        RECT 15.110 44.430 15.390 44.710 ;
        RECT 16.510 44.950 16.790 45.230 ;
        RECT 16.510 44.430 16.790 44.710 ;
        RECT 17.910 44.950 18.190 45.230 ;
        RECT 17.910 44.430 18.190 44.710 ;
        RECT 19.310 51.070 19.590 51.350 ;
        RECT 19.310 50.550 19.590 50.830 ;
        RECT 20.710 51.070 20.990 51.350 ;
        RECT 20.710 50.550 20.990 50.830 ;
        RECT 22.110 54.130 22.390 54.410 ;
        RECT 22.110 53.610 22.390 53.890 ;
        RECT 23.510 57.190 23.790 57.470 ;
        RECT 23.510 56.670 23.790 56.950 ;
        RECT 24.910 48.010 25.190 48.290 ;
        RECT 24.910 47.490 25.190 47.770 ;
        RECT 26.310 54.130 26.590 54.410 ;
        RECT 26.310 53.610 26.590 53.890 ;
        RECT 27.710 51.070 27.990 51.350 ;
        RECT 27.710 50.550 27.990 50.830 ;
        RECT 29.110 51.070 29.390 51.350 ;
        RECT 29.110 50.550 29.390 50.830 ;
        RECT 30.510 44.950 30.790 45.230 ;
        RECT 30.510 44.430 30.790 44.710 ;
        RECT 31.910 44.950 32.190 45.230 ;
        RECT 31.910 44.430 32.190 44.710 ;
        RECT 33.310 44.950 33.590 45.230 ;
        RECT 33.310 44.430 33.590 44.710 ;
        RECT 34.710 44.950 34.990 45.230 ;
        RECT 34.710 44.430 34.990 44.710 ;
        RECT 36.110 44.950 36.390 45.230 ;
        RECT 36.110 44.430 36.390 44.710 ;
        RECT 37.510 44.950 37.790 45.230 ;
        RECT 37.510 44.430 37.790 44.710 ;
        RECT 38.910 44.950 39.190 45.230 ;
        RECT 38.910 44.430 39.190 44.710 ;
        RECT 40.310 44.950 40.590 45.230 ;
        RECT 40.310 44.430 40.590 44.710 ;
        RECT 41.710 51.070 41.990 51.350 ;
        RECT 41.710 50.550 41.990 50.830 ;
        RECT 43.110 51.070 43.390 51.350 ;
        RECT 43.110 50.550 43.390 50.830 ;
        RECT 44.510 54.130 44.790 54.410 ;
        RECT 44.510 53.610 44.790 53.890 ;
        RECT 45.910 48.010 46.190 48.290 ;
        RECT 45.910 47.490 46.190 47.770 ;
        RECT 47.310 41.890 47.590 42.170 ;
        RECT 47.310 41.370 47.590 41.650 ;
        RECT 48.710 54.130 48.990 54.410 ;
        RECT 48.710 53.610 48.990 53.890 ;
        RECT 50.110 51.070 50.390 51.350 ;
        RECT 50.110 50.550 50.390 50.830 ;
        RECT 51.510 51.070 51.790 51.350 ;
        RECT 51.510 50.550 51.790 50.830 ;
        RECT 52.910 44.950 53.190 45.230 ;
        RECT 52.910 44.430 53.190 44.710 ;
        RECT 54.310 44.950 54.590 45.230 ;
        RECT 54.310 44.430 54.590 44.710 ;
        RECT 55.710 44.950 55.990 45.230 ;
        RECT 55.710 44.430 55.990 44.710 ;
        RECT 57.110 44.950 57.390 45.230 ;
        RECT 57.110 44.430 57.390 44.710 ;
        RECT 64.290 91.990 64.570 92.270 ;
        RECT 64.290 91.470 64.570 91.750 ;
        RECT 64.290 88.930 64.570 89.210 ;
        RECT 64.290 88.410 64.570 88.690 ;
        RECT 65.190 85.870 65.470 86.150 ;
        RECT 65.190 85.350 65.470 85.630 ;
        RECT 64.290 82.810 64.570 83.090 ;
        RECT 64.290 82.290 64.570 82.570 ;
        RECT 63.390 79.750 63.670 80.030 ;
        RECT 63.390 79.230 63.670 79.510 ;
        RECT 64.290 76.690 64.570 76.970 ;
        RECT 64.290 76.170 64.570 76.450 ;
        RECT 66.990 71.530 67.270 71.810 ;
        RECT 66.990 71.010 67.270 71.290 ;
        RECT 66.090 68.470 66.370 68.750 ;
        RECT 66.090 67.950 66.370 68.230 ;
        RECT 68.790 74.590 69.070 74.870 ;
        RECT 68.790 74.070 69.070 74.350 ;
        RECT 72.050 74.590 72.330 74.870 ;
        RECT 72.050 74.070 72.330 74.350 ;
        RECT 73.850 71.530 74.130 71.810 ;
        RECT 73.850 71.010 74.130 71.290 ;
        RECT 76.550 91.990 76.830 92.270 ;
        RECT 76.550 91.470 76.830 91.750 ;
        RECT 76.550 88.930 76.830 89.210 ;
        RECT 76.550 88.410 76.830 88.690 ;
        RECT 75.650 85.870 75.930 86.150 ;
        RECT 75.650 85.350 75.930 85.630 ;
        RECT 76.550 82.810 76.830 83.090 ;
        RECT 76.550 82.290 76.830 82.570 ;
        RECT 77.450 79.750 77.730 80.030 ;
        RECT 77.450 79.230 77.730 79.510 ;
        RECT 76.550 76.690 76.830 76.970 ;
        RECT 76.550 76.170 76.830 76.450 ;
        RECT 74.750 68.470 75.030 68.750 ;
        RECT 74.750 67.950 75.030 68.230 ;
        RECT 67.890 65.410 68.170 65.690 ;
        RECT 67.890 64.890 68.170 65.170 ;
        RECT 72.950 65.410 73.230 65.690 ;
        RECT 72.950 64.890 73.230 65.170 ;
        RECT 62.490 62.350 62.770 62.630 ;
        RECT 62.490 61.830 62.770 62.110 ;
        RECT 78.350 62.350 78.630 62.630 ;
        RECT 78.350 61.830 78.630 62.110 ;
        RECT 80.150 109.390 80.430 109.670 ;
        RECT 80.150 108.870 80.430 109.150 ;
        RECT 81.420 109.150 81.700 109.430 ;
        RECT 81.940 109.150 82.220 109.430 ;
        RECT 80.150 106.330 80.430 106.610 ;
        RECT 80.150 105.810 80.430 106.090 ;
        RECT 81.420 106.090 81.700 106.370 ;
        RECT 81.940 106.090 82.220 106.370 ;
        RECT 80.150 103.270 80.430 103.550 ;
        RECT 80.150 102.750 80.430 103.030 ;
        RECT 81.420 103.030 81.700 103.310 ;
        RECT 81.940 103.030 82.220 103.310 ;
        RECT 80.150 100.210 80.430 100.490 ;
        RECT 80.150 99.690 80.430 99.970 ;
        RECT 81.420 99.970 81.700 100.250 ;
        RECT 81.940 99.970 82.220 100.250 ;
        RECT 80.150 97.150 80.430 97.430 ;
        RECT 80.150 96.630 80.430 96.910 ;
        RECT 81.420 96.910 81.700 97.190 ;
        RECT 81.940 96.910 82.220 97.190 ;
        RECT 80.150 94.090 80.430 94.370 ;
        RECT 80.150 93.570 80.430 93.850 ;
        RECT 81.420 93.850 81.700 94.130 ;
        RECT 81.940 93.850 82.220 94.130 ;
        RECT 83.730 97.150 84.010 97.430 ;
        RECT 83.730 96.630 84.010 96.910 ;
        RECT 85.130 97.150 85.410 97.430 ;
        RECT 85.130 96.630 85.410 96.910 ;
        RECT 86.530 97.150 86.810 97.430 ;
        RECT 86.530 96.630 86.810 96.910 ;
        RECT 87.930 97.150 88.210 97.430 ;
        RECT 87.930 96.630 88.210 96.910 ;
        RECT 89.330 103.270 89.610 103.550 ;
        RECT 89.330 102.750 89.610 103.030 ;
        RECT 90.730 103.270 91.010 103.550 ;
        RECT 90.730 102.750 91.010 103.030 ;
        RECT 92.130 106.330 92.410 106.610 ;
        RECT 92.130 105.810 92.410 106.090 ;
        RECT 93.530 94.090 93.810 94.370 ;
        RECT 93.530 93.570 93.810 93.850 ;
        RECT 94.930 100.210 95.210 100.490 ;
        RECT 94.930 99.690 95.210 99.970 ;
        RECT 96.330 106.330 96.610 106.610 ;
        RECT 96.330 105.810 96.610 106.090 ;
        RECT 97.730 103.270 98.010 103.550 ;
        RECT 97.730 102.750 98.010 103.030 ;
        RECT 99.130 103.270 99.410 103.550 ;
        RECT 99.130 102.750 99.410 103.030 ;
        RECT 100.530 97.150 100.810 97.430 ;
        RECT 100.530 96.630 100.810 96.910 ;
        RECT 101.930 97.150 102.210 97.430 ;
        RECT 101.930 96.630 102.210 96.910 ;
        RECT 103.330 97.150 103.610 97.430 ;
        RECT 103.330 96.630 103.610 96.910 ;
        RECT 104.730 97.150 105.010 97.430 ;
        RECT 104.730 96.630 105.010 96.910 ;
        RECT 106.130 97.150 106.410 97.430 ;
        RECT 106.130 96.630 106.410 96.910 ;
        RECT 107.530 97.150 107.810 97.430 ;
        RECT 107.530 96.630 107.810 96.910 ;
        RECT 108.930 97.150 109.210 97.430 ;
        RECT 108.930 96.630 109.210 96.910 ;
        RECT 110.330 97.150 110.610 97.430 ;
        RECT 110.330 96.630 110.610 96.910 ;
        RECT 111.730 103.270 112.010 103.550 ;
        RECT 111.730 102.750 112.010 103.030 ;
        RECT 113.130 103.270 113.410 103.550 ;
        RECT 113.130 102.750 113.410 103.030 ;
        RECT 114.530 106.330 114.810 106.610 ;
        RECT 114.530 105.810 114.810 106.090 ;
        RECT 115.930 100.210 116.210 100.490 ;
        RECT 115.930 99.690 116.210 99.970 ;
        RECT 117.330 109.390 117.610 109.670 ;
        RECT 117.330 108.870 117.610 109.150 ;
        RECT 118.730 106.330 119.010 106.610 ;
        RECT 118.730 105.810 119.010 106.090 ;
        RECT 120.130 103.270 120.410 103.550 ;
        RECT 120.130 102.750 120.410 103.030 ;
        RECT 121.530 103.270 121.810 103.550 ;
        RECT 121.530 102.750 121.810 103.030 ;
        RECT 122.930 97.150 123.210 97.430 ;
        RECT 122.930 96.630 123.210 96.910 ;
        RECT 124.330 97.150 124.610 97.430 ;
        RECT 124.330 96.630 124.610 96.910 ;
        RECT 125.730 97.150 126.010 97.430 ;
        RECT 125.730 96.630 126.010 96.910 ;
        RECT 127.130 97.150 127.410 97.430 ;
        RECT 127.130 96.630 127.410 96.910 ;
        RECT 128.530 101.240 128.810 101.520 ;
        RECT 128.530 100.720 128.810 101.000 ;
        RECT 143.740 115.620 144.020 115.900 ;
        RECT 144.260 115.620 144.540 115.900 ;
        RECT 147.700 117.380 147.980 117.660 ;
        RECT 148.220 117.380 148.500 117.660 ;
        RECT 147.700 116.500 147.980 116.780 ;
        RECT 148.220 116.500 148.500 116.780 ;
        RECT 149.860 114.300 150.140 114.580 ;
        RECT 150.380 114.300 150.660 114.580 ;
        RECT 143.740 112.100 144.020 112.380 ;
        RECT 144.260 112.100 144.540 112.380 ;
        RECT 147.700 112.100 147.980 112.380 ;
        RECT 148.220 112.100 148.500 112.380 ;
        RECT 143.740 110.340 144.020 110.620 ;
        RECT 144.260 110.340 144.540 110.620 ;
        RECT 147.700 110.340 147.980 110.620 ;
        RECT 148.220 110.340 148.500 110.620 ;
        RECT 143.740 106.820 144.020 107.100 ;
        RECT 144.260 106.820 144.540 107.100 ;
        RECT 147.700 106.820 147.980 107.100 ;
        RECT 148.220 106.820 148.500 107.100 ;
        RECT 143.740 103.300 144.020 103.580 ;
        RECT 144.260 103.300 144.540 103.580 ;
        RECT 147.700 103.300 147.980 103.580 ;
        RECT 148.220 103.300 148.500 103.580 ;
        RECT 143.740 101.540 144.020 101.820 ;
        RECT 144.260 101.540 144.540 101.820 ;
        RECT 147.700 101.540 147.980 101.820 ;
        RECT 148.220 101.540 148.500 101.820 ;
        RECT 147.700 100.660 147.980 100.940 ;
        RECT 148.220 100.660 148.500 100.940 ;
        RECT 143.740 98.020 144.020 98.300 ;
        RECT 144.260 98.020 144.540 98.300 ;
        RECT 147.700 98.020 147.980 98.300 ;
        RECT 148.220 98.020 148.500 98.300 ;
        RECT 143.740 96.260 144.020 96.540 ;
        RECT 144.260 96.260 144.540 96.540 ;
        RECT 147.700 96.260 147.980 96.540 ;
        RECT 148.220 96.260 148.500 96.540 ;
        RECT 141.580 94.940 141.860 95.220 ;
        RECT 142.100 94.940 142.380 95.220 ;
        RECT 81.420 91.750 81.700 92.030 ;
        RECT 81.940 91.750 82.220 92.030 ;
        RECT 81.420 88.690 81.700 88.970 ;
        RECT 81.940 88.690 82.220 88.970 ;
        RECT 81.420 85.630 81.700 85.910 ;
        RECT 81.940 85.630 82.220 85.910 ;
        RECT 81.420 82.570 81.700 82.850 ;
        RECT 81.940 82.570 82.220 82.850 ;
        RECT 81.420 79.510 81.700 79.790 ;
        RECT 81.940 79.510 82.220 79.790 ;
        RECT 81.420 76.450 81.700 76.730 ;
        RECT 81.940 76.450 82.220 76.730 ;
        RECT 83.730 79.750 84.010 80.030 ;
        RECT 83.730 79.230 84.010 79.510 ;
        RECT 85.130 79.750 85.410 80.030 ;
        RECT 85.130 79.230 85.410 79.510 ;
        RECT 86.530 79.750 86.810 80.030 ;
        RECT 86.530 79.230 86.810 79.510 ;
        RECT 87.930 79.750 88.210 80.030 ;
        RECT 87.930 79.230 88.210 79.510 ;
        RECT 89.330 85.870 89.610 86.150 ;
        RECT 89.330 85.350 89.610 85.630 ;
        RECT 90.730 85.870 91.010 86.150 ;
        RECT 90.730 85.350 91.010 85.630 ;
        RECT 92.130 88.930 92.410 89.210 ;
        RECT 92.130 88.410 92.410 88.690 ;
        RECT 93.530 76.690 93.810 76.970 ;
        RECT 93.530 76.170 93.810 76.450 ;
        RECT 94.930 82.810 95.210 83.090 ;
        RECT 94.930 82.290 95.210 82.570 ;
        RECT 96.330 88.930 96.610 89.210 ;
        RECT 96.330 88.410 96.610 88.690 ;
        RECT 97.730 85.870 98.010 86.150 ;
        RECT 97.730 85.350 98.010 85.630 ;
        RECT 99.130 85.870 99.410 86.150 ;
        RECT 99.130 85.350 99.410 85.630 ;
        RECT 100.530 79.750 100.810 80.030 ;
        RECT 100.530 79.230 100.810 79.510 ;
        RECT 101.930 79.750 102.210 80.030 ;
        RECT 101.930 79.230 102.210 79.510 ;
        RECT 103.330 79.750 103.610 80.030 ;
        RECT 103.330 79.230 103.610 79.510 ;
        RECT 104.730 79.750 105.010 80.030 ;
        RECT 104.730 79.230 105.010 79.510 ;
        RECT 106.130 79.750 106.410 80.030 ;
        RECT 106.130 79.230 106.410 79.510 ;
        RECT 107.530 79.750 107.810 80.030 ;
        RECT 107.530 79.230 107.810 79.510 ;
        RECT 108.930 79.750 109.210 80.030 ;
        RECT 108.930 79.230 109.210 79.510 ;
        RECT 110.330 79.750 110.610 80.030 ;
        RECT 110.330 79.230 110.610 79.510 ;
        RECT 111.730 85.870 112.010 86.150 ;
        RECT 111.730 85.350 112.010 85.630 ;
        RECT 113.130 85.870 113.410 86.150 ;
        RECT 113.130 85.350 113.410 85.630 ;
        RECT 114.530 88.930 114.810 89.210 ;
        RECT 114.530 88.410 114.810 88.690 ;
        RECT 115.930 82.810 116.210 83.090 ;
        RECT 115.930 82.290 116.210 82.570 ;
        RECT 117.330 91.990 117.610 92.270 ;
        RECT 117.330 91.470 117.610 91.750 ;
        RECT 118.730 88.930 119.010 89.210 ;
        RECT 118.730 88.410 119.010 88.690 ;
        RECT 120.130 85.870 120.410 86.150 ;
        RECT 120.130 85.350 120.410 85.630 ;
        RECT 121.530 85.870 121.810 86.150 ;
        RECT 121.530 85.350 121.810 85.630 ;
        RECT 122.930 79.750 123.210 80.030 ;
        RECT 122.930 79.230 123.210 79.510 ;
        RECT 124.330 79.750 124.610 80.030 ;
        RECT 124.330 79.230 124.610 79.510 ;
        RECT 125.730 79.750 126.010 80.030 ;
        RECT 125.730 79.230 126.010 79.510 ;
        RECT 127.130 79.750 127.410 80.030 ;
        RECT 127.130 79.230 127.410 79.510 ;
        RECT 128.530 83.840 128.810 84.120 ;
        RECT 128.530 83.320 128.810 83.600 ;
        RECT 143.740 90.980 144.020 91.260 ;
        RECT 144.260 90.980 144.540 91.260 ;
        RECT 147.700 92.740 147.980 93.020 ;
        RECT 148.220 92.740 148.500 93.020 ;
        RECT 147.700 91.860 147.980 92.140 ;
        RECT 148.220 91.860 148.500 92.140 ;
        RECT 149.860 89.660 150.140 89.940 ;
        RECT 150.380 89.660 150.660 89.940 ;
        RECT 143.740 87.460 144.020 87.740 ;
        RECT 144.260 87.460 144.540 87.740 ;
        RECT 147.700 87.460 147.980 87.740 ;
        RECT 148.220 87.460 148.500 87.740 ;
        RECT 143.740 85.700 144.020 85.980 ;
        RECT 144.260 85.700 144.540 85.980 ;
        RECT 147.700 85.700 147.980 85.980 ;
        RECT 148.220 85.700 148.500 85.980 ;
        RECT 143.740 82.180 144.020 82.460 ;
        RECT 144.260 82.180 144.540 82.460 ;
        RECT 147.700 82.180 147.980 82.460 ;
        RECT 148.220 82.180 148.500 82.460 ;
        RECT 143.740 78.660 144.020 78.940 ;
        RECT 144.260 78.660 144.540 78.940 ;
        RECT 147.700 78.660 147.980 78.940 ;
        RECT 148.220 78.660 148.500 78.940 ;
        RECT 143.740 76.900 144.020 77.180 ;
        RECT 144.260 76.900 144.540 77.180 ;
        RECT 147.700 76.900 147.980 77.180 ;
        RECT 148.220 76.900 148.500 77.180 ;
        RECT 147.700 76.020 147.980 76.300 ;
        RECT 148.220 76.020 148.500 76.300 ;
        RECT 81.420 74.350 81.700 74.630 ;
        RECT 81.940 74.350 82.220 74.630 ;
        RECT 81.420 71.290 81.700 71.570 ;
        RECT 81.940 71.290 82.220 71.570 ;
        RECT 81.420 68.230 81.700 68.510 ;
        RECT 81.940 68.230 82.220 68.510 ;
        RECT 81.420 65.170 81.700 65.450 ;
        RECT 81.940 65.170 82.220 65.450 ;
        RECT 81.420 62.110 81.700 62.390 ;
        RECT 81.940 62.110 82.220 62.390 ;
        RECT 83.730 62.350 84.010 62.630 ;
        RECT 83.730 61.830 84.010 62.110 ;
        RECT 58.900 56.950 59.180 57.230 ;
        RECT 59.420 56.950 59.700 57.230 ;
        RECT 61.590 57.190 61.870 57.470 ;
        RECT 61.590 56.670 61.870 56.950 ;
        RECT 79.250 57.190 79.530 57.470 ;
        RECT 85.130 62.350 85.410 62.630 ;
        RECT 85.130 61.830 85.410 62.110 ;
        RECT 86.530 62.350 86.810 62.630 ;
        RECT 86.530 61.830 86.810 62.110 ;
        RECT 87.930 62.350 88.210 62.630 ;
        RECT 87.930 61.830 88.210 62.110 ;
        RECT 89.330 68.470 89.610 68.750 ;
        RECT 89.330 67.950 89.610 68.230 ;
        RECT 90.730 68.470 91.010 68.750 ;
        RECT 90.730 67.950 91.010 68.230 ;
        RECT 92.130 71.530 92.410 71.810 ;
        RECT 92.130 71.010 92.410 71.290 ;
        RECT 93.530 59.290 93.810 59.570 ;
        RECT 93.530 58.770 93.810 59.050 ;
        RECT 94.930 65.410 95.210 65.690 ;
        RECT 94.930 64.890 95.210 65.170 ;
        RECT 96.330 71.530 96.610 71.810 ;
        RECT 96.330 71.010 96.610 71.290 ;
        RECT 97.730 68.470 98.010 68.750 ;
        RECT 97.730 67.950 98.010 68.230 ;
        RECT 99.130 68.470 99.410 68.750 ;
        RECT 99.130 67.950 99.410 68.230 ;
        RECT 100.530 62.350 100.810 62.630 ;
        RECT 100.530 61.830 100.810 62.110 ;
        RECT 101.930 62.350 102.210 62.630 ;
        RECT 101.930 61.830 102.210 62.110 ;
        RECT 103.330 62.350 103.610 62.630 ;
        RECT 103.330 61.830 103.610 62.110 ;
        RECT 104.730 62.350 105.010 62.630 ;
        RECT 104.730 61.830 105.010 62.110 ;
        RECT 106.130 62.350 106.410 62.630 ;
        RECT 106.130 61.830 106.410 62.110 ;
        RECT 107.530 62.350 107.810 62.630 ;
        RECT 107.530 61.830 107.810 62.110 ;
        RECT 108.930 62.350 109.210 62.630 ;
        RECT 108.930 61.830 109.210 62.110 ;
        RECT 110.330 62.350 110.610 62.630 ;
        RECT 110.330 61.830 110.610 62.110 ;
        RECT 111.730 68.470 112.010 68.750 ;
        RECT 111.730 67.950 112.010 68.230 ;
        RECT 113.130 68.470 113.410 68.750 ;
        RECT 113.130 67.950 113.410 68.230 ;
        RECT 114.530 71.530 114.810 71.810 ;
        RECT 114.530 71.010 114.810 71.290 ;
        RECT 115.930 65.410 116.210 65.690 ;
        RECT 115.930 64.890 116.210 65.170 ;
        RECT 117.330 74.590 117.610 74.870 ;
        RECT 117.330 74.070 117.610 74.350 ;
        RECT 118.730 71.530 119.010 71.810 ;
        RECT 118.730 71.010 119.010 71.290 ;
        RECT 120.130 68.470 120.410 68.750 ;
        RECT 120.130 67.950 120.410 68.230 ;
        RECT 121.530 68.470 121.810 68.750 ;
        RECT 121.530 67.950 121.810 68.230 ;
        RECT 122.930 62.350 123.210 62.630 ;
        RECT 122.930 61.830 123.210 62.110 ;
        RECT 124.330 62.350 124.610 62.630 ;
        RECT 124.330 61.830 124.610 62.110 ;
        RECT 125.730 62.350 126.010 62.630 ;
        RECT 125.730 61.830 126.010 62.110 ;
        RECT 127.130 62.350 127.410 62.630 ;
        RECT 127.130 61.830 127.410 62.110 ;
        RECT 143.740 73.380 144.020 73.660 ;
        RECT 144.260 73.380 144.540 73.660 ;
        RECT 147.700 73.380 147.980 73.660 ;
        RECT 148.220 73.380 148.500 73.660 ;
        RECT 143.740 71.620 144.020 71.900 ;
        RECT 144.260 71.620 144.540 71.900 ;
        RECT 147.700 71.620 147.980 71.900 ;
        RECT 148.220 71.620 148.500 71.900 ;
        RECT 141.580 70.300 141.860 70.580 ;
        RECT 142.100 70.300 142.380 70.580 ;
        RECT 128.530 66.440 128.810 66.720 ;
        RECT 128.530 65.920 128.810 66.200 ;
        RECT 79.250 56.670 79.530 56.950 ;
        RECT 81.420 56.950 81.700 57.230 ;
        RECT 81.940 56.950 82.220 57.230 ;
        RECT 58.900 53.890 59.180 54.170 ;
        RECT 59.420 53.890 59.700 54.170 ;
        RECT 61.590 54.130 61.870 54.410 ;
        RECT 61.590 53.610 61.870 53.890 ;
        RECT 79.250 54.130 79.530 54.410 ;
        RECT 79.250 53.610 79.530 53.890 ;
        RECT 81.420 53.890 81.700 54.170 ;
        RECT 81.940 53.890 82.220 54.170 ;
        RECT 58.900 50.830 59.180 51.110 ;
        RECT 59.420 50.830 59.700 51.110 ;
        RECT 61.590 51.070 61.870 51.350 ;
        RECT 61.590 50.550 61.870 50.830 ;
        RECT 79.250 51.070 79.530 51.350 ;
        RECT 79.250 50.550 79.530 50.830 ;
        RECT 81.420 50.830 81.700 51.110 ;
        RECT 81.940 50.830 82.220 51.110 ;
        RECT 58.900 47.770 59.180 48.050 ;
        RECT 59.420 47.770 59.700 48.050 ;
        RECT 61.590 48.010 61.870 48.290 ;
        RECT 61.590 47.490 61.870 47.770 ;
        RECT 79.250 48.010 79.530 48.290 ;
        RECT 79.250 47.490 79.530 47.770 ;
        RECT 81.420 47.770 81.700 48.050 ;
        RECT 81.940 47.770 82.220 48.050 ;
        RECT 58.900 44.710 59.180 44.990 ;
        RECT 59.420 44.710 59.700 44.990 ;
        RECT 61.590 44.950 61.870 45.230 ;
        RECT 61.590 44.430 61.870 44.710 ;
        RECT 79.250 44.950 79.530 45.230 ;
        RECT 79.250 44.430 79.530 44.710 ;
        RECT 81.420 44.710 81.700 44.990 ;
        RECT 81.940 44.710 82.220 44.990 ;
        RECT 58.900 41.650 59.180 41.930 ;
        RECT 59.420 41.650 59.700 41.930 ;
        RECT 61.590 41.890 61.870 42.170 ;
        RECT 61.590 41.370 61.870 41.650 ;
        RECT 79.250 41.890 79.530 42.170 ;
        RECT 79.250 41.370 79.530 41.650 ;
        RECT 81.420 41.650 81.700 41.930 ;
        RECT 81.940 41.650 82.220 41.930 ;
        RECT 83.730 44.950 84.010 45.230 ;
        RECT 83.730 44.430 84.010 44.710 ;
        RECT 85.130 44.950 85.410 45.230 ;
        RECT 85.130 44.430 85.410 44.710 ;
        RECT 86.530 44.950 86.810 45.230 ;
        RECT 86.530 44.430 86.810 44.710 ;
        RECT 87.930 44.950 88.210 45.230 ;
        RECT 87.930 44.430 88.210 44.710 ;
        RECT 89.330 51.070 89.610 51.350 ;
        RECT 89.330 50.550 89.610 50.830 ;
        RECT 90.730 51.070 91.010 51.350 ;
        RECT 90.730 50.550 91.010 50.830 ;
        RECT 92.130 54.130 92.410 54.410 ;
        RECT 92.130 53.610 92.410 53.890 ;
        RECT 93.530 41.890 93.810 42.170 ;
        RECT 93.530 41.370 93.810 41.650 ;
        RECT 94.930 48.010 95.210 48.290 ;
        RECT 94.930 47.490 95.210 47.770 ;
        RECT 96.330 54.130 96.610 54.410 ;
        RECT 96.330 53.610 96.610 53.890 ;
        RECT 97.730 51.070 98.010 51.350 ;
        RECT 97.730 50.550 98.010 50.830 ;
        RECT 99.130 51.070 99.410 51.350 ;
        RECT 99.130 50.550 99.410 50.830 ;
        RECT 100.530 44.950 100.810 45.230 ;
        RECT 100.530 44.430 100.810 44.710 ;
        RECT 101.930 44.950 102.210 45.230 ;
        RECT 101.930 44.430 102.210 44.710 ;
        RECT 103.330 44.950 103.610 45.230 ;
        RECT 103.330 44.430 103.610 44.710 ;
        RECT 104.730 44.950 105.010 45.230 ;
        RECT 104.730 44.430 105.010 44.710 ;
        RECT 106.130 44.950 106.410 45.230 ;
        RECT 106.130 44.430 106.410 44.710 ;
        RECT 107.530 44.950 107.810 45.230 ;
        RECT 107.530 44.430 107.810 44.710 ;
        RECT 108.930 44.950 109.210 45.230 ;
        RECT 108.930 44.430 109.210 44.710 ;
        RECT 110.330 44.950 110.610 45.230 ;
        RECT 110.330 44.430 110.610 44.710 ;
        RECT 111.730 51.070 112.010 51.350 ;
        RECT 111.730 50.550 112.010 50.830 ;
        RECT 113.130 51.070 113.410 51.350 ;
        RECT 113.130 50.550 113.410 50.830 ;
        RECT 114.530 54.130 114.810 54.410 ;
        RECT 114.530 53.610 114.810 53.890 ;
        RECT 115.930 48.010 116.210 48.290 ;
        RECT 115.930 47.490 116.210 47.770 ;
        RECT 117.330 57.190 117.610 57.470 ;
        RECT 117.330 56.670 117.610 56.950 ;
        RECT 118.730 54.130 119.010 54.410 ;
        RECT 118.730 53.610 119.010 53.890 ;
        RECT 120.130 51.070 120.410 51.350 ;
        RECT 120.130 50.550 120.410 50.830 ;
        RECT 121.530 51.070 121.810 51.350 ;
        RECT 121.530 50.550 121.810 50.830 ;
        RECT 122.930 44.950 123.210 45.230 ;
        RECT 122.930 44.430 123.210 44.710 ;
        RECT 124.330 44.950 124.610 45.230 ;
        RECT 124.330 44.430 124.610 44.710 ;
        RECT 125.730 44.950 126.010 45.230 ;
        RECT 125.730 44.430 126.010 44.710 ;
        RECT 127.130 44.950 127.410 45.230 ;
        RECT 127.130 44.430 127.410 44.710 ;
        RECT 143.740 66.340 144.020 66.620 ;
        RECT 144.260 66.340 144.540 66.620 ;
        RECT 147.700 68.100 147.980 68.380 ;
        RECT 148.220 68.100 148.500 68.380 ;
        RECT 147.700 67.220 147.980 67.500 ;
        RECT 148.220 67.220 148.500 67.500 ;
        RECT 149.860 65.020 150.140 65.300 ;
        RECT 150.380 65.020 150.660 65.300 ;
        RECT 143.740 62.820 144.020 63.100 ;
        RECT 144.260 62.820 144.540 63.100 ;
        RECT 147.700 62.820 147.980 63.100 ;
        RECT 148.220 62.820 148.500 63.100 ;
        RECT 143.740 61.060 144.020 61.340 ;
        RECT 144.260 61.060 144.540 61.340 ;
        RECT 147.700 61.060 147.980 61.340 ;
        RECT 148.220 61.060 148.500 61.340 ;
        RECT 143.740 57.540 144.020 57.820 ;
        RECT 144.260 57.540 144.540 57.820 ;
        RECT 147.700 57.540 147.980 57.820 ;
        RECT 148.220 57.540 148.500 57.820 ;
        RECT 143.740 54.020 144.020 54.300 ;
        RECT 144.260 54.020 144.540 54.300 ;
        RECT 147.700 54.020 147.980 54.300 ;
        RECT 148.220 54.020 148.500 54.300 ;
        RECT 143.740 52.260 144.020 52.540 ;
        RECT 144.260 52.260 144.540 52.540 ;
        RECT 147.700 52.260 147.980 52.540 ;
        RECT 148.220 52.260 148.500 52.540 ;
        RECT 147.700 51.380 147.980 51.660 ;
        RECT 148.220 51.380 148.500 51.660 ;
        RECT 128.530 49.040 128.810 49.320 ;
        RECT 128.530 48.520 128.810 48.800 ;
        RECT 143.740 48.740 144.020 49.020 ;
        RECT 144.260 48.740 144.540 49.020 ;
        RECT 147.700 48.740 147.980 49.020 ;
        RECT 148.220 48.740 148.500 49.020 ;
        RECT 143.740 46.980 144.020 47.260 ;
        RECT 144.260 46.980 144.540 47.260 ;
        RECT 147.700 46.980 147.980 47.260 ;
        RECT 148.220 46.980 148.500 47.260 ;
        RECT 141.580 45.660 141.860 45.940 ;
        RECT 142.100 45.660 142.380 45.940 ;
        RECT 47.080 38.580 48.160 38.935 ;
        RECT 14.320 37.700 15.400 38.055 ;
        RECT 47.080 36.820 48.160 37.175 ;
        RECT 14.320 35.940 15.400 36.295 ;
        RECT 47.080 35.060 48.160 35.415 ;
        RECT 93.160 38.580 94.240 38.935 ;
        RECT 125.920 37.700 127.000 38.055 ;
        RECT 93.160 36.820 94.240 37.175 ;
        RECT 125.920 35.940 127.000 36.295 ;
        RECT 93.160 35.060 94.240 35.415 ;
        RECT 14.320 34.185 15.400 34.535 ;
        RECT 125.920 34.185 127.000 34.535 ;
        RECT 47.080 33.300 48.160 33.655 ;
        RECT 14.320 32.420 15.400 32.775 ;
        RECT 93.160 33.300 94.240 33.655 ;
        RECT 54.860 32.040 55.140 32.320 ;
        RECT 55.380 32.040 55.660 32.320 ;
        RECT 58.820 32.040 59.100 32.320 ;
        RECT 59.340 32.040 59.620 32.320 ;
        RECT 81.700 32.040 81.980 32.320 ;
        RECT 82.220 32.040 82.500 32.320 ;
        RECT 85.660 32.040 85.940 32.320 ;
        RECT 86.180 32.040 86.460 32.320 ;
        RECT 47.080 31.540 48.160 31.895 ;
        RECT 14.320 30.660 15.400 31.015 ;
        RECT 125.920 32.420 127.000 32.775 ;
        RECT 93.160 31.540 94.240 31.895 ;
        RECT 54.860 31.160 55.140 31.440 ;
        RECT 55.380 31.160 55.660 31.440 ;
        RECT 58.820 31.160 59.100 31.440 ;
        RECT 59.340 31.160 59.620 31.440 ;
        RECT 81.700 31.160 81.980 31.440 ;
        RECT 82.220 31.160 82.500 31.440 ;
        RECT 85.660 31.160 85.940 31.440 ;
        RECT 86.180 31.160 86.460 31.440 ;
        RECT 61.740 30.240 62.020 30.520 ;
        RECT 62.260 30.240 62.540 30.520 ;
        RECT 47.080 29.780 48.160 30.135 ;
        RECT 54.860 29.400 55.140 29.680 ;
        RECT 55.380 29.400 55.660 29.680 ;
        RECT 58.820 29.400 59.100 29.680 ;
        RECT 59.340 29.400 59.620 29.680 ;
        RECT 14.320 28.905 15.400 29.255 ;
        RECT 54.860 28.520 55.140 28.800 ;
        RECT 55.380 28.520 55.660 28.800 ;
        RECT 58.820 28.520 59.100 28.800 ;
        RECT 59.340 28.520 59.620 28.800 ;
        RECT 47.080 28.020 48.160 28.375 ;
        RECT 14.320 27.140 15.400 27.495 ;
        RECT 54.860 27.640 55.140 27.920 ;
        RECT 55.380 27.640 55.660 27.920 ;
        RECT 58.820 27.640 59.100 27.920 ;
        RECT 59.340 27.640 59.620 27.920 ;
        RECT 47.080 26.260 48.160 26.615 ;
        RECT 14.320 25.380 15.400 25.735 ;
        RECT 54.860 25.880 55.140 26.160 ;
        RECT 55.380 25.880 55.660 26.160 ;
        RECT 58.820 25.880 59.100 26.160 ;
        RECT 59.340 25.880 59.620 26.160 ;
        RECT 54.860 25.000 55.140 25.280 ;
        RECT 55.380 25.000 55.660 25.280 ;
        RECT 58.740 25.000 59.020 25.280 ;
        RECT 59.260 25.000 59.540 25.280 ;
        RECT 47.080 24.500 48.160 24.855 ;
        RECT 78.780 30.240 79.060 30.520 ;
        RECT 79.300 30.240 79.580 30.520 ;
        RECT 125.920 30.660 127.000 31.015 ;
        RECT 93.160 29.780 94.240 30.135 ;
        RECT 81.700 29.400 81.980 29.680 ;
        RECT 82.220 29.400 82.500 29.680 ;
        RECT 85.660 29.400 85.940 29.680 ;
        RECT 86.180 29.400 86.460 29.680 ;
        RECT 125.920 28.905 127.000 29.255 ;
        RECT 81.700 28.520 81.980 28.800 ;
        RECT 82.220 28.520 82.500 28.800 ;
        RECT 85.660 28.520 85.940 28.800 ;
        RECT 86.180 28.520 86.460 28.800 ;
        RECT 93.160 28.020 94.240 28.375 ;
        RECT 81.700 27.640 81.980 27.920 ;
        RECT 82.220 27.640 82.500 27.920 ;
        RECT 85.660 27.640 85.940 27.920 ;
        RECT 86.180 27.640 86.460 27.920 ;
        RECT 65.860 25.880 66.140 26.160 ;
        RECT 66.380 25.880 66.660 26.160 ;
        RECT 74.500 25.880 74.780 26.160 ;
        RECT 75.020 25.880 75.300 26.160 ;
        RECT 125.920 27.140 127.000 27.495 ;
        RECT 93.160 26.260 94.240 26.615 ;
        RECT 81.700 25.880 81.980 26.160 ;
        RECT 82.220 25.880 82.500 26.160 ;
        RECT 85.660 25.880 85.940 26.160 ;
        RECT 86.180 25.880 86.460 26.160 ;
        RECT 81.780 25.000 82.060 25.280 ;
        RECT 82.300 25.000 82.580 25.280 ;
        RECT 85.660 25.000 85.940 25.280 ;
        RECT 86.180 25.000 86.460 25.280 ;
        RECT 143.740 41.700 144.020 41.980 ;
        RECT 144.260 41.700 144.540 41.980 ;
        RECT 147.700 43.460 147.980 43.740 ;
        RECT 148.220 43.460 148.500 43.740 ;
        RECT 147.700 42.580 147.980 42.860 ;
        RECT 148.220 42.580 148.500 42.860 ;
        RECT 149.860 40.380 150.140 40.660 ;
        RECT 150.380 40.380 150.660 40.660 ;
        RECT 143.740 38.180 144.020 38.460 ;
        RECT 144.260 38.180 144.540 38.460 ;
        RECT 147.700 38.180 147.980 38.460 ;
        RECT 148.220 38.180 148.500 38.460 ;
        RECT 143.740 36.420 144.020 36.700 ;
        RECT 144.260 36.420 144.540 36.700 ;
        RECT 147.700 36.420 147.980 36.700 ;
        RECT 148.220 36.420 148.500 36.700 ;
        RECT 143.740 32.900 144.020 33.180 ;
        RECT 144.260 32.900 144.540 33.180 ;
        RECT 147.700 32.900 147.980 33.180 ;
        RECT 148.220 32.900 148.500 33.180 ;
        RECT 143.740 29.380 144.020 29.660 ;
        RECT 144.260 29.380 144.540 29.660 ;
        RECT 147.700 29.380 147.980 29.660 ;
        RECT 148.220 29.380 148.500 29.660 ;
        RECT 143.740 27.620 144.020 27.900 ;
        RECT 144.260 27.620 144.540 27.900 ;
        RECT 147.700 27.620 147.980 27.900 ;
        RECT 148.220 27.620 148.500 27.900 ;
        RECT 147.700 26.740 147.980 27.020 ;
        RECT 148.220 26.740 148.500 27.020 ;
        RECT 125.920 25.380 127.000 25.735 ;
        RECT 93.160 24.500 94.240 24.855 ;
        RECT 143.740 24.100 144.020 24.380 ;
        RECT 144.260 24.100 144.540 24.380 ;
        RECT 147.700 24.100 147.980 24.380 ;
        RECT 148.220 24.100 148.500 24.380 ;
        RECT 14.320 23.625 15.400 23.975 ;
        RECT 125.920 23.625 127.000 23.975 ;
        RECT 52.700 23.240 52.980 23.520 ;
        RECT 53.220 23.240 53.500 23.520 ;
        RECT 87.820 23.240 88.100 23.520 ;
        RECT 88.340 23.240 88.620 23.520 ;
        RECT 47.080 22.740 48.160 23.095 ;
        RECT 60.980 22.800 61.260 23.080 ;
        RECT 61.500 22.800 61.780 23.080 ;
        RECT 79.540 22.800 79.820 23.080 ;
        RECT 80.060 22.800 80.340 23.080 ;
        RECT 14.320 21.860 15.400 22.215 ;
        RECT 93.160 22.740 94.240 23.095 ;
        RECT 58.820 22.360 59.100 22.640 ;
        RECT 59.340 22.360 59.620 22.640 ;
        RECT 81.700 22.360 81.980 22.640 ;
        RECT 82.220 22.360 82.500 22.640 ;
        RECT 47.080 20.980 48.160 21.335 ;
        RECT 14.320 20.100 15.400 20.455 ;
        RECT 54.860 20.600 55.140 20.880 ;
        RECT 55.380 20.600 55.660 20.880 ;
        RECT 47.080 19.220 48.160 19.575 ;
        RECT 52.700 19.280 52.980 19.560 ;
        RECT 53.220 19.280 53.500 19.560 ;
        RECT 54.860 18.840 55.140 19.120 ;
        RECT 55.380 18.840 55.660 19.120 ;
        RECT 58.820 18.840 59.100 19.120 ;
        RECT 59.340 18.840 59.620 19.120 ;
        RECT 14.320 18.345 15.400 18.695 ;
        RECT 54.860 17.960 55.140 18.240 ;
        RECT 55.380 17.960 55.660 18.240 ;
        RECT 58.820 17.960 59.100 18.240 ;
        RECT 59.340 17.960 59.620 18.240 ;
        RECT 65.860 18.840 66.140 19.120 ;
        RECT 66.380 18.840 66.660 19.120 ;
        RECT 74.500 18.840 74.780 19.120 ;
        RECT 75.020 18.840 75.300 19.120 ;
        RECT 143.740 22.340 144.020 22.620 ;
        RECT 144.260 22.340 144.540 22.620 ;
        RECT 147.700 22.340 147.980 22.620 ;
        RECT 148.220 22.340 148.500 22.620 ;
        RECT 125.920 21.860 127.000 22.215 ;
        RECT 93.160 20.980 94.240 21.335 ;
        RECT 85.660 20.600 85.940 20.880 ;
        RECT 86.180 20.600 86.460 20.880 ;
        RECT 147.700 21.460 147.980 21.740 ;
        RECT 148.220 21.460 148.500 21.740 ;
        RECT 125.920 20.100 127.000 20.455 ;
        RECT 87.820 19.280 88.100 19.560 ;
        RECT 88.340 19.280 88.620 19.560 ;
        RECT 93.160 19.220 94.240 19.575 ;
        RECT 81.700 18.840 81.980 19.120 ;
        RECT 82.220 18.840 82.500 19.120 ;
        RECT 85.660 18.840 85.940 19.120 ;
        RECT 86.180 18.840 86.460 19.120 ;
        RECT 143.740 18.820 144.020 19.100 ;
        RECT 144.260 18.820 144.540 19.100 ;
        RECT 147.700 18.820 147.980 19.100 ;
        RECT 148.220 18.820 148.500 19.100 ;
        RECT 125.920 18.345 127.000 18.695 ;
        RECT 81.700 17.960 81.980 18.240 ;
        RECT 82.220 17.960 82.500 18.240 ;
        RECT 85.660 17.960 85.940 18.240 ;
        RECT 86.180 17.960 86.460 18.240 ;
        RECT 47.080 17.460 48.160 17.815 ;
        RECT 68.100 17.520 68.380 17.800 ;
        RECT 68.620 17.520 68.900 17.800 ;
        RECT 72.420 17.520 72.700 17.800 ;
        RECT 72.940 17.520 73.220 17.800 ;
        RECT 14.320 16.580 15.400 16.935 ;
        RECT 58.820 16.390 59.100 16.670 ;
        RECT 59.340 16.390 59.620 16.670 ;
        RECT 81.700 16.390 81.980 16.670 ;
        RECT 82.220 16.390 82.500 16.670 ;
        RECT 93.160 17.460 94.240 17.815 ;
        RECT 143.740 17.060 144.020 17.340 ;
        RECT 144.260 17.060 144.540 17.340 ;
        RECT 147.700 17.060 147.980 17.340 ;
        RECT 148.220 17.060 148.500 17.340 ;
        RECT 125.920 16.580 127.000 16.935 ;
        RECT 47.080 15.700 48.160 16.055 ;
        RECT 14.320 14.820 15.400 15.175 ;
        RECT 54.860 15.320 55.140 15.600 ;
        RECT 55.380 15.320 55.660 15.600 ;
        RECT 58.820 15.320 59.100 15.600 ;
        RECT 59.340 15.320 59.620 15.600 ;
        RECT 54.860 14.440 55.140 14.720 ;
        RECT 55.380 14.440 55.660 14.720 ;
        RECT 58.820 14.440 59.100 14.720 ;
        RECT 59.340 14.440 59.620 14.720 ;
        RECT 47.080 13.940 48.160 14.295 ;
        RECT 54.860 13.560 55.140 13.840 ;
        RECT 55.380 13.560 55.660 13.840 ;
        RECT 58.820 13.560 59.100 13.840 ;
        RECT 59.340 13.560 59.620 13.840 ;
        RECT 14.320 13.065 15.400 13.415 ;
        RECT 58.740 10.220 59.020 10.500 ;
        RECT 59.260 10.220 59.540 10.500 ;
        RECT 58.740 9.700 59.020 9.980 ;
        RECT 59.260 9.700 59.540 9.980 ;
        RECT 54.780 6.620 55.060 6.900 ;
        RECT 55.300 6.620 55.580 6.900 ;
        RECT 54.780 6.100 55.060 6.380 ;
        RECT 55.300 6.100 55.580 6.380 ;
        RECT 65.940 14.400 66.220 14.680 ;
        RECT 66.460 14.400 66.740 14.680 ;
        RECT 74.580 14.400 74.860 14.680 ;
        RECT 75.100 14.400 75.380 14.680 ;
        RECT 93.160 15.700 94.240 16.055 ;
        RECT 81.700 15.320 81.980 15.600 ;
        RECT 82.220 15.320 82.500 15.600 ;
        RECT 85.660 15.320 85.940 15.600 ;
        RECT 86.180 15.320 86.460 15.600 ;
        RECT 81.700 14.440 81.980 14.720 ;
        RECT 82.220 14.440 82.500 14.720 ;
        RECT 85.660 14.440 85.940 14.720 ;
        RECT 86.180 14.440 86.460 14.720 ;
        RECT 143.740 15.300 144.020 15.580 ;
        RECT 144.260 15.300 144.540 15.580 ;
        RECT 147.700 15.300 147.980 15.580 ;
        RECT 148.220 15.300 148.500 15.580 ;
        RECT 125.920 14.820 127.000 15.175 ;
        RECT 93.160 13.940 94.240 14.295 ;
        RECT 81.700 13.560 81.980 13.840 ;
        RECT 82.220 13.560 82.500 13.840 ;
        RECT 85.660 13.560 85.940 13.840 ;
        RECT 86.180 13.560 86.460 13.840 ;
        RECT 143.740 14.420 144.020 14.700 ;
        RECT 144.260 14.420 144.540 14.700 ;
        RECT 125.920 13.065 127.000 13.415 ;
        RECT 143.740 11.780 144.020 12.060 ;
        RECT 144.260 11.780 144.540 12.060 ;
        RECT 147.700 11.780 147.980 12.060 ;
        RECT 148.220 11.780 148.500 12.060 ;
        RECT 81.700 10.220 81.980 10.500 ;
        RECT 82.220 10.220 82.500 10.500 ;
        RECT 143.740 10.020 144.020 10.300 ;
        RECT 144.260 10.020 144.540 10.300 ;
        RECT 147.700 10.020 147.980 10.300 ;
        RECT 148.220 10.020 148.500 10.300 ;
        RECT 81.700 9.700 81.980 9.980 ;
        RECT 82.220 9.700 82.500 9.980 ;
        RECT 143.740 9.140 144.020 9.420 ;
        RECT 144.260 9.140 144.540 9.420 ;
        RECT 147.700 9.140 147.980 9.420 ;
        RECT 148.220 9.140 148.500 9.420 ;
        RECT 85.660 6.620 85.940 6.900 ;
        RECT 86.180 6.620 86.460 6.900 ;
        RECT 143.740 6.500 144.020 6.780 ;
        RECT 144.260 6.500 144.540 6.780 ;
        RECT 147.700 6.500 147.980 6.780 ;
        RECT 148.220 6.500 148.500 6.780 ;
        RECT 85.660 6.100 85.940 6.380 ;
        RECT 86.180 6.100 86.460 6.380 ;
        RECT 143.740 4.740 144.020 5.020 ;
        RECT 144.260 4.740 144.540 5.020 ;
        RECT 147.700 4.740 147.980 5.020 ;
        RECT 148.220 4.740 148.500 5.020 ;
        RECT 61.660 4.030 61.940 4.310 ;
        RECT 62.180 4.030 62.460 4.310 ;
        RECT 78.780 4.030 79.060 4.310 ;
        RECT 79.300 4.030 79.580 4.310 ;
        RECT 143.740 3.860 144.020 4.140 ;
        RECT 144.260 3.860 144.540 4.140 ;
        RECT 147.700 3.860 147.980 4.140 ;
        RECT 148.220 3.860 148.500 4.140 ;
        RECT 143.740 2.980 144.020 3.260 ;
        RECT 144.260 2.980 144.540 3.260 ;
        RECT 147.700 2.980 147.980 3.260 ;
        RECT 148.220 2.980 148.500 3.260 ;
      LAYER met2 ;
        RECT 24.580 221.190 25.580 222.190 ;
        RECT 27.540 221.190 28.540 222.190 ;
        RECT 49.780 221.190 50.780 222.190 ;
        RECT 52.740 221.190 53.740 222.190 ;
        RECT 74.980 221.190 75.980 222.190 ;
        RECT 77.940 221.190 78.940 222.190 ;
        RECT 100.180 221.190 101.180 222.190 ;
        RECT 103.140 221.190 104.140 222.190 ;
        RECT 143.680 222.070 144.680 222.450 ;
        RECT 147.640 222.070 148.640 222.450 ;
        RECT 143.680 221.190 144.680 221.570 ;
        RECT 147.640 221.190 148.640 221.570 ;
        RECT 143.680 219.430 144.680 219.810 ;
        RECT 147.640 219.430 148.640 219.810 ;
        RECT 21.700 217.590 22.700 218.590 ;
        RECT 30.420 217.590 31.420 218.590 ;
        RECT 46.900 217.590 47.900 218.590 ;
        RECT 55.620 217.590 56.620 218.590 ;
        RECT 72.100 217.590 73.100 218.590 ;
        RECT 80.820 217.590 81.820 218.590 ;
        RECT 97.300 217.590 98.300 218.590 ;
        RECT 106.020 217.590 107.020 218.590 ;
        RECT 122.500 217.590 123.500 218.590 ;
        RECT 141.520 218.110 143.300 218.490 ;
        RECT 17.740 213.990 18.740 214.990 ;
        RECT 34.380 213.990 35.380 214.990 ;
        RECT 42.940 213.990 43.940 214.990 ;
        RECT 59.580 213.990 60.580 214.990 ;
        RECT 68.140 213.990 69.140 214.990 ;
        RECT 84.780 213.990 85.780 214.990 ;
        RECT 93.340 213.990 94.340 214.990 ;
        RECT 109.980 213.990 110.980 214.990 ;
        RECT 118.540 213.990 119.540 214.990 ;
        RECT 142.920 213.210 143.300 218.110 ;
        RECT 147.640 215.910 148.640 216.290 ;
        RECT 147.640 215.030 148.640 215.410 ;
        RECT 143.680 214.150 144.680 214.530 ;
        RECT 142.920 212.830 150.800 213.210 ;
        RECT 17.740 210.800 18.740 211.180 ;
        RECT 21.700 210.800 22.700 211.180 ;
        RECT 30.420 210.800 31.420 211.180 ;
        RECT 34.380 210.800 35.380 211.180 ;
        RECT 42.940 210.800 43.940 211.180 ;
        RECT 46.900 210.800 47.900 211.180 ;
        RECT 55.620 210.800 56.620 211.180 ;
        RECT 59.580 210.800 60.580 211.180 ;
        RECT 68.140 210.800 69.140 211.180 ;
        RECT 72.100 210.800 73.100 211.180 ;
        RECT 80.820 210.800 81.820 211.180 ;
        RECT 84.780 210.800 85.780 211.180 ;
        RECT 93.340 210.800 94.340 211.180 ;
        RECT 97.300 210.800 98.300 211.180 ;
        RECT 106.020 210.800 107.020 211.180 ;
        RECT 109.980 210.800 110.980 211.180 ;
        RECT 143.680 210.630 144.680 211.010 ;
        RECT 147.640 210.630 148.640 211.010 ;
        RECT 17.740 209.920 18.740 210.300 ;
        RECT 21.700 209.920 22.700 210.300 ;
        RECT 30.420 209.920 31.420 210.300 ;
        RECT 34.380 209.920 35.380 210.300 ;
        RECT 42.940 209.920 43.940 210.300 ;
        RECT 46.900 209.920 47.900 210.300 ;
        RECT 55.620 209.920 56.620 210.300 ;
        RECT 59.580 209.920 60.580 210.300 ;
        RECT 68.140 209.920 69.140 210.300 ;
        RECT 72.100 209.920 73.100 210.300 ;
        RECT 80.820 209.920 81.820 210.300 ;
        RECT 84.780 209.920 85.780 210.300 ;
        RECT 93.340 209.920 94.340 210.300 ;
        RECT 97.300 209.920 98.300 210.300 ;
        RECT 106.020 209.920 107.020 210.300 ;
        RECT 109.980 209.920 110.980 210.300 ;
        RECT 21.700 209.570 22.700 209.610 ;
        RECT 23.420 209.570 23.800 209.610 ;
        RECT 21.700 209.190 23.800 209.570 ;
        RECT 46.900 209.570 47.900 209.610 ;
        RECT 48.620 209.570 49.000 209.610 ;
        RECT 46.900 209.190 49.000 209.570 ;
        RECT 72.100 209.570 73.100 209.610 ;
        RECT 73.820 209.570 74.200 209.610 ;
        RECT 72.100 209.190 74.200 209.570 ;
        RECT 97.300 209.570 98.300 209.610 ;
        RECT 99.020 209.570 99.400 209.610 ;
        RECT 97.300 209.190 99.400 209.570 ;
        RECT 17.740 208.160 18.740 208.540 ;
        RECT 21.700 208.160 22.700 208.540 ;
        RECT 17.740 207.280 18.740 207.660 ;
        RECT 23.420 206.520 23.800 209.190 ;
        RECT 30.420 208.160 31.420 208.540 ;
        RECT 34.380 208.160 35.380 208.540 ;
        RECT 42.940 208.160 43.940 208.540 ;
        RECT 46.900 208.160 47.900 208.540 ;
        RECT 34.380 207.280 35.380 207.660 ;
        RECT 42.940 207.280 43.940 207.660 ;
        RECT 36.460 207.140 37.460 207.220 ;
        RECT 36.080 206.840 37.460 207.140 ;
        RECT 36.080 206.520 36.460 206.840 ;
        RECT 23.420 206.140 36.460 206.520 ;
        RECT 48.620 206.520 49.000 209.190 ;
        RECT 55.620 208.160 56.620 208.540 ;
        RECT 59.580 208.160 60.580 208.540 ;
        RECT 68.140 208.160 69.140 208.540 ;
        RECT 72.100 208.160 73.100 208.540 ;
        RECT 59.580 207.280 60.580 207.660 ;
        RECT 68.140 207.280 69.140 207.660 ;
        RECT 61.660 207.140 62.660 207.220 ;
        RECT 61.280 206.840 62.660 207.140 ;
        RECT 61.280 206.520 61.660 206.840 ;
        RECT 48.620 206.140 61.660 206.520 ;
        RECT 73.820 206.520 74.200 209.190 ;
        RECT 80.820 208.160 81.820 208.540 ;
        RECT 84.780 208.160 85.780 208.540 ;
        RECT 93.340 208.160 94.340 208.540 ;
        RECT 97.300 208.160 98.300 208.540 ;
        RECT 84.780 207.280 85.780 207.660 ;
        RECT 93.340 207.280 94.340 207.660 ;
        RECT 86.860 207.140 87.860 207.220 ;
        RECT 86.480 206.840 87.860 207.140 ;
        RECT 86.480 206.520 86.860 206.840 ;
        RECT 73.820 206.140 86.860 206.520 ;
        RECT 99.020 206.520 99.400 209.190 ;
        RECT 105.940 209.040 114.520 209.420 ;
        RECT 118.540 209.040 119.540 209.420 ;
        RECT 122.500 209.040 123.500 209.420 ;
        RECT 106.020 208.160 107.020 208.540 ;
        RECT 109.980 208.160 110.980 208.540 ;
        RECT 109.980 207.280 110.980 207.660 ;
        RECT 114.140 207.370 114.520 209.040 ;
        RECT 143.680 208.870 144.680 209.250 ;
        RECT 147.640 208.870 148.640 209.250 ;
        RECT 118.540 208.160 119.540 208.540 ;
        RECT 122.500 208.160 123.500 208.540 ;
        RECT 116.380 207.370 117.380 207.410 ;
        RECT 112.060 207.140 113.060 207.220 ;
        RECT 111.680 206.840 113.060 207.140 ;
        RECT 114.140 207.030 117.380 207.370 ;
        RECT 114.140 206.990 116.920 207.030 ;
        RECT 111.680 206.520 112.060 206.840 ;
        RECT 99.020 206.140 112.060 206.520 ;
        RECT 118.540 206.400 119.540 206.780 ;
        RECT 122.500 206.400 123.500 206.780 ;
        RECT 118.540 205.520 119.540 205.900 ;
        RECT 123.960 205.080 125.740 205.460 ;
        RECT 143.680 205.350 144.680 205.730 ;
        RECT 147.640 205.350 148.640 205.730 ;
        RECT 17.740 204.640 18.740 205.020 ;
        RECT 21.700 204.640 22.700 205.020 ;
        RECT 30.420 204.640 31.420 205.020 ;
        RECT 34.380 204.640 35.380 205.020 ;
        RECT 42.940 204.640 43.940 205.020 ;
        RECT 46.900 204.640 47.900 205.020 ;
        RECT 55.620 204.640 56.620 205.020 ;
        RECT 59.580 204.640 60.580 205.020 ;
        RECT 68.140 204.640 69.140 205.020 ;
        RECT 72.100 204.640 73.100 205.020 ;
        RECT 80.820 204.640 81.820 205.020 ;
        RECT 84.780 204.640 85.780 205.020 ;
        RECT 93.340 204.640 94.340 205.020 ;
        RECT 97.300 204.640 98.300 205.020 ;
        RECT 106.020 204.640 107.020 205.020 ;
        RECT 109.980 204.640 110.980 205.020 ;
        RECT 17.740 202.880 18.740 203.260 ;
        RECT 21.700 202.880 22.700 203.260 ;
        RECT 30.420 202.880 31.420 203.260 ;
        RECT 34.380 202.880 35.380 203.260 ;
        RECT 42.940 202.880 43.940 203.260 ;
        RECT 46.900 202.880 47.900 203.260 ;
        RECT 55.620 202.880 56.620 203.260 ;
        RECT 59.580 202.880 60.580 203.260 ;
        RECT 68.140 202.880 69.140 203.260 ;
        RECT 72.100 202.880 73.100 203.260 ;
        RECT 80.820 202.880 81.820 203.260 ;
        RECT 84.780 202.880 85.780 203.260 ;
        RECT 93.340 202.880 94.340 203.260 ;
        RECT 97.300 202.880 98.300 203.260 ;
        RECT 106.020 202.880 107.020 203.260 ;
        RECT 109.980 202.880 110.980 203.260 ;
        RECT 118.540 202.880 119.540 203.260 ;
        RECT 122.500 202.880 123.500 203.260 ;
        RECT 21.700 202.000 22.700 202.380 ;
        RECT 30.420 202.000 31.420 202.380 ;
        RECT 46.900 202.000 47.900 202.380 ;
        RECT 55.620 202.000 56.620 202.380 ;
        RECT 72.100 202.000 73.100 202.380 ;
        RECT 80.820 202.000 81.820 202.380 ;
        RECT 97.300 202.000 98.300 202.380 ;
        RECT 106.020 202.000 107.020 202.380 ;
        RECT 122.500 202.000 123.500 202.380 ;
        RECT 17.740 199.360 18.740 199.740 ;
        RECT 21.700 199.360 22.700 199.740 ;
        RECT 30.420 199.360 31.420 199.740 ;
        RECT 34.380 199.360 35.380 199.740 ;
        RECT 42.940 199.360 43.940 199.740 ;
        RECT 46.900 199.360 47.900 199.740 ;
        RECT 55.620 199.360 56.620 199.740 ;
        RECT 59.580 199.360 60.580 199.740 ;
        RECT 68.140 199.360 69.140 199.740 ;
        RECT 72.100 199.360 73.100 199.740 ;
        RECT 80.820 199.360 81.820 199.740 ;
        RECT 84.780 199.360 85.780 199.740 ;
        RECT 93.340 199.360 94.340 199.740 ;
        RECT 97.300 199.360 98.300 199.740 ;
        RECT 106.020 199.360 107.020 199.740 ;
        RECT 109.980 199.360 110.980 199.740 ;
        RECT 118.540 199.360 119.540 199.740 ;
        RECT 122.500 199.360 123.500 199.740 ;
        RECT 123.960 198.860 124.340 205.080 ;
        RECT 124.660 203.320 126.440 203.700 ;
        RECT 109.980 198.480 124.340 198.860 ;
        RECT 17.740 197.600 18.740 197.980 ;
        RECT 21.700 197.600 22.700 197.980 ;
        RECT 30.420 197.600 31.420 197.980 ;
        RECT 34.380 197.600 35.380 197.980 ;
        RECT 42.940 197.600 43.940 197.980 ;
        RECT 46.900 197.600 47.900 197.980 ;
        RECT 55.620 197.600 56.620 197.980 ;
        RECT 59.580 197.600 60.580 197.980 ;
        RECT 68.140 197.600 69.140 197.980 ;
        RECT 72.100 197.600 73.100 197.980 ;
        RECT 80.820 197.600 81.820 197.980 ;
        RECT 84.780 197.600 85.780 197.980 ;
        RECT 93.340 197.600 94.340 197.980 ;
        RECT 97.300 197.600 98.300 197.980 ;
        RECT 106.020 197.600 107.020 197.980 ;
        RECT 109.980 197.600 110.980 197.980 ;
        RECT 118.540 197.600 119.540 197.980 ;
        RECT 122.500 197.600 123.500 197.980 ;
        RECT 17.740 195.840 18.740 196.220 ;
        RECT 21.700 195.840 22.700 196.220 ;
        RECT 30.420 195.840 31.420 196.220 ;
        RECT 34.380 195.840 35.380 196.220 ;
        RECT 42.940 195.840 43.940 196.220 ;
        RECT 46.900 195.840 47.900 196.220 ;
        RECT 55.620 195.840 56.620 196.220 ;
        RECT 59.580 195.840 60.580 196.220 ;
        RECT 68.140 195.840 69.140 196.220 ;
        RECT 72.100 195.840 73.100 196.220 ;
        RECT 80.820 195.840 81.820 196.220 ;
        RECT 84.780 195.840 85.780 196.220 ;
        RECT 93.340 195.840 94.340 196.220 ;
        RECT 97.300 195.840 98.300 196.220 ;
        RECT 106.020 195.840 107.020 196.220 ;
        RECT 109.980 195.840 110.980 196.220 ;
        RECT 126.060 194.900 126.440 203.320 ;
        RECT 143.680 201.830 144.680 202.210 ;
        RECT 147.640 201.830 148.640 202.210 ;
        RECT 143.680 200.070 144.680 200.450 ;
        RECT 147.640 200.070 148.640 200.450 ;
        RECT 147.640 199.190 148.640 199.570 ;
        RECT 143.680 196.550 144.680 196.930 ;
        RECT 147.640 196.550 148.640 196.930 ;
        RECT 112.060 194.520 126.440 194.900 ;
        RECT 143.680 194.790 144.680 195.170 ;
        RECT 147.640 194.790 148.640 195.170 ;
        RECT 141.520 193.470 143.300 193.850 ;
        RECT 17.740 192.320 18.740 192.700 ;
        RECT 21.700 192.320 22.700 192.700 ;
        RECT 30.420 192.320 31.420 192.700 ;
        RECT 34.380 192.320 35.380 192.700 ;
        RECT 42.940 192.320 43.940 192.700 ;
        RECT 46.900 192.320 47.900 192.700 ;
        RECT 55.620 192.320 56.620 192.700 ;
        RECT 59.580 192.320 60.580 192.700 ;
        RECT 68.140 192.320 69.140 192.700 ;
        RECT 72.100 192.320 73.100 192.700 ;
        RECT 80.820 192.320 81.820 192.700 ;
        RECT 84.780 192.320 85.780 192.700 ;
        RECT 93.340 192.320 94.340 192.700 ;
        RECT 97.300 192.320 98.300 192.700 ;
        RECT 106.020 192.320 107.020 192.700 ;
        RECT 109.980 192.320 110.980 192.700 ;
        RECT 17.740 191.440 18.740 191.820 ;
        RECT 21.700 191.440 22.700 191.820 ;
        RECT 30.420 191.440 31.420 191.820 ;
        RECT 34.380 191.440 35.380 191.820 ;
        RECT 42.940 191.440 43.940 191.820 ;
        RECT 46.900 191.440 47.900 191.820 ;
        RECT 55.620 191.440 56.620 191.820 ;
        RECT 59.580 191.440 60.580 191.820 ;
        RECT 68.140 191.440 69.140 191.820 ;
        RECT 72.100 191.440 73.100 191.820 ;
        RECT 80.820 191.440 81.820 191.820 ;
        RECT 84.780 191.440 85.780 191.820 ;
        RECT 93.340 191.440 94.340 191.820 ;
        RECT 97.300 191.440 98.300 191.820 ;
        RECT 106.020 191.440 107.020 191.820 ;
        RECT 109.980 191.440 110.980 191.820 ;
        RECT 15.580 191.300 16.580 191.380 ;
        RECT 36.460 191.300 37.460 191.380 ;
        RECT 40.780 191.300 41.780 191.380 ;
        RECT 61.660 191.300 62.660 191.380 ;
        RECT 65.980 191.300 66.980 191.380 ;
        RECT 86.860 191.300 87.860 191.380 ;
        RECT 91.180 191.300 92.180 191.380 ;
        RECT 112.060 191.300 113.060 191.380 ;
        RECT 15.200 191.000 16.580 191.300 ;
        RECT 36.080 191.000 37.460 191.300 ;
        RECT 40.400 191.000 41.780 191.300 ;
        RECT 61.280 191.000 62.660 191.300 ;
        RECT 65.600 191.000 66.980 191.300 ;
        RECT 86.480 191.000 87.860 191.300 ;
        RECT 90.800 191.000 92.180 191.300 ;
        RECT 111.680 191.000 113.060 191.300 ;
        RECT 15.200 190.680 15.580 191.000 ;
        RECT 36.080 190.680 36.460 191.000 ;
        RECT 40.400 190.680 40.780 191.000 ;
        RECT 61.280 190.680 61.660 191.000 ;
        RECT 65.600 190.680 65.980 191.000 ;
        RECT 86.480 190.680 86.860 191.000 ;
        RECT 90.800 190.680 91.180 191.000 ;
        RECT 111.680 190.680 112.060 191.000 ;
        RECT 15.200 190.300 113.140 190.680 ;
        RECT 17.740 188.800 18.740 189.180 ;
        RECT 34.380 188.800 35.380 189.180 ;
        RECT 42.940 188.800 43.940 189.180 ;
        RECT 59.580 188.800 60.580 189.180 ;
        RECT 68.140 188.800 69.140 189.180 ;
        RECT 84.780 188.800 85.780 189.180 ;
        RECT 93.340 188.800 94.340 189.180 ;
        RECT 109.980 188.800 110.980 189.180 ;
        RECT 142.920 188.570 143.300 193.470 ;
        RECT 147.640 191.270 148.640 191.650 ;
        RECT 147.640 190.390 148.640 190.770 ;
        RECT 143.680 189.510 144.680 189.890 ;
        RECT 17.740 187.920 18.740 188.300 ;
        RECT 21.700 187.920 23.480 188.300 ;
        RECT 17.740 185.280 18.740 185.660 ;
        RECT 23.100 184.780 23.480 187.920 ;
        RECT 29.640 187.920 31.420 188.300 ;
        RECT 34.380 187.920 35.380 188.300 ;
        RECT 42.940 187.920 43.940 188.300 ;
        RECT 46.900 187.920 48.680 188.300 ;
        RECT 24.580 184.780 25.580 185.400 ;
        RECT 17.740 184.400 18.740 184.780 ;
        RECT 21.700 184.400 25.580 184.780 ;
        RECT 27.540 184.780 28.540 185.400 ;
        RECT 29.640 184.780 30.020 187.920 ;
        RECT 34.380 185.280 35.380 185.660 ;
        RECT 42.940 185.280 43.940 185.660 ;
        RECT 48.300 184.780 48.680 187.920 ;
        RECT 54.840 187.920 56.620 188.300 ;
        RECT 59.580 187.920 60.580 188.300 ;
        RECT 68.140 187.920 69.140 188.300 ;
        RECT 72.100 187.920 73.880 188.300 ;
        RECT 49.780 184.780 50.780 185.400 ;
        RECT 27.540 184.400 31.420 184.780 ;
        RECT 34.380 184.400 35.380 184.780 ;
        RECT 42.940 184.400 43.940 184.780 ;
        RECT 46.900 184.400 50.780 184.780 ;
        RECT 52.740 184.780 53.740 185.400 ;
        RECT 54.840 184.780 55.220 187.920 ;
        RECT 59.580 185.280 60.580 185.660 ;
        RECT 68.140 185.280 69.140 185.660 ;
        RECT 73.500 184.780 73.880 187.920 ;
        RECT 80.040 187.920 81.820 188.300 ;
        RECT 84.780 187.920 85.780 188.300 ;
        RECT 93.340 187.920 94.340 188.300 ;
        RECT 97.300 187.920 99.080 188.300 ;
        RECT 74.980 184.780 75.980 185.400 ;
        RECT 52.740 184.400 56.620 184.780 ;
        RECT 59.580 184.400 60.580 184.780 ;
        RECT 68.140 184.400 69.140 184.780 ;
        RECT 72.100 184.400 75.980 184.780 ;
        RECT 77.940 184.780 78.940 185.400 ;
        RECT 80.040 184.780 80.420 187.920 ;
        RECT 84.780 185.280 85.780 185.660 ;
        RECT 93.340 185.280 94.340 185.660 ;
        RECT 98.700 184.780 99.080 187.920 ;
        RECT 105.240 187.920 107.020 188.300 ;
        RECT 109.980 187.920 110.980 188.300 ;
        RECT 142.920 188.190 150.800 188.570 ;
        RECT 100.180 184.780 101.180 185.400 ;
        RECT 77.940 184.400 81.820 184.780 ;
        RECT 84.780 184.400 85.780 184.780 ;
        RECT 93.340 184.400 94.340 184.780 ;
        RECT 97.300 184.400 101.180 184.780 ;
        RECT 103.140 184.780 104.140 185.400 ;
        RECT 105.240 184.780 105.620 187.920 ;
        RECT 122.500 186.160 123.500 186.540 ;
        RECT 143.680 185.990 144.680 186.370 ;
        RECT 147.640 185.990 148.640 186.370 ;
        RECT 109.980 185.280 110.980 185.660 ;
        RECT 118.540 185.280 119.540 185.660 ;
        RECT 103.140 184.400 107.020 184.780 ;
        RECT 109.980 184.400 110.980 184.780 ;
        RECT 122.500 184.400 123.500 184.780 ;
        RECT 20.910 182.290 21.290 183.290 ;
        RECT 23.100 182.140 23.480 184.400 ;
        RECT 17.740 181.760 18.740 182.140 ;
        RECT 21.700 181.760 23.480 182.140 ;
        RECT 29.640 182.140 30.020 184.400 ;
        RECT 31.830 182.290 32.210 183.290 ;
        RECT 46.110 182.290 46.490 183.290 ;
        RECT 48.300 182.140 48.680 184.400 ;
        RECT 29.640 181.760 31.420 182.140 ;
        RECT 34.380 181.760 35.380 182.140 ;
        RECT 42.940 181.760 43.940 182.140 ;
        RECT 46.900 181.760 48.680 182.140 ;
        RECT 54.840 182.140 55.220 184.400 ;
        RECT 57.030 182.290 57.410 183.290 ;
        RECT 71.310 182.290 71.690 183.290 ;
        RECT 73.500 182.140 73.880 184.400 ;
        RECT 54.840 181.760 56.620 182.140 ;
        RECT 59.580 181.760 60.580 182.140 ;
        RECT 68.140 181.760 69.140 182.140 ;
        RECT 72.100 181.760 73.880 182.140 ;
        RECT 80.040 182.140 80.420 184.400 ;
        RECT 82.230 182.290 82.610 183.290 ;
        RECT 96.510 182.290 96.890 183.290 ;
        RECT 98.700 182.140 99.080 184.400 ;
        RECT 80.040 181.760 81.820 182.140 ;
        RECT 84.780 181.760 85.780 182.140 ;
        RECT 93.340 181.760 94.340 182.140 ;
        RECT 97.300 181.760 99.080 182.140 ;
        RECT 105.240 182.140 105.620 184.400 ;
        RECT 143.680 184.230 144.680 184.610 ;
        RECT 147.640 184.230 148.640 184.610 ;
        RECT 107.430 182.290 107.810 183.290 ;
        RECT 116.380 182.200 118.160 182.580 ;
        RECT 105.240 181.760 107.020 182.140 ;
        RECT 109.980 181.760 110.980 182.140 ;
        RECT 122.500 181.760 123.500 182.140 ;
        RECT 17.740 180.880 18.740 181.260 ;
        RECT 21.700 180.880 23.480 181.260 ;
        RECT 17.740 178.240 18.740 178.620 ;
        RECT 23.100 177.740 23.480 180.880 ;
        RECT 29.640 180.880 31.420 181.260 ;
        RECT 34.380 180.880 35.380 181.260 ;
        RECT 42.940 180.880 43.940 181.260 ;
        RECT 46.900 180.880 48.680 181.260 ;
        RECT 24.580 177.740 25.580 178.360 ;
        RECT 17.740 177.360 18.740 177.740 ;
        RECT 21.700 177.360 25.580 177.740 ;
        RECT 27.540 177.740 28.540 178.360 ;
        RECT 29.640 177.740 30.020 180.880 ;
        RECT 34.380 178.240 35.380 178.620 ;
        RECT 42.940 178.240 43.940 178.620 ;
        RECT 48.300 177.740 48.680 180.880 ;
        RECT 54.840 180.880 56.620 181.260 ;
        RECT 59.580 180.880 60.580 181.260 ;
        RECT 68.140 180.880 69.140 181.260 ;
        RECT 72.100 180.880 73.880 181.260 ;
        RECT 49.780 177.740 50.780 178.360 ;
        RECT 27.540 177.360 31.420 177.740 ;
        RECT 34.380 177.360 35.380 177.740 ;
        RECT 42.940 177.360 43.940 177.740 ;
        RECT 46.900 177.360 50.780 177.740 ;
        RECT 52.740 177.740 53.740 178.360 ;
        RECT 54.840 177.740 55.220 180.880 ;
        RECT 59.580 178.240 60.580 178.620 ;
        RECT 68.140 178.240 69.140 178.620 ;
        RECT 73.500 177.740 73.880 180.880 ;
        RECT 80.040 180.880 81.820 181.260 ;
        RECT 84.780 180.880 85.780 181.260 ;
        RECT 93.340 180.880 94.340 181.260 ;
        RECT 97.300 180.880 99.080 181.260 ;
        RECT 74.980 177.740 75.980 178.360 ;
        RECT 52.740 177.360 56.620 177.740 ;
        RECT 59.580 177.360 60.580 177.740 ;
        RECT 68.140 177.360 69.140 177.740 ;
        RECT 72.100 177.360 75.980 177.740 ;
        RECT 77.940 177.740 78.940 178.360 ;
        RECT 80.040 177.740 80.420 180.880 ;
        RECT 84.780 178.240 85.780 178.620 ;
        RECT 93.340 178.240 94.340 178.620 ;
        RECT 98.700 177.740 99.080 180.880 ;
        RECT 105.240 180.880 107.020 181.260 ;
        RECT 109.980 180.880 110.980 181.260 ;
        RECT 122.500 180.880 123.500 181.260 ;
        RECT 100.180 177.740 101.180 178.360 ;
        RECT 77.940 177.360 81.820 177.740 ;
        RECT 84.780 177.360 85.780 177.740 ;
        RECT 93.340 177.360 94.340 177.740 ;
        RECT 97.300 177.360 101.180 177.740 ;
        RECT 103.140 177.740 104.140 178.360 ;
        RECT 105.240 177.740 105.620 180.880 ;
        RECT 143.680 180.710 144.680 181.090 ;
        RECT 147.640 180.710 148.640 181.090 ;
        RECT 109.980 178.240 110.980 178.620 ;
        RECT 122.500 178.240 123.500 178.620 ;
        RECT 103.140 177.360 107.020 177.740 ;
        RECT 109.980 177.360 110.980 177.740 ;
        RECT 122.500 177.360 123.500 177.740 ;
        RECT 20.035 175.250 20.415 176.250 ;
        RECT 23.100 175.100 23.480 177.360 ;
        RECT 17.740 174.720 18.740 175.100 ;
        RECT 21.700 174.720 23.480 175.100 ;
        RECT 29.640 175.100 30.020 177.360 ;
        RECT 32.705 175.250 33.085 176.250 ;
        RECT 45.235 175.250 45.615 176.250 ;
        RECT 48.300 175.100 48.680 177.360 ;
        RECT 29.640 174.720 31.420 175.100 ;
        RECT 34.380 174.720 35.380 175.100 ;
        RECT 42.940 174.720 43.940 175.100 ;
        RECT 46.900 174.720 48.680 175.100 ;
        RECT 54.840 175.100 55.220 177.360 ;
        RECT 57.905 175.250 58.285 176.250 ;
        RECT 70.435 175.250 70.815 176.250 ;
        RECT 73.500 175.100 73.880 177.360 ;
        RECT 54.840 174.720 56.620 175.100 ;
        RECT 59.580 174.720 60.580 175.100 ;
        RECT 68.140 174.720 69.140 175.100 ;
        RECT 72.100 174.720 73.880 175.100 ;
        RECT 80.040 175.100 80.420 177.360 ;
        RECT 83.105 175.250 83.485 176.250 ;
        RECT 95.635 175.250 96.015 176.250 ;
        RECT 98.700 175.100 99.080 177.360 ;
        RECT 80.040 174.720 81.820 175.100 ;
        RECT 84.780 174.720 85.780 175.100 ;
        RECT 93.340 174.720 94.340 175.100 ;
        RECT 97.300 174.720 99.080 175.100 ;
        RECT 105.240 175.100 105.620 177.360 ;
        RECT 124.660 176.920 125.660 177.300 ;
        RECT 143.680 177.190 144.680 177.570 ;
        RECT 147.640 177.190 148.640 177.570 ;
        RECT 108.305 175.250 108.685 176.250 ;
        RECT 143.680 175.430 144.680 175.810 ;
        RECT 147.640 175.430 148.640 175.810 ;
        RECT 105.240 174.720 107.020 175.100 ;
        RECT 109.980 174.720 110.980 175.100 ;
        RECT 122.500 174.720 123.500 175.100 ;
        RECT 147.640 174.550 148.640 174.930 ;
        RECT 17.740 173.840 18.740 174.220 ;
        RECT 21.700 173.840 23.480 174.220 ;
        RECT 17.740 171.200 18.740 171.580 ;
        RECT 23.100 170.700 23.480 173.840 ;
        RECT 29.640 173.840 31.420 174.220 ;
        RECT 34.380 173.840 35.380 174.220 ;
        RECT 42.940 173.840 43.940 174.220 ;
        RECT 46.900 173.840 48.680 174.220 ;
        RECT 24.580 170.700 25.580 171.320 ;
        RECT 17.740 170.320 18.740 170.700 ;
        RECT 21.700 170.320 25.580 170.700 ;
        RECT 27.540 170.700 28.540 171.320 ;
        RECT 29.640 170.700 30.020 173.840 ;
        RECT 34.380 171.200 35.380 171.580 ;
        RECT 42.940 171.200 43.940 171.580 ;
        RECT 48.300 170.700 48.680 173.840 ;
        RECT 54.840 173.840 56.620 174.220 ;
        RECT 59.580 173.840 60.580 174.220 ;
        RECT 68.140 173.840 69.140 174.220 ;
        RECT 72.100 173.840 73.880 174.220 ;
        RECT 49.780 170.700 50.780 171.320 ;
        RECT 27.540 170.320 31.420 170.700 ;
        RECT 34.380 170.320 35.380 170.700 ;
        RECT 42.940 170.320 43.940 170.700 ;
        RECT 46.900 170.320 50.780 170.700 ;
        RECT 52.740 170.700 53.740 171.320 ;
        RECT 54.840 170.700 55.220 173.840 ;
        RECT 59.580 171.200 60.580 171.580 ;
        RECT 68.140 171.200 69.140 171.580 ;
        RECT 73.500 170.700 73.880 173.840 ;
        RECT 80.040 173.840 81.820 174.220 ;
        RECT 84.780 173.840 85.780 174.220 ;
        RECT 93.340 173.840 94.340 174.220 ;
        RECT 97.300 173.840 99.080 174.220 ;
        RECT 74.980 170.700 75.980 171.320 ;
        RECT 52.740 170.320 56.620 170.700 ;
        RECT 59.580 170.320 60.580 170.700 ;
        RECT 68.140 170.320 69.140 170.700 ;
        RECT 72.100 170.320 75.980 170.700 ;
        RECT 77.940 170.700 78.940 171.320 ;
        RECT 80.040 170.700 80.420 173.840 ;
        RECT 84.780 171.200 85.780 171.580 ;
        RECT 93.340 171.200 94.340 171.580 ;
        RECT 98.700 170.700 99.080 173.840 ;
        RECT 105.240 173.840 107.020 174.220 ;
        RECT 109.980 173.840 110.980 174.220 ;
        RECT 122.500 173.840 123.500 174.220 ;
        RECT 100.180 170.700 101.180 171.320 ;
        RECT 77.940 170.320 81.820 170.700 ;
        RECT 84.780 170.320 85.780 170.700 ;
        RECT 93.340 170.320 94.340 170.700 ;
        RECT 97.300 170.320 101.180 170.700 ;
        RECT 103.140 170.700 104.140 171.320 ;
        RECT 105.240 170.700 105.620 173.840 ;
        RECT 118.540 172.960 119.540 173.340 ;
        RECT 118.540 172.080 119.540 172.460 ;
        RECT 122.500 172.080 123.500 172.460 ;
        RECT 143.680 171.910 144.680 172.290 ;
        RECT 147.640 171.910 148.640 172.290 ;
        RECT 109.980 171.200 110.980 171.580 ;
        RECT 113.460 170.700 122.800 171.080 ;
        RECT 103.140 170.320 107.020 170.700 ;
        RECT 109.980 170.320 110.980 170.700 ;
        RECT 15.660 168.080 16.660 168.460 ;
        RECT 19.235 168.210 19.615 169.210 ;
        RECT 23.100 168.060 23.480 170.320 ;
        RECT 17.740 167.680 18.740 168.060 ;
        RECT 21.700 167.680 23.480 168.060 ;
        RECT 29.640 168.060 30.020 170.320 ;
        RECT 33.505 168.210 33.885 169.210 ;
        RECT 36.460 168.080 37.460 168.460 ;
        RECT 40.860 168.080 41.860 168.460 ;
        RECT 44.435 168.210 44.815 169.210 ;
        RECT 48.300 168.060 48.680 170.320 ;
        RECT 29.640 167.680 31.420 168.060 ;
        RECT 34.380 167.680 35.380 168.060 ;
        RECT 42.940 167.680 43.940 168.060 ;
        RECT 46.900 167.680 48.680 168.060 ;
        RECT 54.840 168.060 55.220 170.320 ;
        RECT 58.705 168.210 59.085 169.210 ;
        RECT 61.660 168.080 62.660 168.460 ;
        RECT 66.060 168.080 67.060 168.460 ;
        RECT 69.635 168.210 70.015 169.210 ;
        RECT 73.500 168.060 73.880 170.320 ;
        RECT 54.840 167.680 56.620 168.060 ;
        RECT 59.580 167.680 60.580 168.060 ;
        RECT 68.140 167.680 69.140 168.060 ;
        RECT 72.100 167.680 73.880 168.060 ;
        RECT 80.040 168.060 80.420 170.320 ;
        RECT 83.905 168.210 84.285 169.210 ;
        RECT 86.860 168.080 87.860 168.460 ;
        RECT 91.260 168.080 92.260 168.460 ;
        RECT 94.835 168.210 95.215 169.210 ;
        RECT 98.700 168.060 99.080 170.320 ;
        RECT 80.040 167.680 81.820 168.060 ;
        RECT 84.780 167.680 85.780 168.060 ;
        RECT 93.340 167.680 94.340 168.060 ;
        RECT 97.300 167.680 99.080 168.060 ;
        RECT 105.240 168.060 105.620 170.320 ;
        RECT 109.105 168.210 109.485 169.210 ;
        RECT 112.060 168.080 113.060 168.460 ;
        RECT 105.240 167.680 107.020 168.060 ;
        RECT 109.980 167.680 110.980 168.060 ;
        RECT 17.740 166.800 18.740 167.180 ;
        RECT 21.700 166.800 23.480 167.180 ;
        RECT 17.740 164.160 18.740 164.540 ;
        RECT 23.100 163.660 23.480 166.800 ;
        RECT 29.640 166.800 31.420 167.180 ;
        RECT 34.380 166.800 35.380 167.180 ;
        RECT 42.940 166.800 43.940 167.180 ;
        RECT 46.900 166.800 48.680 167.180 ;
        RECT 24.580 163.660 25.580 164.280 ;
        RECT 17.740 163.280 18.740 163.660 ;
        RECT 21.700 163.280 25.580 163.660 ;
        RECT 27.540 163.660 28.540 164.280 ;
        RECT 29.640 163.660 30.020 166.800 ;
        RECT 34.380 164.160 35.380 164.540 ;
        RECT 42.940 164.160 43.940 164.540 ;
        RECT 48.300 163.660 48.680 166.800 ;
        RECT 54.840 166.800 56.620 167.180 ;
        RECT 59.580 166.800 60.580 167.180 ;
        RECT 68.140 166.800 69.140 167.180 ;
        RECT 72.100 166.800 73.880 167.180 ;
        RECT 49.780 163.660 50.780 164.280 ;
        RECT 27.540 163.280 31.420 163.660 ;
        RECT 34.380 163.280 35.380 163.660 ;
        RECT 42.940 163.280 43.940 163.660 ;
        RECT 46.900 163.280 50.780 163.660 ;
        RECT 52.740 163.660 53.740 164.280 ;
        RECT 54.840 163.660 55.220 166.800 ;
        RECT 59.580 164.160 60.580 164.540 ;
        RECT 68.140 164.160 69.140 164.540 ;
        RECT 73.500 163.660 73.880 166.800 ;
        RECT 80.040 166.800 81.820 167.180 ;
        RECT 84.780 166.800 85.780 167.180 ;
        RECT 93.340 166.800 94.340 167.180 ;
        RECT 97.300 166.800 99.080 167.180 ;
        RECT 74.980 163.660 75.980 164.280 ;
        RECT 52.740 163.280 56.620 163.660 ;
        RECT 59.580 163.280 60.580 163.660 ;
        RECT 68.140 163.280 69.140 163.660 ;
        RECT 72.100 163.280 75.980 163.660 ;
        RECT 77.940 163.660 78.940 164.280 ;
        RECT 80.040 163.660 80.420 166.800 ;
        RECT 84.780 164.160 85.780 164.540 ;
        RECT 93.340 164.160 94.340 164.540 ;
        RECT 98.700 163.660 99.080 166.800 ;
        RECT 105.240 166.800 107.020 167.180 ;
        RECT 109.980 166.800 110.980 167.180 ;
        RECT 100.180 163.660 101.180 164.280 ;
        RECT 77.940 163.280 81.820 163.660 ;
        RECT 84.780 163.280 85.780 163.660 ;
        RECT 93.340 163.280 94.340 163.660 ;
        RECT 97.300 163.280 101.180 163.660 ;
        RECT 103.140 163.660 104.140 164.280 ;
        RECT 105.240 163.660 105.620 166.800 ;
        RECT 109.980 164.160 110.980 164.540 ;
        RECT 103.140 163.280 107.020 163.660 ;
        RECT 109.980 163.280 110.980 163.660 ;
        RECT 23.100 161.020 23.480 163.280 ;
        RECT 17.740 160.640 18.740 161.020 ;
        RECT 21.700 160.640 23.480 161.020 ;
        RECT 29.640 161.020 30.020 163.280 ;
        RECT 48.300 161.020 48.680 163.280 ;
        RECT 29.640 160.640 31.420 161.020 ;
        RECT 34.380 160.640 35.380 161.020 ;
        RECT 42.940 160.640 43.940 161.020 ;
        RECT 46.900 160.640 48.680 161.020 ;
        RECT 54.840 161.020 55.220 163.280 ;
        RECT 73.500 161.020 73.880 163.280 ;
        RECT 54.840 160.640 56.620 161.020 ;
        RECT 59.580 160.640 60.580 161.020 ;
        RECT 68.140 160.640 69.140 161.020 ;
        RECT 72.100 160.640 73.880 161.020 ;
        RECT 80.040 161.020 80.420 163.280 ;
        RECT 98.700 161.020 99.080 163.280 ;
        RECT 80.040 160.640 81.820 161.020 ;
        RECT 84.780 160.640 85.780 161.020 ;
        RECT 93.340 160.640 94.340 161.020 ;
        RECT 97.300 160.640 99.080 161.020 ;
        RECT 105.240 161.020 105.620 163.280 ;
        RECT 105.240 160.640 107.020 161.020 ;
        RECT 109.980 160.640 110.980 161.020 ;
        RECT 15.580 159.620 16.580 159.700 ;
        RECT 23.860 159.620 24.860 159.700 ;
        RECT 28.180 159.620 29.180 159.700 ;
        RECT 49.060 159.620 50.060 159.700 ;
        RECT 53.380 159.620 54.380 159.700 ;
        RECT 74.260 159.620 75.260 159.700 ;
        RECT 78.580 159.620 79.580 159.700 ;
        RECT 99.460 159.620 100.460 159.700 ;
        RECT 103.780 159.620 104.780 159.700 ;
        RECT 15.580 159.320 104.860 159.620 ;
        RECT 113.460 156.180 113.840 170.700 ;
        RECT 122.500 170.320 123.500 170.700 ;
        RECT 143.680 170.150 144.680 170.530 ;
        RECT 147.640 170.150 148.640 170.530 ;
        RECT 118.540 169.440 119.540 169.820 ;
        RECT 122.500 169.440 123.500 169.820 ;
        RECT 118.540 168.560 119.540 168.940 ;
        RECT 122.500 168.560 123.500 168.940 ;
        RECT 141.520 168.830 143.300 169.210 ;
        RECT 118.620 167.330 119.620 167.370 ;
        RECT 15.580 156.100 16.580 156.180 ;
        RECT 36.460 156.100 37.460 156.180 ;
        RECT 40.780 156.100 41.780 156.180 ;
        RECT 61.660 156.100 62.660 156.180 ;
        RECT 65.980 156.100 66.980 156.180 ;
        RECT 86.860 156.100 87.860 156.180 ;
        RECT 91.180 156.100 92.180 156.180 ;
        RECT 112.060 156.100 113.840 156.180 ;
        RECT 15.200 155.800 16.580 156.100 ;
        RECT 36.080 155.800 37.460 156.100 ;
        RECT 40.400 155.800 41.780 156.100 ;
        RECT 61.280 155.800 62.660 156.100 ;
        RECT 65.600 155.800 66.980 156.100 ;
        RECT 86.480 155.800 87.860 156.100 ;
        RECT 90.800 155.800 92.180 156.100 ;
        RECT 111.680 155.800 113.840 156.100 ;
        RECT 115.720 166.990 119.620 167.330 ;
        RECT 115.720 166.950 119.080 166.990 ;
        RECT 15.200 154.720 15.580 155.800 ;
        RECT 17.740 155.360 18.740 155.740 ;
        RECT 21.700 155.360 22.700 155.740 ;
        RECT 30.420 155.360 31.420 155.740 ;
        RECT 34.380 155.360 35.380 155.740 ;
        RECT 36.080 154.720 36.460 155.800 ;
        RECT 40.400 154.720 40.780 155.800 ;
        RECT 42.940 155.360 43.940 155.740 ;
        RECT 46.900 155.360 47.900 155.740 ;
        RECT 55.620 155.360 56.620 155.740 ;
        RECT 59.580 155.360 60.580 155.740 ;
        RECT 61.280 154.720 61.660 155.800 ;
        RECT 65.600 154.720 65.980 155.800 ;
        RECT 68.140 155.360 69.140 155.740 ;
        RECT 72.100 155.360 73.100 155.740 ;
        RECT 80.820 155.360 81.820 155.740 ;
        RECT 84.780 155.360 85.780 155.740 ;
        RECT 86.480 154.720 86.860 155.800 ;
        RECT 90.800 154.720 91.180 155.800 ;
        RECT 93.340 155.360 94.340 155.740 ;
        RECT 97.300 155.360 98.300 155.740 ;
        RECT 106.020 155.360 107.020 155.740 ;
        RECT 109.980 155.360 110.980 155.740 ;
        RECT 111.680 154.720 112.060 155.800 ;
        RECT 15.200 154.340 113.140 154.720 ;
        RECT 15.280 151.940 113.060 152.320 ;
        RECT 15.280 150.860 15.660 151.940 ;
        RECT 36.080 150.860 36.460 151.940 ;
        RECT 40.480 150.860 40.860 151.940 ;
        RECT 61.280 150.860 61.660 151.940 ;
        RECT 65.680 150.860 66.060 151.940 ;
        RECT 86.480 150.860 86.860 151.940 ;
        RECT 90.880 150.860 91.260 151.940 ;
        RECT 111.680 150.860 112.060 151.940 ;
        RECT 115.720 151.240 116.100 166.950 ;
        RECT 118.540 165.920 119.540 166.300 ;
        RECT 122.500 165.920 123.500 166.300 ;
        RECT 122.500 165.040 123.500 165.420 ;
        RECT 142.920 163.930 143.300 168.830 ;
        RECT 147.640 166.630 148.640 167.010 ;
        RECT 147.640 165.750 148.640 166.130 ;
        RECT 143.680 164.870 144.680 165.250 ;
        RECT 142.920 163.550 150.800 163.930 ;
        RECT 122.500 162.400 123.500 162.780 ;
        RECT 122.500 161.520 123.500 161.900 ;
        RECT 143.680 161.350 144.680 161.730 ;
        RECT 147.640 161.350 148.640 161.730 ;
        RECT 143.680 159.590 144.680 159.970 ;
        RECT 147.640 159.590 148.640 159.970 ;
        RECT 122.500 158.880 123.500 159.260 ;
        RECT 122.500 158.000 123.500 158.380 ;
        RECT 124.660 157.560 125.660 157.940 ;
        RECT 143.680 156.070 144.680 156.450 ;
        RECT 147.640 156.070 148.640 156.450 ;
        RECT 122.500 155.360 123.500 155.740 ;
        RECT 122.500 154.480 123.500 154.860 ;
        RECT 118.540 153.600 119.540 153.980 ;
        RECT 143.680 152.550 144.680 152.930 ;
        RECT 147.640 152.550 148.640 152.930 ;
        RECT 112.760 150.860 116.100 151.240 ;
        RECT 15.280 150.480 16.660 150.860 ;
        RECT 36.080 150.480 37.460 150.860 ;
        RECT 40.480 150.480 41.860 150.860 ;
        RECT 61.280 150.480 62.660 150.860 ;
        RECT 65.680 150.480 67.060 150.860 ;
        RECT 86.480 150.480 87.860 150.860 ;
        RECT 90.880 150.480 92.260 150.860 ;
        RECT 111.680 150.480 113.060 150.860 ;
        RECT 116.380 150.520 117.380 150.900 ;
        RECT 143.680 150.790 144.680 151.170 ;
        RECT 147.640 150.790 148.640 151.170 ;
        RECT 17.740 150.080 18.740 150.460 ;
        RECT 21.700 150.080 22.700 150.460 ;
        RECT 30.420 150.080 31.420 150.460 ;
        RECT 34.380 150.080 35.380 150.460 ;
        RECT 42.940 150.080 43.940 150.460 ;
        RECT 46.900 150.080 47.900 150.460 ;
        RECT 55.620 150.080 56.620 150.460 ;
        RECT 59.580 150.080 60.580 150.460 ;
        RECT 68.140 150.080 69.140 150.460 ;
        RECT 72.100 150.080 73.100 150.460 ;
        RECT 80.820 150.080 81.820 150.460 ;
        RECT 84.780 150.080 85.780 150.460 ;
        RECT 93.340 150.080 94.340 150.460 ;
        RECT 97.300 150.080 98.300 150.460 ;
        RECT 106.020 150.080 107.020 150.460 ;
        RECT 109.980 150.080 110.980 150.460 ;
        RECT 147.640 149.910 148.640 150.290 ;
        RECT 17.740 148.320 18.740 148.700 ;
        RECT 21.700 148.320 22.700 148.700 ;
        RECT 30.420 148.320 31.420 148.700 ;
        RECT 34.380 148.320 35.380 148.700 ;
        RECT 42.940 148.320 43.940 148.700 ;
        RECT 46.900 148.320 47.900 148.700 ;
        RECT 55.620 148.320 56.620 148.700 ;
        RECT 59.580 148.320 60.580 148.700 ;
        RECT 68.140 148.320 69.140 148.700 ;
        RECT 72.100 148.320 73.100 148.700 ;
        RECT 80.820 148.320 81.820 148.700 ;
        RECT 84.780 148.320 85.780 148.700 ;
        RECT 93.340 148.320 94.340 148.700 ;
        RECT 97.300 148.320 98.300 148.700 ;
        RECT 106.020 148.320 107.020 148.700 ;
        RECT 109.980 148.320 110.980 148.700 ;
        RECT 21.700 147.440 22.700 147.820 ;
        RECT 30.420 147.440 31.420 147.820 ;
        RECT 46.900 147.440 47.900 147.820 ;
        RECT 55.620 147.440 56.620 147.820 ;
        RECT 72.100 147.440 73.100 147.820 ;
        RECT 80.820 147.440 81.820 147.820 ;
        RECT 97.300 147.440 98.300 147.820 ;
        RECT 106.020 147.440 107.020 147.820 ;
        RECT 143.680 147.270 144.680 147.650 ;
        RECT 147.640 147.270 148.640 147.650 ;
        RECT 17.740 146.560 18.740 146.940 ;
        RECT 34.380 146.560 35.380 146.940 ;
        RECT 42.940 146.560 43.940 146.940 ;
        RECT 59.580 146.560 60.580 146.940 ;
        RECT 68.140 146.560 69.140 146.940 ;
        RECT 84.780 146.560 85.780 146.940 ;
        RECT 93.340 146.560 94.340 146.940 ;
        RECT 109.980 146.560 110.980 146.940 ;
        RECT 17.740 145.680 18.740 146.060 ;
        RECT 34.380 145.680 35.380 146.060 ;
        RECT 42.940 145.680 43.940 146.060 ;
        RECT 59.580 145.680 60.580 146.060 ;
        RECT 68.140 145.680 69.140 146.060 ;
        RECT 84.780 145.680 85.780 146.060 ;
        RECT 93.340 145.680 94.340 146.060 ;
        RECT 109.980 145.680 110.980 146.060 ;
        RECT 143.680 145.510 144.680 145.890 ;
        RECT 147.640 145.510 148.640 145.890 ;
        RECT 141.520 144.190 143.300 144.570 ;
        RECT 31.980 143.700 40.860 144.080 ;
        RECT 17.740 143.040 18.740 143.420 ;
        RECT 31.980 143.380 32.360 143.700 ;
        RECT 21.780 143.000 23.800 143.380 ;
        RECT 30.340 143.000 32.360 143.380 ;
        RECT 34.380 143.040 35.380 143.420 ;
        RECT 21.700 142.160 22.700 142.540 ;
        RECT 15.660 141.680 16.660 142.060 ;
        RECT 23.420 141.360 23.800 143.000 ;
        RECT 30.420 142.160 31.420 142.540 ;
        RECT 40.480 142.060 40.860 143.700 ;
        RECT 57.180 143.700 66.060 144.080 ;
        RECT 42.940 143.040 43.940 143.420 ;
        RECT 57.180 143.380 57.560 143.700 ;
        RECT 46.980 143.000 49.000 143.380 ;
        RECT 55.540 143.000 57.560 143.380 ;
        RECT 59.580 143.040 60.580 143.420 ;
        RECT 46.900 142.160 47.900 142.540 ;
        RECT 36.080 141.680 37.460 142.060 ;
        RECT 40.480 141.680 41.860 142.060 ;
        RECT 36.080 141.360 36.460 141.680 ;
        RECT 23.420 140.980 36.460 141.360 ;
        RECT 48.620 141.360 49.000 143.000 ;
        RECT 55.620 142.160 56.620 142.540 ;
        RECT 65.680 142.060 66.060 143.700 ;
        RECT 82.380 143.700 91.260 144.080 ;
        RECT 68.140 143.040 69.140 143.420 ;
        RECT 82.380 143.380 82.760 143.700 ;
        RECT 72.180 143.000 74.200 143.380 ;
        RECT 80.740 143.000 82.760 143.380 ;
        RECT 84.780 143.040 85.780 143.420 ;
        RECT 72.100 142.160 73.100 142.540 ;
        RECT 61.280 141.680 62.660 142.060 ;
        RECT 65.680 141.680 67.060 142.060 ;
        RECT 61.280 141.360 61.660 141.680 ;
        RECT 48.620 140.980 61.660 141.360 ;
        RECT 73.820 141.360 74.200 143.000 ;
        RECT 80.820 142.160 81.820 142.540 ;
        RECT 90.880 142.060 91.260 143.700 ;
        RECT 93.340 143.040 94.340 143.420 ;
        RECT 107.580 143.380 107.960 143.700 ;
        RECT 97.380 143.000 99.400 143.380 ;
        RECT 105.940 143.000 107.960 143.380 ;
        RECT 109.980 143.040 110.980 143.420 ;
        RECT 97.300 142.160 98.300 142.540 ;
        RECT 86.480 141.680 87.860 142.060 ;
        RECT 90.880 141.680 92.260 142.060 ;
        RECT 86.480 141.360 86.860 141.680 ;
        RECT 73.820 140.980 86.860 141.360 ;
        RECT 99.020 141.360 99.400 143.000 ;
        RECT 106.020 142.160 107.020 142.540 ;
        RECT 122.500 142.160 123.500 142.540 ;
        RECT 111.680 141.680 113.060 142.060 ;
        RECT 111.680 141.360 112.060 141.680 ;
        RECT 99.020 140.980 112.060 141.360 ;
        RECT 118.540 141.280 119.540 141.660 ;
        RECT 17.740 140.400 18.740 140.780 ;
        RECT 21.700 140.400 22.700 140.780 ;
        RECT 30.420 140.400 31.420 140.780 ;
        RECT 34.380 140.400 35.380 140.780 ;
        RECT 42.940 140.400 43.940 140.780 ;
        RECT 46.900 140.400 47.900 140.780 ;
        RECT 55.620 140.400 56.620 140.780 ;
        RECT 59.580 140.400 60.580 140.780 ;
        RECT 68.140 140.400 69.140 140.780 ;
        RECT 72.100 140.400 73.100 140.780 ;
        RECT 80.820 140.400 81.820 140.780 ;
        RECT 84.780 140.400 85.780 140.780 ;
        RECT 93.340 140.400 94.340 140.780 ;
        RECT 97.300 140.400 98.300 140.780 ;
        RECT 106.020 140.400 107.020 140.780 ;
        RECT 109.980 140.400 110.980 140.780 ;
        RECT 118.540 140.400 119.540 140.780 ;
        RECT 122.500 140.400 123.500 140.780 ;
        RECT 17.740 139.520 18.740 139.900 ;
        RECT 21.700 139.520 22.700 139.900 ;
        RECT 30.420 139.520 31.420 139.900 ;
        RECT 34.380 139.520 35.380 139.900 ;
        RECT 42.940 139.520 43.940 139.900 ;
        RECT 46.900 139.520 47.900 139.900 ;
        RECT 55.620 139.520 56.620 139.900 ;
        RECT 59.580 139.520 60.580 139.900 ;
        RECT 68.140 139.520 69.140 139.900 ;
        RECT 72.100 139.520 73.100 139.900 ;
        RECT 80.820 139.520 81.820 139.900 ;
        RECT 84.780 139.520 85.780 139.900 ;
        RECT 93.340 139.520 94.340 139.900 ;
        RECT 97.300 139.520 98.300 139.900 ;
        RECT 106.020 139.520 107.020 139.900 ;
        RECT 109.980 139.520 110.980 139.900 ;
        RECT 118.540 139.520 119.540 139.900 ;
        RECT 122.500 139.520 123.500 139.900 ;
        RECT 142.920 139.290 143.300 144.190 ;
        RECT 147.640 141.990 148.640 142.370 ;
        RECT 147.640 141.110 148.640 141.490 ;
        RECT 143.680 140.230 144.680 140.610 ;
        RECT 142.920 138.910 150.800 139.290 ;
        RECT 143.680 136.710 144.680 137.090 ;
        RECT 147.640 136.710 148.640 137.090 ;
        RECT 72.020 135.730 72.400 136.040 ;
        RECT 96.510 135.730 96.890 136.040 ;
        RECT 72.020 135.350 96.890 135.730 ;
        RECT 72.020 135.040 72.400 135.350 ;
        RECT 72.920 134.760 73.300 135.070 ;
        RECT 82.230 134.760 82.610 135.070 ;
        RECT 96.510 135.040 96.890 135.350 ;
        RECT 143.680 134.950 144.680 135.330 ;
        RECT 147.640 134.950 148.640 135.330 ;
        RECT 72.920 134.380 82.610 134.760 ;
        RECT 71.310 133.790 71.690 134.100 ;
        RECT 72.920 134.070 73.300 134.380 ;
        RECT 73.820 133.790 74.200 134.100 ;
        RECT 82.230 134.070 82.610 134.380 ;
        RECT 71.310 133.410 74.240 133.790 ;
        RECT 57.030 132.820 57.410 133.130 ;
        RECT 71.310 133.100 71.690 133.410 ;
        RECT 73.820 133.100 74.200 133.410 ;
        RECT 74.720 132.820 75.100 133.130 ;
        RECT 57.030 132.440 75.140 132.820 ;
        RECT 46.110 131.850 46.490 132.160 ;
        RECT 57.030 132.130 57.410 132.440 ;
        RECT 74.720 132.130 75.100 132.440 ;
        RECT 75.620 131.850 76.000 132.160 ;
        RECT 46.110 131.470 76.040 131.850 ;
        RECT 31.830 130.880 32.210 131.190 ;
        RECT 46.110 131.160 46.490 131.470 ;
        RECT 75.620 131.160 76.000 131.470 ;
        RECT 143.680 131.430 144.680 131.810 ;
        RECT 147.640 131.430 148.640 131.810 ;
        RECT 77.420 130.880 77.800 131.190 ;
        RECT 31.830 130.500 77.840 130.880 ;
        RECT 20.910 129.910 21.290 130.220 ;
        RECT 31.830 130.190 32.210 130.500 ;
        RECT 77.420 130.190 77.800 130.500 ;
        RECT 79.220 129.910 79.600 130.220 ;
        RECT 20.910 129.530 79.640 129.910 ;
        RECT 20.910 129.220 21.290 129.530 ;
        RECT 45.235 128.940 45.615 129.250 ;
        RECT 65.120 128.940 65.500 129.250 ;
        RECT 79.220 129.220 79.600 129.530 ;
        RECT 45.235 128.560 65.540 128.940 ;
        RECT 32.700 127.970 33.080 128.280 ;
        RECT 45.235 128.250 45.615 128.560 ;
        RECT 63.320 127.970 63.700 128.280 ;
        RECT 65.120 128.250 65.500 128.560 ;
        RECT 32.700 127.590 63.740 127.970 ;
        RECT 143.680 127.910 144.680 128.290 ;
        RECT 147.640 127.910 148.640 128.290 ;
        RECT 20.035 127.000 20.415 127.310 ;
        RECT 32.700 127.280 33.080 127.590 ;
        RECT 61.520 127.000 61.900 127.310 ;
        RECT 63.320 127.280 63.700 127.590 ;
        RECT 20.035 126.620 61.940 127.000 ;
        RECT 20.035 126.310 20.415 126.620 ;
        RECT 61.520 126.310 61.900 126.620 ;
        RECT 68.720 126.030 69.100 126.340 ;
        RECT 94.835 126.030 95.215 126.340 ;
        RECT 143.680 126.150 144.680 126.530 ;
        RECT 147.640 126.150 148.640 126.530 ;
        RECT 68.720 125.650 95.215 126.030 ;
        RECT 67.820 125.060 68.200 125.370 ;
        RECT 68.720 125.340 69.100 125.650 ;
        RECT 83.900 125.060 84.280 125.370 ;
        RECT 94.835 125.340 95.215 125.650 ;
        RECT 147.640 125.270 148.640 125.650 ;
        RECT 67.820 124.680 84.280 125.060 ;
        RECT 66.920 124.090 67.300 124.400 ;
        RECT 67.820 124.370 68.200 124.680 ;
        RECT 69.635 124.090 70.015 124.400 ;
        RECT 83.900 124.370 84.280 124.680 ;
        RECT 66.920 123.710 70.015 124.090 ;
        RECT 58.700 123.120 59.080 123.430 ;
        RECT 66.020 123.120 66.400 123.430 ;
        RECT 66.920 123.400 67.300 123.710 ;
        RECT 69.635 123.400 70.015 123.710 ;
        RECT 58.700 122.740 66.440 123.120 ;
        RECT 44.435 122.150 44.815 122.460 ;
        RECT 58.700 122.430 59.080 122.740 ;
        RECT 64.220 122.150 64.600 122.460 ;
        RECT 66.020 122.430 66.400 122.740 ;
        RECT 143.680 122.630 144.680 123.010 ;
        RECT 147.640 122.630 148.640 123.010 ;
        RECT 44.435 121.770 64.640 122.150 ;
        RECT 33.500 121.180 33.880 121.490 ;
        RECT 44.435 121.460 44.815 121.770 ;
        RECT 62.420 121.180 62.800 121.490 ;
        RECT 64.220 121.460 64.600 121.770 ;
        RECT 33.500 120.800 62.840 121.180 ;
        RECT 143.680 120.870 144.680 121.250 ;
        RECT 147.640 120.870 148.640 121.250 ;
        RECT 19.235 120.210 19.615 120.520 ;
        RECT 33.500 120.490 33.880 120.800 ;
        RECT 60.620 120.210 61.000 120.520 ;
        RECT 62.420 120.490 62.800 120.800 ;
        RECT 19.235 119.830 61.040 120.210 ;
        RECT 19.235 119.520 19.615 119.830 ;
        RECT 40.860 119.240 41.240 119.550 ;
        RECT 60.620 119.520 61.000 119.830 ;
        RECT 141.520 119.550 143.300 119.930 ;
        RECT 76.520 119.240 76.900 119.550 ;
        RECT 40.860 118.860 76.940 119.240 ;
        RECT 36.460 118.270 36.840 118.580 ;
        RECT 40.860 118.550 41.240 118.860 ;
        RECT 76.520 118.550 76.900 118.860 ;
        RECT 78.320 118.270 78.700 118.580 ;
        RECT 36.460 117.890 78.740 118.270 ;
        RECT 15.660 117.300 16.040 117.610 ;
        RECT 36.460 117.580 36.840 117.890 ;
        RECT 78.320 117.580 78.700 117.890 ;
        RECT 80.120 117.300 80.500 117.610 ;
        RECT 15.660 116.920 80.540 117.300 ;
        RECT 15.660 116.610 16.040 116.920 ;
        RECT 80.120 116.610 80.500 116.920 ;
        RECT 116.380 115.360 116.760 117.880 ;
        RECT 57.740 114.980 58.740 115.360 ;
        RECT 116.380 114.980 117.380 115.360 ;
        RECT 57.740 110.510 58.120 114.980 ;
        RECT 117.780 113.420 118.160 117.880 ;
        RECT 142.920 114.650 143.300 119.550 ;
        RECT 147.640 117.350 148.640 117.730 ;
        RECT 147.640 116.470 148.640 116.850 ;
        RECT 143.680 115.590 144.680 115.970 ;
        RECT 142.920 114.270 150.800 114.650 ;
        RECT 83.000 113.040 84.000 113.420 ;
        RECT 117.780 113.040 118.780 113.420 ;
        RECT 83.000 110.510 83.380 113.040 ;
        RECT 143.680 112.070 144.680 112.450 ;
        RECT 147.640 112.070 148.640 112.450 ;
        RECT 12.240 40.610 12.620 110.510 ;
        RECT 23.440 108.810 23.820 109.810 ;
        RECT 60.620 109.500 61.000 109.810 ;
        RECT 58.760 109.120 61.000 109.500 ;
        RECT 60.620 108.810 61.000 109.120 ;
        RECT 80.120 109.500 80.500 109.810 ;
        RECT 80.120 109.120 82.360 109.500 ;
        RECT 80.120 108.810 80.500 109.120 ;
        RECT 117.300 108.810 117.680 109.810 ;
        RECT 22.040 105.750 22.420 106.750 ;
        RECT 26.240 105.750 26.620 106.750 ;
        RECT 44.440 105.750 44.820 106.750 ;
        RECT 48.640 105.750 49.020 106.750 ;
        RECT 60.620 106.440 61.000 106.750 ;
        RECT 58.760 106.060 61.000 106.440 ;
        RECT 60.620 105.750 61.000 106.060 ;
        RECT 80.120 106.440 80.500 106.750 ;
        RECT 80.120 106.060 82.360 106.440 ;
        RECT 80.120 105.750 80.500 106.060 ;
        RECT 92.100 105.750 92.480 106.750 ;
        RECT 96.300 105.750 96.680 106.750 ;
        RECT 114.500 105.750 114.880 106.750 ;
        RECT 118.700 105.750 119.080 106.750 ;
        RECT 19.240 102.690 19.620 103.690 ;
        RECT 20.640 102.690 21.020 103.690 ;
        RECT 27.640 102.690 28.020 103.690 ;
        RECT 29.040 102.690 29.420 103.690 ;
        RECT 41.640 102.690 42.020 103.690 ;
        RECT 43.040 102.690 43.420 103.690 ;
        RECT 50.040 102.690 50.420 103.690 ;
        RECT 51.440 102.690 51.820 103.690 ;
        RECT 60.620 103.380 61.000 103.690 ;
        RECT 58.760 103.000 61.000 103.380 ;
        RECT 60.620 102.690 61.000 103.000 ;
        RECT 80.120 103.380 80.500 103.690 ;
        RECT 80.120 103.000 82.360 103.380 ;
        RECT 80.120 102.690 80.500 103.000 ;
        RECT 89.300 102.690 89.680 103.690 ;
        RECT 90.700 102.690 91.080 103.690 ;
        RECT 97.700 102.690 98.080 103.690 ;
        RECT 99.100 102.690 99.480 103.690 ;
        RECT 111.700 102.690 112.080 103.690 ;
        RECT 113.100 102.690 113.480 103.690 ;
        RECT 120.100 102.690 120.480 103.690 ;
        RECT 121.500 102.690 121.880 103.690 ;
        RECT 24.840 99.630 25.220 100.630 ;
        RECT 45.840 99.630 46.220 100.630 ;
        RECT 60.620 100.320 61.000 100.630 ;
        RECT 58.760 99.940 61.000 100.320 ;
        RECT 60.620 99.630 61.000 99.940 ;
        RECT 80.120 100.320 80.500 100.630 ;
        RECT 80.120 99.940 82.360 100.320 ;
        RECT 80.120 99.630 80.500 99.940 ;
        RECT 94.900 99.630 95.280 100.630 ;
        RECT 115.900 99.630 116.280 100.630 ;
        RECT 13.640 96.570 14.020 97.570 ;
        RECT 15.040 96.570 15.420 97.570 ;
        RECT 16.440 96.570 16.820 97.570 ;
        RECT 17.840 96.570 18.220 97.570 ;
        RECT 30.440 96.570 30.820 97.570 ;
        RECT 31.840 96.570 32.220 97.570 ;
        RECT 33.240 96.570 33.620 97.570 ;
        RECT 34.640 96.570 35.020 97.570 ;
        RECT 36.040 96.570 36.420 97.570 ;
        RECT 37.440 96.570 37.820 97.570 ;
        RECT 38.840 96.570 39.220 97.570 ;
        RECT 40.240 96.570 40.620 97.570 ;
        RECT 52.840 96.570 53.220 97.570 ;
        RECT 54.240 96.570 54.620 97.570 ;
        RECT 55.640 96.570 56.020 97.570 ;
        RECT 57.040 96.570 57.420 97.570 ;
        RECT 60.620 97.260 61.000 97.570 ;
        RECT 58.760 96.880 61.000 97.260 ;
        RECT 60.620 96.570 61.000 96.880 ;
        RECT 80.120 97.260 80.500 97.570 ;
        RECT 80.120 96.880 82.360 97.260 ;
        RECT 80.120 96.570 80.500 96.880 ;
        RECT 83.700 96.570 84.080 97.570 ;
        RECT 85.100 96.570 85.480 97.570 ;
        RECT 86.500 96.570 86.880 97.570 ;
        RECT 87.900 96.570 88.280 97.570 ;
        RECT 100.500 96.570 100.880 97.570 ;
        RECT 101.900 96.570 102.280 97.570 ;
        RECT 103.300 96.570 103.680 97.570 ;
        RECT 104.700 96.570 105.080 97.570 ;
        RECT 106.100 96.570 106.480 97.570 ;
        RECT 107.500 96.570 107.880 97.570 ;
        RECT 108.900 96.570 109.280 97.570 ;
        RECT 110.300 96.570 110.680 97.570 ;
        RECT 122.900 96.570 123.280 97.570 ;
        RECT 124.300 96.570 124.680 97.570 ;
        RECT 125.700 96.570 126.080 97.570 ;
        RECT 127.100 96.570 127.480 97.570 ;
        RECT 47.240 93.510 47.620 94.510 ;
        RECT 60.620 94.200 61.000 94.510 ;
        RECT 58.760 93.820 61.000 94.200 ;
        RECT 60.620 93.510 61.000 93.820 ;
        RECT 80.120 94.200 80.500 94.510 ;
        RECT 80.120 93.820 82.360 94.200 ;
        RECT 80.120 93.510 80.500 93.820 ;
        RECT 93.500 93.510 93.880 94.510 ;
        RECT 23.440 91.410 23.820 92.410 ;
        RECT 64.220 92.100 64.600 92.410 ;
        RECT 58.760 91.720 64.600 92.100 ;
        RECT 64.220 91.410 64.600 91.720 ;
        RECT 76.520 92.100 76.900 92.410 ;
        RECT 76.520 91.720 82.360 92.100 ;
        RECT 76.520 91.410 76.900 91.720 ;
        RECT 117.300 91.410 117.680 92.410 ;
        RECT 22.040 88.350 22.420 89.350 ;
        RECT 26.240 88.350 26.620 89.350 ;
        RECT 44.440 88.350 44.820 89.350 ;
        RECT 48.640 88.350 49.020 89.350 ;
        RECT 64.220 89.040 64.600 89.350 ;
        RECT 58.760 88.660 64.600 89.040 ;
        RECT 64.220 88.350 64.600 88.660 ;
        RECT 76.520 89.040 76.900 89.350 ;
        RECT 76.520 88.660 82.360 89.040 ;
        RECT 76.520 88.350 76.900 88.660 ;
        RECT 92.100 88.350 92.480 89.350 ;
        RECT 96.300 88.350 96.680 89.350 ;
        RECT 114.500 88.350 114.880 89.350 ;
        RECT 118.700 88.350 119.080 89.350 ;
        RECT 19.240 85.290 19.620 86.290 ;
        RECT 20.640 85.290 21.020 86.290 ;
        RECT 27.640 85.290 28.020 86.290 ;
        RECT 29.040 85.290 29.420 86.290 ;
        RECT 41.640 85.290 42.020 86.290 ;
        RECT 43.040 85.290 43.420 86.290 ;
        RECT 50.040 85.290 50.420 86.290 ;
        RECT 51.440 85.290 51.820 86.290 ;
        RECT 65.120 85.980 65.500 86.290 ;
        RECT 58.760 85.600 65.500 85.980 ;
        RECT 65.120 85.290 65.500 85.600 ;
        RECT 75.620 85.980 76.000 86.290 ;
        RECT 75.620 85.600 82.360 85.980 ;
        RECT 75.620 85.290 76.000 85.600 ;
        RECT 89.300 85.290 89.680 86.290 ;
        RECT 90.700 85.290 91.080 86.290 ;
        RECT 97.700 85.290 98.080 86.290 ;
        RECT 99.100 85.290 99.480 86.290 ;
        RECT 111.700 85.290 112.080 86.290 ;
        RECT 113.100 85.290 113.480 86.290 ;
        RECT 120.100 85.290 120.480 86.290 ;
        RECT 121.500 85.290 121.880 86.290 ;
        RECT 24.840 82.230 25.220 83.230 ;
        RECT 45.840 82.230 46.220 83.230 ;
        RECT 64.220 82.920 64.600 83.230 ;
        RECT 58.760 82.540 64.600 82.920 ;
        RECT 64.220 82.230 64.600 82.540 ;
        RECT 76.520 82.920 76.900 83.230 ;
        RECT 76.520 82.540 82.360 82.920 ;
        RECT 76.520 82.230 76.900 82.540 ;
        RECT 94.900 82.230 95.280 83.230 ;
        RECT 115.900 82.230 116.280 83.230 ;
        RECT 13.640 79.170 14.020 80.170 ;
        RECT 15.040 79.170 15.420 80.170 ;
        RECT 16.440 79.170 16.820 80.170 ;
        RECT 17.840 79.170 18.220 80.170 ;
        RECT 30.440 79.170 30.820 80.170 ;
        RECT 31.840 79.170 32.220 80.170 ;
        RECT 33.240 79.170 33.620 80.170 ;
        RECT 34.640 79.170 35.020 80.170 ;
        RECT 36.040 79.170 36.420 80.170 ;
        RECT 37.440 79.170 37.820 80.170 ;
        RECT 38.840 79.170 39.220 80.170 ;
        RECT 40.240 79.170 40.620 80.170 ;
        RECT 52.840 79.170 53.220 80.170 ;
        RECT 54.240 79.170 54.620 80.170 ;
        RECT 55.640 79.170 56.020 80.170 ;
        RECT 57.040 79.170 57.420 80.170 ;
        RECT 63.320 79.860 63.700 80.170 ;
        RECT 58.760 79.480 63.700 79.860 ;
        RECT 63.320 79.170 63.700 79.480 ;
        RECT 77.420 79.860 77.800 80.170 ;
        RECT 77.420 79.480 82.360 79.860 ;
        RECT 77.420 79.170 77.800 79.480 ;
        RECT 83.700 79.170 84.080 80.170 ;
        RECT 85.100 79.170 85.480 80.170 ;
        RECT 86.500 79.170 86.880 80.170 ;
        RECT 87.900 79.170 88.280 80.170 ;
        RECT 100.500 79.170 100.880 80.170 ;
        RECT 101.900 79.170 102.280 80.170 ;
        RECT 103.300 79.170 103.680 80.170 ;
        RECT 104.700 79.170 105.080 80.170 ;
        RECT 106.100 79.170 106.480 80.170 ;
        RECT 107.500 79.170 107.880 80.170 ;
        RECT 108.900 79.170 109.280 80.170 ;
        RECT 110.300 79.170 110.680 80.170 ;
        RECT 122.900 79.170 123.280 80.170 ;
        RECT 124.300 79.170 124.680 80.170 ;
        RECT 125.700 79.170 126.080 80.170 ;
        RECT 127.100 79.170 127.480 80.170 ;
        RECT 47.240 76.110 47.620 77.110 ;
        RECT 64.220 76.800 64.600 77.110 ;
        RECT 58.760 76.420 64.600 76.800 ;
        RECT 64.220 76.110 64.600 76.420 ;
        RECT 76.520 76.800 76.900 77.110 ;
        RECT 76.520 76.420 82.360 76.800 ;
        RECT 76.520 76.110 76.900 76.420 ;
        RECT 93.500 76.110 93.880 77.110 ;
        RECT 23.440 74.010 23.820 75.010 ;
        RECT 68.720 74.700 69.100 75.010 ;
        RECT 58.760 74.320 69.100 74.700 ;
        RECT 68.720 74.010 69.100 74.320 ;
        RECT 72.020 74.700 72.400 75.010 ;
        RECT 72.020 74.320 82.360 74.700 ;
        RECT 72.020 74.010 72.400 74.320 ;
        RECT 117.300 74.010 117.680 75.010 ;
        RECT 22.040 70.950 22.420 71.950 ;
        RECT 26.240 70.950 26.620 71.950 ;
        RECT 44.440 70.950 44.820 71.950 ;
        RECT 48.640 70.950 49.020 71.950 ;
        RECT 66.920 71.640 67.300 71.950 ;
        RECT 58.760 71.260 67.300 71.640 ;
        RECT 66.920 70.950 67.300 71.260 ;
        RECT 73.820 71.640 74.200 71.950 ;
        RECT 73.820 71.260 82.360 71.640 ;
        RECT 73.820 70.950 74.200 71.260 ;
        RECT 92.100 70.950 92.480 71.950 ;
        RECT 96.300 70.950 96.680 71.950 ;
        RECT 114.500 70.950 114.880 71.950 ;
        RECT 118.700 70.950 119.080 71.950 ;
        RECT 19.240 67.890 19.620 68.890 ;
        RECT 20.640 67.890 21.020 68.890 ;
        RECT 27.640 67.890 28.020 68.890 ;
        RECT 29.040 67.890 29.420 68.890 ;
        RECT 41.640 67.890 42.020 68.890 ;
        RECT 43.040 67.890 43.420 68.890 ;
        RECT 50.040 67.890 50.420 68.890 ;
        RECT 51.440 67.890 51.820 68.890 ;
        RECT 66.020 68.580 66.400 68.890 ;
        RECT 58.760 68.200 66.400 68.580 ;
        RECT 66.020 67.890 66.400 68.200 ;
        RECT 74.720 68.580 75.100 68.890 ;
        RECT 74.720 68.200 82.360 68.580 ;
        RECT 74.720 67.890 75.100 68.200 ;
        RECT 89.300 67.890 89.680 68.890 ;
        RECT 90.700 67.890 91.080 68.890 ;
        RECT 97.700 67.890 98.080 68.890 ;
        RECT 99.100 67.890 99.480 68.890 ;
        RECT 111.700 67.890 112.080 68.890 ;
        RECT 113.100 67.890 113.480 68.890 ;
        RECT 120.100 67.890 120.480 68.890 ;
        RECT 121.500 67.890 121.880 68.890 ;
        RECT 24.840 64.830 25.220 65.830 ;
        RECT 45.840 64.830 46.220 65.830 ;
        RECT 67.820 65.520 68.200 65.830 ;
        RECT 58.760 65.140 68.200 65.520 ;
        RECT 67.820 64.830 68.200 65.140 ;
        RECT 72.920 65.520 73.300 65.830 ;
        RECT 72.920 65.140 82.360 65.520 ;
        RECT 72.920 64.830 73.300 65.140 ;
        RECT 94.900 64.830 95.280 65.830 ;
        RECT 115.900 64.830 116.280 65.830 ;
        RECT 13.640 61.770 14.020 62.770 ;
        RECT 15.040 61.770 15.420 62.770 ;
        RECT 16.440 61.770 16.820 62.770 ;
        RECT 17.840 61.770 18.220 62.770 ;
        RECT 30.440 61.770 30.820 62.770 ;
        RECT 31.840 61.770 32.220 62.770 ;
        RECT 33.240 61.770 33.620 62.770 ;
        RECT 34.640 61.770 35.020 62.770 ;
        RECT 36.040 61.770 36.420 62.770 ;
        RECT 37.440 61.770 37.820 62.770 ;
        RECT 38.840 61.770 39.220 62.770 ;
        RECT 40.240 61.770 40.620 62.770 ;
        RECT 52.840 61.770 53.220 62.770 ;
        RECT 54.240 61.770 54.620 62.770 ;
        RECT 55.640 61.770 56.020 62.770 ;
        RECT 57.040 61.770 57.420 62.770 ;
        RECT 62.420 62.460 62.800 62.770 ;
        RECT 58.760 62.080 62.800 62.460 ;
        RECT 62.420 61.770 62.800 62.080 ;
        RECT 78.320 62.460 78.700 62.770 ;
        RECT 78.320 62.080 82.360 62.460 ;
        RECT 78.320 61.770 78.700 62.080 ;
        RECT 83.700 61.770 84.080 62.770 ;
        RECT 85.100 61.770 85.480 62.770 ;
        RECT 86.500 61.770 86.880 62.770 ;
        RECT 87.900 61.770 88.280 62.770 ;
        RECT 100.500 61.770 100.880 62.770 ;
        RECT 101.900 61.770 102.280 62.770 ;
        RECT 103.300 61.770 103.680 62.770 ;
        RECT 104.700 61.770 105.080 62.770 ;
        RECT 106.100 61.770 106.480 62.770 ;
        RECT 107.500 61.770 107.880 62.770 ;
        RECT 108.900 61.770 109.280 62.770 ;
        RECT 110.300 61.770 110.680 62.770 ;
        RECT 122.900 61.770 123.280 62.770 ;
        RECT 124.300 61.770 124.680 62.770 ;
        RECT 125.700 61.770 126.080 62.770 ;
        RECT 127.100 61.770 127.480 62.770 ;
        RECT 47.240 58.710 47.620 59.710 ;
        RECT 93.500 58.710 93.880 59.710 ;
        RECT 23.440 56.610 23.820 57.610 ;
        RECT 61.520 57.300 61.900 57.610 ;
        RECT 58.760 56.920 61.900 57.300 ;
        RECT 61.520 56.610 61.900 56.920 ;
        RECT 79.220 57.300 79.600 57.610 ;
        RECT 79.220 56.920 82.360 57.300 ;
        RECT 79.220 56.610 79.600 56.920 ;
        RECT 117.300 56.610 117.680 57.610 ;
        RECT 22.040 53.550 22.420 54.550 ;
        RECT 26.240 53.550 26.620 54.550 ;
        RECT 44.440 53.550 44.820 54.550 ;
        RECT 48.640 53.550 49.020 54.550 ;
        RECT 61.520 54.240 61.900 54.550 ;
        RECT 58.760 53.860 61.900 54.240 ;
        RECT 61.520 53.550 61.900 53.860 ;
        RECT 79.220 54.240 79.600 54.550 ;
        RECT 79.220 53.860 82.360 54.240 ;
        RECT 79.220 53.550 79.600 53.860 ;
        RECT 92.100 53.550 92.480 54.550 ;
        RECT 96.300 53.550 96.680 54.550 ;
        RECT 114.500 53.550 114.880 54.550 ;
        RECT 118.700 53.550 119.080 54.550 ;
        RECT 19.240 50.490 19.620 51.490 ;
        RECT 20.640 50.490 21.020 51.490 ;
        RECT 27.640 50.490 28.020 51.490 ;
        RECT 29.040 50.490 29.420 51.490 ;
        RECT 41.640 50.490 42.020 51.490 ;
        RECT 43.040 50.490 43.420 51.490 ;
        RECT 50.040 50.490 50.420 51.490 ;
        RECT 51.440 50.490 51.820 51.490 ;
        RECT 61.520 51.180 61.900 51.490 ;
        RECT 58.760 50.800 61.900 51.180 ;
        RECT 61.520 50.490 61.900 50.800 ;
        RECT 79.220 51.180 79.600 51.490 ;
        RECT 79.220 50.800 82.360 51.180 ;
        RECT 79.220 50.490 79.600 50.800 ;
        RECT 89.300 50.490 89.680 51.490 ;
        RECT 90.700 50.490 91.080 51.490 ;
        RECT 97.700 50.490 98.080 51.490 ;
        RECT 99.100 50.490 99.480 51.490 ;
        RECT 111.700 50.490 112.080 51.490 ;
        RECT 113.100 50.490 113.480 51.490 ;
        RECT 120.100 50.490 120.480 51.490 ;
        RECT 121.500 50.490 121.880 51.490 ;
        RECT 24.840 47.430 25.220 48.430 ;
        RECT 45.840 47.430 46.220 48.430 ;
        RECT 61.520 48.120 61.900 48.430 ;
        RECT 58.760 47.740 61.900 48.120 ;
        RECT 61.520 47.430 61.900 47.740 ;
        RECT 79.220 48.120 79.600 48.430 ;
        RECT 79.220 47.740 82.360 48.120 ;
        RECT 79.220 47.430 79.600 47.740 ;
        RECT 94.900 47.430 95.280 48.430 ;
        RECT 115.900 47.430 116.280 48.430 ;
        RECT 13.640 44.370 14.020 45.370 ;
        RECT 15.040 44.370 15.420 45.370 ;
        RECT 16.440 44.370 16.820 45.370 ;
        RECT 17.840 44.370 18.220 45.370 ;
        RECT 30.440 44.370 30.820 45.370 ;
        RECT 31.840 44.370 32.220 45.370 ;
        RECT 33.240 44.370 33.620 45.370 ;
        RECT 34.640 44.370 35.020 45.370 ;
        RECT 36.040 44.370 36.420 45.370 ;
        RECT 37.440 44.370 37.820 45.370 ;
        RECT 38.840 44.370 39.220 45.370 ;
        RECT 40.240 44.370 40.620 45.370 ;
        RECT 52.840 44.370 53.220 45.370 ;
        RECT 54.240 44.370 54.620 45.370 ;
        RECT 55.640 44.370 56.020 45.370 ;
        RECT 57.040 44.370 57.420 45.370 ;
        RECT 61.520 45.060 61.900 45.370 ;
        RECT 58.760 44.680 61.900 45.060 ;
        RECT 61.520 44.370 61.900 44.680 ;
        RECT 79.220 45.060 79.600 45.370 ;
        RECT 79.220 44.680 82.360 45.060 ;
        RECT 79.220 44.370 79.600 44.680 ;
        RECT 83.700 44.370 84.080 45.370 ;
        RECT 85.100 44.370 85.480 45.370 ;
        RECT 86.500 44.370 86.880 45.370 ;
        RECT 87.900 44.370 88.280 45.370 ;
        RECT 100.500 44.370 100.880 45.370 ;
        RECT 101.900 44.370 102.280 45.370 ;
        RECT 103.300 44.370 103.680 45.370 ;
        RECT 104.700 44.370 105.080 45.370 ;
        RECT 106.100 44.370 106.480 45.370 ;
        RECT 107.500 44.370 107.880 45.370 ;
        RECT 108.900 44.370 109.280 45.370 ;
        RECT 110.300 44.370 110.680 45.370 ;
        RECT 122.900 44.370 123.280 45.370 ;
        RECT 124.300 44.370 124.680 45.370 ;
        RECT 125.700 44.370 126.080 45.370 ;
        RECT 127.100 44.370 127.480 45.370 ;
        RECT 47.240 41.310 47.620 42.310 ;
        RECT 61.520 42.000 61.900 42.310 ;
        RECT 58.760 41.620 61.900 42.000 ;
        RECT 61.520 41.310 61.900 41.620 ;
        RECT 79.220 42.000 79.600 42.310 ;
        RECT 79.220 41.620 82.360 42.000 ;
        RECT 79.220 41.310 79.600 41.620 ;
        RECT 93.500 41.310 93.880 42.310 ;
        RECT 128.500 40.610 128.880 110.510 ;
        RECT 143.680 110.310 144.680 110.690 ;
        RECT 147.640 110.310 148.640 110.690 ;
        RECT 143.680 106.790 144.680 107.170 ;
        RECT 147.640 106.790 148.640 107.170 ;
        RECT 143.680 103.270 144.680 103.650 ;
        RECT 147.640 103.270 148.640 103.650 ;
        RECT 143.680 101.510 144.680 101.890 ;
        RECT 147.640 101.510 148.640 101.890 ;
        RECT 147.640 100.630 148.640 101.010 ;
        RECT 143.680 97.990 144.680 98.370 ;
        RECT 147.640 97.990 148.640 98.370 ;
        RECT 143.680 96.230 144.680 96.610 ;
        RECT 147.640 96.230 148.640 96.610 ;
        RECT 141.520 94.910 143.300 95.290 ;
        RECT 142.920 90.010 143.300 94.910 ;
        RECT 147.640 92.710 148.640 93.090 ;
        RECT 147.640 91.830 148.640 92.210 ;
        RECT 143.680 90.950 144.680 91.330 ;
        RECT 142.920 89.630 150.800 90.010 ;
        RECT 143.680 87.430 144.680 87.810 ;
        RECT 147.640 87.430 148.640 87.810 ;
        RECT 143.680 85.670 144.680 86.050 ;
        RECT 147.640 85.670 148.640 86.050 ;
        RECT 143.680 82.150 144.680 82.530 ;
        RECT 147.640 82.150 148.640 82.530 ;
        RECT 143.680 78.630 144.680 79.010 ;
        RECT 147.640 78.630 148.640 79.010 ;
        RECT 143.680 76.870 144.680 77.250 ;
        RECT 147.640 76.870 148.640 77.250 ;
        RECT 147.640 75.990 148.640 76.370 ;
        RECT 143.680 73.350 144.680 73.730 ;
        RECT 147.640 73.350 148.640 73.730 ;
        RECT 143.680 71.590 144.680 71.970 ;
        RECT 147.640 71.590 148.640 71.970 ;
        RECT 141.520 70.270 143.300 70.650 ;
        RECT 142.920 65.370 143.300 70.270 ;
        RECT 147.640 68.070 148.640 68.450 ;
        RECT 147.640 67.190 148.640 67.570 ;
        RECT 143.680 66.310 144.680 66.690 ;
        RECT 142.920 64.990 150.800 65.370 ;
        RECT 143.680 62.790 144.680 63.170 ;
        RECT 147.640 62.790 148.640 63.170 ;
        RECT 143.680 61.030 144.680 61.410 ;
        RECT 147.640 61.030 148.640 61.410 ;
        RECT 143.680 57.510 144.680 57.890 ;
        RECT 147.640 57.510 148.640 57.890 ;
        RECT 143.680 53.990 144.680 54.370 ;
        RECT 147.640 53.990 148.640 54.370 ;
        RECT 143.680 52.230 144.680 52.610 ;
        RECT 147.640 52.230 148.640 52.610 ;
        RECT 147.640 51.350 148.640 51.730 ;
        RECT 143.680 48.710 144.680 49.090 ;
        RECT 147.640 48.710 148.640 49.090 ;
        RECT 143.680 46.950 144.680 47.330 ;
        RECT 147.640 46.950 148.640 47.330 ;
        RECT 141.520 45.630 143.300 46.010 ;
        RECT 142.920 40.730 143.300 45.630 ;
        RECT 147.640 43.430 148.640 43.810 ;
        RECT 147.640 42.550 148.640 42.930 ;
        RECT 143.680 41.670 144.680 42.050 ;
        RECT 142.920 40.350 150.800 40.730 ;
        RECT 13.600 38.540 49.240 38.980 ;
        RECT 13.600 37.660 48.520 38.100 ;
        RECT 13.600 36.340 13.960 37.660 ;
        RECT 48.880 37.220 49.240 38.540 ;
        RECT 14.320 36.780 49.240 37.220 ;
        RECT 13.600 35.900 48.520 36.340 ;
        RECT 13.600 34.580 13.960 35.900 ;
        RECT 48.880 35.460 49.240 36.780 ;
        RECT 14.320 35.020 49.240 35.460 ;
        RECT 92.080 38.540 127.720 38.980 ;
        RECT 92.080 37.220 92.440 38.540 ;
        RECT 143.680 38.150 144.680 38.530 ;
        RECT 147.640 38.150 148.640 38.530 ;
        RECT 92.800 37.660 127.720 38.100 ;
        RECT 92.080 36.780 127.000 37.220 ;
        RECT 92.080 35.460 92.440 36.780 ;
        RECT 127.360 36.340 127.720 37.660 ;
        RECT 143.680 36.390 144.680 36.770 ;
        RECT 147.640 36.390 148.640 36.770 ;
        RECT 92.800 35.900 127.720 36.340 ;
        RECT 92.080 35.020 127.000 35.460 ;
        RECT 127.360 34.580 127.720 35.900 ;
        RECT 13.600 34.140 49.240 34.580 ;
        RECT 92.080 34.140 127.720 34.580 ;
        RECT 13.600 33.260 49.240 33.700 ;
        RECT 13.600 32.380 48.520 32.820 ;
        RECT 13.600 31.060 13.960 32.380 ;
        RECT 48.880 31.940 49.240 33.260 ;
        RECT 92.080 33.260 127.720 33.700 ;
        RECT 54.720 32.010 55.720 32.390 ;
        RECT 58.680 32.010 59.680 32.390 ;
        RECT 81.640 32.010 82.640 32.390 ;
        RECT 85.600 32.010 86.600 32.390 ;
        RECT 14.320 31.500 49.240 31.940 ;
        RECT 92.080 31.940 92.440 33.260 ;
        RECT 143.680 32.870 144.680 33.250 ;
        RECT 147.640 32.870 148.640 33.250 ;
        RECT 92.800 32.380 127.720 32.820 ;
        RECT 13.600 30.620 48.520 31.060 ;
        RECT 13.600 29.300 13.960 30.620 ;
        RECT 48.880 30.180 49.240 31.500 ;
        RECT 54.720 31.130 55.720 31.510 ;
        RECT 58.680 31.130 59.680 31.510 ;
        RECT 81.640 31.130 82.640 31.510 ;
        RECT 85.600 31.130 86.600 31.510 ;
        RECT 92.080 31.500 127.000 31.940 ;
        RECT 61.600 30.210 62.600 30.590 ;
        RECT 78.720 30.210 79.720 30.590 ;
        RECT 14.320 29.740 49.240 30.180 ;
        RECT 92.080 30.180 92.440 31.500 ;
        RECT 127.360 31.060 127.720 32.380 ;
        RECT 92.800 30.620 127.720 31.060 ;
        RECT 54.720 29.370 55.720 29.750 ;
        RECT 58.680 29.370 59.680 29.750 ;
        RECT 81.640 29.370 82.640 29.750 ;
        RECT 85.600 29.370 86.600 29.750 ;
        RECT 92.080 29.740 127.000 30.180 ;
        RECT 127.360 29.300 127.720 30.620 ;
        RECT 143.680 29.350 144.680 29.730 ;
        RECT 147.640 29.350 148.640 29.730 ;
        RECT 13.600 28.860 49.240 29.300 ;
        RECT 54.720 28.490 55.720 28.870 ;
        RECT 58.680 28.490 59.680 28.870 ;
        RECT 81.640 28.490 82.640 28.870 ;
        RECT 85.600 28.490 86.600 28.870 ;
        RECT 92.080 28.860 127.720 29.300 ;
        RECT 13.600 27.980 49.240 28.420 ;
        RECT 13.600 27.100 48.520 27.540 ;
        RECT 13.600 25.780 13.960 27.100 ;
        RECT 48.880 26.660 49.240 27.980 ;
        RECT 54.720 27.610 55.720 27.990 ;
        RECT 58.680 27.610 59.680 27.990 ;
        RECT 81.640 27.610 82.640 27.990 ;
        RECT 85.600 27.610 86.600 27.990 ;
        RECT 92.080 27.980 127.720 28.420 ;
        RECT 14.320 26.220 49.240 26.660 ;
        RECT 92.080 26.660 92.440 27.980 ;
        RECT 143.680 27.590 144.680 27.970 ;
        RECT 147.640 27.590 148.640 27.970 ;
        RECT 92.800 27.100 127.720 27.540 ;
        RECT 13.600 25.340 48.520 25.780 ;
        RECT 13.600 24.020 13.960 25.340 ;
        RECT 48.880 24.900 49.240 26.220 ;
        RECT 54.720 25.850 55.720 26.230 ;
        RECT 58.680 25.850 59.680 26.230 ;
        RECT 65.800 25.850 67.580 26.230 ;
        RECT 74.440 25.850 75.440 26.230 ;
        RECT 81.640 25.850 82.640 26.230 ;
        RECT 85.600 25.850 86.600 26.230 ;
        RECT 92.080 26.220 127.000 26.660 ;
        RECT 54.720 24.970 55.720 25.350 ;
        RECT 58.600 24.970 63.580 25.350 ;
        RECT 14.320 24.460 49.240 24.900 ;
        RECT 13.600 23.580 49.240 24.020 ;
        RECT 52.560 23.210 53.560 23.590 ;
        RECT 13.600 22.700 49.240 23.140 ;
        RECT 60.060 22.770 61.840 23.150 ;
        RECT 13.600 21.820 48.520 22.260 ;
        RECT 13.600 20.500 13.960 21.820 ;
        RECT 48.880 21.380 49.240 22.700 ;
        RECT 58.680 22.330 59.680 22.710 ;
        RECT 14.320 20.940 49.240 21.380 ;
        RECT 13.600 20.060 48.520 20.500 ;
        RECT 13.600 18.740 13.960 20.060 ;
        RECT 48.880 19.620 49.240 20.940 ;
        RECT 53.940 20.570 55.720 20.950 ;
        RECT 14.320 19.180 49.240 19.620 ;
        RECT 52.560 19.250 53.560 19.630 ;
        RECT 13.600 18.300 49.240 18.740 ;
        RECT 13.600 17.420 49.240 17.860 ;
        RECT 13.600 16.540 48.520 16.980 ;
        RECT 13.600 15.220 13.960 16.540 ;
        RECT 48.880 16.100 49.240 17.420 ;
        RECT 14.320 15.660 49.240 16.100 ;
        RECT 13.600 14.780 48.520 15.220 ;
        RECT 13.600 13.460 13.960 14.780 ;
        RECT 48.880 14.340 49.240 15.660 ;
        RECT 14.320 13.900 49.240 14.340 ;
        RECT 13.600 13.400 49.240 13.460 ;
        RECT 53.940 13.400 54.320 20.570 ;
        RECT 54.720 18.810 55.720 19.190 ;
        RECT 58.680 18.810 59.680 19.190 ;
        RECT 54.720 17.930 55.720 18.310 ;
        RECT 58.680 17.930 59.680 18.310 ;
        RECT 58.680 16.700 59.680 16.740 ;
        RECT 60.060 16.700 60.440 22.770 ;
        RECT 63.200 17.870 63.580 24.970 ;
        RECT 67.200 19.190 67.580 25.850 ;
        RECT 77.740 24.970 82.720 25.350 ;
        RECT 85.600 24.970 86.600 25.350 ;
        RECT 65.800 18.810 66.800 19.190 ;
        RECT 67.200 18.810 75.440 19.190 ;
        RECT 77.740 17.870 78.120 24.970 ;
        RECT 92.080 24.900 92.440 26.220 ;
        RECT 127.360 25.780 127.720 27.100 ;
        RECT 147.640 26.710 148.640 27.090 ;
        RECT 92.800 25.340 127.720 25.780 ;
        RECT 92.080 24.460 127.000 24.900 ;
        RECT 127.360 24.020 127.720 25.340 ;
        RECT 143.680 24.070 144.680 24.450 ;
        RECT 147.640 24.070 148.640 24.450 ;
        RECT 87.760 23.210 88.760 23.590 ;
        RECT 92.080 23.580 127.720 24.020 ;
        RECT 79.480 22.770 81.260 23.150 ;
        RECT 63.200 17.490 68.960 17.870 ;
        RECT 72.360 17.490 78.120 17.870 ;
        RECT 58.680 16.360 60.440 16.700 ;
        RECT 59.140 16.320 60.440 16.360 ;
        RECT 80.880 16.700 81.260 22.770 ;
        RECT 81.640 22.330 82.640 22.710 ;
        RECT 92.080 22.700 127.720 23.140 ;
        RECT 92.080 21.380 92.440 22.700 ;
        RECT 143.680 22.310 144.680 22.690 ;
        RECT 147.640 22.310 148.640 22.690 ;
        RECT 92.800 21.820 127.720 22.260 ;
        RECT 85.600 20.570 87.380 20.950 ;
        RECT 81.640 18.810 82.640 19.190 ;
        RECT 85.600 18.810 86.600 19.190 ;
        RECT 81.640 17.930 82.640 18.310 ;
        RECT 85.600 17.930 86.600 18.310 ;
        RECT 81.640 16.700 82.640 16.740 ;
        RECT 80.880 16.360 82.640 16.700 ;
        RECT 80.880 16.320 82.180 16.360 ;
        RECT 54.720 15.290 55.720 15.670 ;
        RECT 58.680 15.290 59.680 15.670 ;
        RECT 81.640 15.290 82.640 15.670 ;
        RECT 85.600 15.290 86.600 15.670 ;
        RECT 54.720 14.410 55.720 14.790 ;
        RECT 58.680 14.410 59.680 14.790 ;
        RECT 65.800 14.370 66.800 14.750 ;
        RECT 74.520 14.370 75.520 14.750 ;
        RECT 81.640 14.410 82.640 14.790 ;
        RECT 85.600 14.410 86.600 14.790 ;
        RECT 54.720 13.530 55.720 13.910 ;
        RECT 58.680 13.530 59.680 13.910 ;
        RECT 81.640 13.530 82.640 13.910 ;
        RECT 85.600 13.530 86.600 13.910 ;
        RECT 13.600 13.020 54.320 13.400 ;
        RECT 87.000 13.400 87.380 20.570 ;
        RECT 92.080 20.940 127.000 21.380 ;
        RECT 87.760 19.250 88.760 19.630 ;
        RECT 92.080 19.620 92.440 20.940 ;
        RECT 127.360 20.500 127.720 21.820 ;
        RECT 147.640 21.430 148.640 21.810 ;
        RECT 92.800 20.060 127.720 20.500 ;
        RECT 92.080 19.180 127.000 19.620 ;
        RECT 127.360 18.740 127.720 20.060 ;
        RECT 143.680 18.790 144.680 19.170 ;
        RECT 147.640 18.790 148.640 19.170 ;
        RECT 92.080 18.300 127.720 18.740 ;
        RECT 92.080 17.420 127.720 17.860 ;
        RECT 92.080 16.100 92.440 17.420 ;
        RECT 143.680 17.030 144.680 17.410 ;
        RECT 147.640 17.030 148.640 17.410 ;
        RECT 92.800 16.540 127.720 16.980 ;
        RECT 92.080 15.660 127.000 16.100 ;
        RECT 92.080 14.340 92.440 15.660 ;
        RECT 127.360 15.220 127.720 16.540 ;
        RECT 143.680 15.270 144.680 15.650 ;
        RECT 147.640 15.270 148.640 15.650 ;
        RECT 92.800 14.780 127.720 15.220 ;
        RECT 92.080 13.900 127.000 14.340 ;
        RECT 127.360 13.460 127.720 14.780 ;
        RECT 143.680 14.390 144.680 14.770 ;
        RECT 92.080 13.400 127.720 13.460 ;
        RECT 87.000 13.020 127.720 13.400 ;
        RECT 143.680 11.750 144.680 12.130 ;
        RECT 147.640 11.750 148.640 12.130 ;
        RECT 58.680 9.640 59.680 10.640 ;
        RECT 81.640 9.640 82.640 10.640 ;
        RECT 143.680 9.990 144.680 10.370 ;
        RECT 147.640 9.990 148.640 10.370 ;
        RECT 143.680 9.110 144.680 9.490 ;
        RECT 147.640 9.110 148.640 9.490 ;
        RECT 54.720 6.040 55.720 7.040 ;
        RECT 85.600 6.040 86.600 7.040 ;
        RECT 143.680 6.470 144.680 6.850 ;
        RECT 147.640 6.470 148.640 6.850 ;
        RECT 143.680 4.710 144.680 5.090 ;
        RECT 147.640 4.710 148.640 5.090 ;
        RECT 61.600 4.000 62.600 4.380 ;
        RECT 78.720 4.000 79.720 4.380 ;
        RECT 143.680 3.830 144.680 4.210 ;
        RECT 147.640 3.830 148.640 4.210 ;
        RECT 143.680 2.950 144.680 3.330 ;
        RECT 147.640 2.950 148.640 3.330 ;
      LAYER via2 ;
        RECT 24.640 221.810 24.960 222.130 ;
        RECT 25.200 221.810 25.520 222.130 ;
        RECT 24.640 221.250 24.960 221.570 ;
        RECT 25.200 221.250 25.520 221.570 ;
        RECT 27.600 221.810 27.920 222.130 ;
        RECT 28.160 221.810 28.480 222.130 ;
        RECT 27.600 221.250 27.920 221.570 ;
        RECT 28.160 221.250 28.480 221.570 ;
        RECT 49.840 221.810 50.160 222.130 ;
        RECT 50.400 221.810 50.720 222.130 ;
        RECT 49.840 221.250 50.160 221.570 ;
        RECT 50.400 221.250 50.720 221.570 ;
        RECT 52.800 221.810 53.120 222.130 ;
        RECT 53.360 221.810 53.680 222.130 ;
        RECT 52.800 221.250 53.120 221.570 ;
        RECT 53.360 221.250 53.680 221.570 ;
        RECT 75.040 221.810 75.360 222.130 ;
        RECT 75.600 221.810 75.920 222.130 ;
        RECT 75.040 221.250 75.360 221.570 ;
        RECT 75.600 221.250 75.920 221.570 ;
        RECT 78.000 221.810 78.320 222.130 ;
        RECT 78.560 221.810 78.880 222.130 ;
        RECT 78.000 221.250 78.320 221.570 ;
        RECT 78.560 221.250 78.880 221.570 ;
        RECT 100.240 221.810 100.560 222.130 ;
        RECT 100.800 221.810 101.120 222.130 ;
        RECT 100.240 221.250 100.560 221.570 ;
        RECT 100.800 221.250 101.120 221.570 ;
        RECT 103.200 221.810 103.520 222.130 ;
        RECT 103.760 221.810 104.080 222.130 ;
        RECT 143.740 222.100 144.060 222.420 ;
        RECT 144.300 222.100 144.620 222.420 ;
        RECT 147.700 222.100 148.020 222.420 ;
        RECT 148.260 222.100 148.580 222.420 ;
        RECT 103.200 221.250 103.520 221.570 ;
        RECT 103.760 221.250 104.080 221.570 ;
        RECT 143.740 221.220 144.060 221.540 ;
        RECT 144.300 221.220 144.620 221.540 ;
        RECT 147.700 221.220 148.020 221.540 ;
        RECT 148.260 221.220 148.580 221.540 ;
        RECT 143.740 219.460 144.060 219.780 ;
        RECT 144.300 219.460 144.620 219.780 ;
        RECT 147.700 219.460 148.020 219.780 ;
        RECT 148.260 219.460 148.580 219.780 ;
        RECT 21.760 218.210 22.080 218.530 ;
        RECT 22.320 218.210 22.640 218.530 ;
        RECT 21.760 217.650 22.080 217.970 ;
        RECT 22.320 217.650 22.640 217.970 ;
        RECT 30.480 218.210 30.800 218.530 ;
        RECT 31.040 218.210 31.360 218.530 ;
        RECT 30.480 217.650 30.800 217.970 ;
        RECT 31.040 217.650 31.360 217.970 ;
        RECT 46.960 218.210 47.280 218.530 ;
        RECT 47.520 218.210 47.840 218.530 ;
        RECT 46.960 217.650 47.280 217.970 ;
        RECT 47.520 217.650 47.840 217.970 ;
        RECT 55.680 218.210 56.000 218.530 ;
        RECT 56.240 218.210 56.560 218.530 ;
        RECT 55.680 217.650 56.000 217.970 ;
        RECT 56.240 217.650 56.560 217.970 ;
        RECT 72.160 218.210 72.480 218.530 ;
        RECT 72.720 218.210 73.040 218.530 ;
        RECT 72.160 217.650 72.480 217.970 ;
        RECT 72.720 217.650 73.040 217.970 ;
        RECT 80.880 218.210 81.200 218.530 ;
        RECT 81.440 218.210 81.760 218.530 ;
        RECT 80.880 217.650 81.200 217.970 ;
        RECT 81.440 217.650 81.760 217.970 ;
        RECT 97.360 218.210 97.680 218.530 ;
        RECT 97.920 218.210 98.240 218.530 ;
        RECT 97.360 217.650 97.680 217.970 ;
        RECT 97.920 217.650 98.240 217.970 ;
        RECT 106.080 218.210 106.400 218.530 ;
        RECT 106.640 218.210 106.960 218.530 ;
        RECT 106.080 217.650 106.400 217.970 ;
        RECT 106.640 217.650 106.960 217.970 ;
        RECT 122.560 218.210 122.880 218.530 ;
        RECT 123.120 218.210 123.440 218.530 ;
        RECT 122.560 217.650 122.880 217.970 ;
        RECT 123.120 217.650 123.440 217.970 ;
        RECT 17.800 214.610 18.120 214.930 ;
        RECT 18.360 214.610 18.680 214.930 ;
        RECT 17.800 214.050 18.120 214.370 ;
        RECT 18.360 214.050 18.680 214.370 ;
        RECT 34.440 214.610 34.760 214.930 ;
        RECT 35.000 214.610 35.320 214.930 ;
        RECT 34.440 214.050 34.760 214.370 ;
        RECT 35.000 214.050 35.320 214.370 ;
        RECT 43.000 214.610 43.320 214.930 ;
        RECT 43.560 214.610 43.880 214.930 ;
        RECT 43.000 214.050 43.320 214.370 ;
        RECT 43.560 214.050 43.880 214.370 ;
        RECT 59.640 214.610 59.960 214.930 ;
        RECT 60.200 214.610 60.520 214.930 ;
        RECT 59.640 214.050 59.960 214.370 ;
        RECT 60.200 214.050 60.520 214.370 ;
        RECT 68.200 214.610 68.520 214.930 ;
        RECT 68.760 214.610 69.080 214.930 ;
        RECT 68.200 214.050 68.520 214.370 ;
        RECT 68.760 214.050 69.080 214.370 ;
        RECT 84.840 214.610 85.160 214.930 ;
        RECT 85.400 214.610 85.720 214.930 ;
        RECT 84.840 214.050 85.160 214.370 ;
        RECT 85.400 214.050 85.720 214.370 ;
        RECT 93.400 214.610 93.720 214.930 ;
        RECT 93.960 214.610 94.280 214.930 ;
        RECT 93.400 214.050 93.720 214.370 ;
        RECT 93.960 214.050 94.280 214.370 ;
        RECT 110.040 214.610 110.360 214.930 ;
        RECT 110.600 214.610 110.920 214.930 ;
        RECT 110.040 214.050 110.360 214.370 ;
        RECT 110.600 214.050 110.920 214.370 ;
        RECT 118.600 214.610 118.920 214.930 ;
        RECT 119.160 214.610 119.480 214.930 ;
        RECT 118.600 214.050 118.920 214.370 ;
        RECT 119.160 214.050 119.480 214.370 ;
        RECT 147.700 215.940 148.020 216.260 ;
        RECT 148.260 215.940 148.580 216.260 ;
        RECT 147.700 215.060 148.020 215.380 ;
        RECT 148.260 215.060 148.580 215.380 ;
        RECT 143.740 214.180 144.060 214.500 ;
        RECT 144.300 214.180 144.620 214.500 ;
        RECT 17.800 210.830 18.120 211.150 ;
        RECT 18.360 210.830 18.680 211.150 ;
        RECT 21.760 210.830 22.080 211.150 ;
        RECT 22.320 210.830 22.640 211.150 ;
        RECT 30.480 210.830 30.800 211.150 ;
        RECT 31.040 210.830 31.360 211.150 ;
        RECT 34.440 210.830 34.760 211.150 ;
        RECT 35.000 210.830 35.320 211.150 ;
        RECT 43.000 210.830 43.320 211.150 ;
        RECT 43.560 210.830 43.880 211.150 ;
        RECT 46.960 210.830 47.280 211.150 ;
        RECT 47.520 210.830 47.840 211.150 ;
        RECT 55.680 210.830 56.000 211.150 ;
        RECT 56.240 210.830 56.560 211.150 ;
        RECT 59.640 210.830 59.960 211.150 ;
        RECT 60.200 210.830 60.520 211.150 ;
        RECT 68.200 210.830 68.520 211.150 ;
        RECT 68.760 210.830 69.080 211.150 ;
        RECT 72.160 210.830 72.480 211.150 ;
        RECT 72.720 210.830 73.040 211.150 ;
        RECT 80.880 210.830 81.200 211.150 ;
        RECT 81.440 210.830 81.760 211.150 ;
        RECT 84.840 210.830 85.160 211.150 ;
        RECT 85.400 210.830 85.720 211.150 ;
        RECT 93.400 210.830 93.720 211.150 ;
        RECT 93.960 210.830 94.280 211.150 ;
        RECT 97.360 210.830 97.680 211.150 ;
        RECT 97.920 210.830 98.240 211.150 ;
        RECT 106.080 210.830 106.400 211.150 ;
        RECT 106.640 210.830 106.960 211.150 ;
        RECT 110.040 210.830 110.360 211.150 ;
        RECT 110.600 210.830 110.920 211.150 ;
        RECT 143.740 210.660 144.060 210.980 ;
        RECT 144.300 210.660 144.620 210.980 ;
        RECT 147.700 210.660 148.020 210.980 ;
        RECT 148.260 210.660 148.580 210.980 ;
        RECT 17.800 209.950 18.120 210.270 ;
        RECT 18.360 209.950 18.680 210.270 ;
        RECT 21.760 209.950 22.080 210.270 ;
        RECT 22.320 209.950 22.640 210.270 ;
        RECT 30.480 209.950 30.800 210.270 ;
        RECT 31.040 209.950 31.360 210.270 ;
        RECT 34.440 209.950 34.760 210.270 ;
        RECT 35.000 209.950 35.320 210.270 ;
        RECT 43.000 209.950 43.320 210.270 ;
        RECT 43.560 209.950 43.880 210.270 ;
        RECT 46.960 209.950 47.280 210.270 ;
        RECT 47.520 209.950 47.840 210.270 ;
        RECT 55.680 209.950 56.000 210.270 ;
        RECT 56.240 209.950 56.560 210.270 ;
        RECT 59.640 209.950 59.960 210.270 ;
        RECT 60.200 209.950 60.520 210.270 ;
        RECT 68.200 209.950 68.520 210.270 ;
        RECT 68.760 209.950 69.080 210.270 ;
        RECT 72.160 209.950 72.480 210.270 ;
        RECT 72.720 209.950 73.040 210.270 ;
        RECT 80.880 209.950 81.200 210.270 ;
        RECT 81.440 209.950 81.760 210.270 ;
        RECT 84.840 209.950 85.160 210.270 ;
        RECT 85.400 209.950 85.720 210.270 ;
        RECT 93.400 209.950 93.720 210.270 ;
        RECT 93.960 209.950 94.280 210.270 ;
        RECT 97.360 209.950 97.680 210.270 ;
        RECT 97.920 209.950 98.240 210.270 ;
        RECT 106.080 209.950 106.400 210.270 ;
        RECT 106.640 209.950 106.960 210.270 ;
        RECT 110.040 209.950 110.360 210.270 ;
        RECT 110.600 209.950 110.920 210.270 ;
        RECT 17.800 208.190 18.120 208.510 ;
        RECT 18.360 208.190 18.680 208.510 ;
        RECT 21.760 208.190 22.080 208.510 ;
        RECT 22.320 208.190 22.640 208.510 ;
        RECT 17.800 207.310 18.120 207.630 ;
        RECT 18.360 207.310 18.680 207.630 ;
        RECT 30.480 208.190 30.800 208.510 ;
        RECT 31.040 208.190 31.360 208.510 ;
        RECT 34.440 208.190 34.760 208.510 ;
        RECT 35.000 208.190 35.320 208.510 ;
        RECT 43.000 208.190 43.320 208.510 ;
        RECT 43.560 208.190 43.880 208.510 ;
        RECT 46.960 208.190 47.280 208.510 ;
        RECT 47.520 208.190 47.840 208.510 ;
        RECT 34.440 207.310 34.760 207.630 ;
        RECT 35.000 207.310 35.320 207.630 ;
        RECT 43.000 207.310 43.320 207.630 ;
        RECT 43.560 207.310 43.880 207.630 ;
        RECT 55.680 208.190 56.000 208.510 ;
        RECT 56.240 208.190 56.560 208.510 ;
        RECT 59.640 208.190 59.960 208.510 ;
        RECT 60.200 208.190 60.520 208.510 ;
        RECT 68.200 208.190 68.520 208.510 ;
        RECT 68.760 208.190 69.080 208.510 ;
        RECT 72.160 208.190 72.480 208.510 ;
        RECT 72.720 208.190 73.040 208.510 ;
        RECT 59.640 207.310 59.960 207.630 ;
        RECT 60.200 207.310 60.520 207.630 ;
        RECT 68.200 207.310 68.520 207.630 ;
        RECT 68.760 207.310 69.080 207.630 ;
        RECT 80.880 208.190 81.200 208.510 ;
        RECT 81.440 208.190 81.760 208.510 ;
        RECT 84.840 208.190 85.160 208.510 ;
        RECT 85.400 208.190 85.720 208.510 ;
        RECT 93.400 208.190 93.720 208.510 ;
        RECT 93.960 208.190 94.280 208.510 ;
        RECT 97.360 208.190 97.680 208.510 ;
        RECT 97.920 208.190 98.240 208.510 ;
        RECT 84.840 207.310 85.160 207.630 ;
        RECT 85.400 207.310 85.720 207.630 ;
        RECT 93.400 207.310 93.720 207.630 ;
        RECT 93.960 207.310 94.280 207.630 ;
        RECT 118.600 209.070 118.920 209.390 ;
        RECT 119.160 209.070 119.480 209.390 ;
        RECT 122.560 209.070 122.880 209.390 ;
        RECT 123.120 209.070 123.440 209.390 ;
        RECT 106.080 208.190 106.400 208.510 ;
        RECT 106.640 208.190 106.960 208.510 ;
        RECT 110.040 208.190 110.360 208.510 ;
        RECT 110.600 208.190 110.920 208.510 ;
        RECT 110.040 207.310 110.360 207.630 ;
        RECT 110.600 207.310 110.920 207.630 ;
        RECT 143.740 208.900 144.060 209.220 ;
        RECT 144.300 208.900 144.620 209.220 ;
        RECT 147.700 208.900 148.020 209.220 ;
        RECT 148.260 208.900 148.580 209.220 ;
        RECT 118.600 208.190 118.920 208.510 ;
        RECT 119.160 208.190 119.480 208.510 ;
        RECT 122.560 208.190 122.880 208.510 ;
        RECT 123.120 208.190 123.440 208.510 ;
        RECT 118.600 206.430 118.920 206.750 ;
        RECT 119.160 206.430 119.480 206.750 ;
        RECT 122.560 206.430 122.880 206.750 ;
        RECT 123.120 206.430 123.440 206.750 ;
        RECT 118.600 205.550 118.920 205.870 ;
        RECT 119.160 205.550 119.480 205.870 ;
        RECT 143.740 205.380 144.060 205.700 ;
        RECT 144.300 205.380 144.620 205.700 ;
        RECT 147.700 205.380 148.020 205.700 ;
        RECT 148.260 205.380 148.580 205.700 ;
        RECT 17.800 204.670 18.120 204.990 ;
        RECT 18.360 204.670 18.680 204.990 ;
        RECT 21.760 204.670 22.080 204.990 ;
        RECT 22.320 204.670 22.640 204.990 ;
        RECT 30.480 204.670 30.800 204.990 ;
        RECT 31.040 204.670 31.360 204.990 ;
        RECT 34.440 204.670 34.760 204.990 ;
        RECT 35.000 204.670 35.320 204.990 ;
        RECT 43.000 204.670 43.320 204.990 ;
        RECT 43.560 204.670 43.880 204.990 ;
        RECT 46.960 204.670 47.280 204.990 ;
        RECT 47.520 204.670 47.840 204.990 ;
        RECT 55.680 204.670 56.000 204.990 ;
        RECT 56.240 204.670 56.560 204.990 ;
        RECT 59.640 204.670 59.960 204.990 ;
        RECT 60.200 204.670 60.520 204.990 ;
        RECT 68.200 204.670 68.520 204.990 ;
        RECT 68.760 204.670 69.080 204.990 ;
        RECT 72.160 204.670 72.480 204.990 ;
        RECT 72.720 204.670 73.040 204.990 ;
        RECT 80.880 204.670 81.200 204.990 ;
        RECT 81.440 204.670 81.760 204.990 ;
        RECT 84.840 204.670 85.160 204.990 ;
        RECT 85.400 204.670 85.720 204.990 ;
        RECT 93.400 204.670 93.720 204.990 ;
        RECT 93.960 204.670 94.280 204.990 ;
        RECT 97.360 204.670 97.680 204.990 ;
        RECT 97.920 204.670 98.240 204.990 ;
        RECT 106.080 204.670 106.400 204.990 ;
        RECT 106.640 204.670 106.960 204.990 ;
        RECT 110.040 204.670 110.360 204.990 ;
        RECT 110.600 204.670 110.920 204.990 ;
        RECT 17.800 202.910 18.120 203.230 ;
        RECT 18.360 202.910 18.680 203.230 ;
        RECT 21.760 202.910 22.080 203.230 ;
        RECT 22.320 202.910 22.640 203.230 ;
        RECT 30.480 202.910 30.800 203.230 ;
        RECT 31.040 202.910 31.360 203.230 ;
        RECT 34.440 202.910 34.760 203.230 ;
        RECT 35.000 202.910 35.320 203.230 ;
        RECT 43.000 202.910 43.320 203.230 ;
        RECT 43.560 202.910 43.880 203.230 ;
        RECT 46.960 202.910 47.280 203.230 ;
        RECT 47.520 202.910 47.840 203.230 ;
        RECT 55.680 202.910 56.000 203.230 ;
        RECT 56.240 202.910 56.560 203.230 ;
        RECT 59.640 202.910 59.960 203.230 ;
        RECT 60.200 202.910 60.520 203.230 ;
        RECT 68.200 202.910 68.520 203.230 ;
        RECT 68.760 202.910 69.080 203.230 ;
        RECT 72.160 202.910 72.480 203.230 ;
        RECT 72.720 202.910 73.040 203.230 ;
        RECT 80.880 202.910 81.200 203.230 ;
        RECT 81.440 202.910 81.760 203.230 ;
        RECT 84.840 202.910 85.160 203.230 ;
        RECT 85.400 202.910 85.720 203.230 ;
        RECT 93.400 202.910 93.720 203.230 ;
        RECT 93.960 202.910 94.280 203.230 ;
        RECT 97.360 202.910 97.680 203.230 ;
        RECT 97.920 202.910 98.240 203.230 ;
        RECT 106.080 202.910 106.400 203.230 ;
        RECT 106.640 202.910 106.960 203.230 ;
        RECT 110.040 202.910 110.360 203.230 ;
        RECT 110.600 202.910 110.920 203.230 ;
        RECT 118.600 202.910 118.920 203.230 ;
        RECT 119.160 202.910 119.480 203.230 ;
        RECT 122.560 202.910 122.880 203.230 ;
        RECT 123.120 202.910 123.440 203.230 ;
        RECT 21.760 202.030 22.080 202.350 ;
        RECT 22.320 202.030 22.640 202.350 ;
        RECT 30.480 202.030 30.800 202.350 ;
        RECT 31.040 202.030 31.360 202.350 ;
        RECT 46.960 202.030 47.280 202.350 ;
        RECT 47.520 202.030 47.840 202.350 ;
        RECT 55.680 202.030 56.000 202.350 ;
        RECT 56.240 202.030 56.560 202.350 ;
        RECT 72.160 202.030 72.480 202.350 ;
        RECT 72.720 202.030 73.040 202.350 ;
        RECT 80.880 202.030 81.200 202.350 ;
        RECT 81.440 202.030 81.760 202.350 ;
        RECT 97.360 202.030 97.680 202.350 ;
        RECT 97.920 202.030 98.240 202.350 ;
        RECT 106.080 202.030 106.400 202.350 ;
        RECT 106.640 202.030 106.960 202.350 ;
        RECT 122.560 202.030 122.880 202.350 ;
        RECT 123.120 202.030 123.440 202.350 ;
        RECT 17.800 199.390 18.120 199.710 ;
        RECT 18.360 199.390 18.680 199.710 ;
        RECT 21.760 199.390 22.080 199.710 ;
        RECT 22.320 199.390 22.640 199.710 ;
        RECT 30.480 199.390 30.800 199.710 ;
        RECT 31.040 199.390 31.360 199.710 ;
        RECT 34.440 199.390 34.760 199.710 ;
        RECT 35.000 199.390 35.320 199.710 ;
        RECT 43.000 199.390 43.320 199.710 ;
        RECT 43.560 199.390 43.880 199.710 ;
        RECT 46.960 199.390 47.280 199.710 ;
        RECT 47.520 199.390 47.840 199.710 ;
        RECT 55.680 199.390 56.000 199.710 ;
        RECT 56.240 199.390 56.560 199.710 ;
        RECT 59.640 199.390 59.960 199.710 ;
        RECT 60.200 199.390 60.520 199.710 ;
        RECT 68.200 199.390 68.520 199.710 ;
        RECT 68.760 199.390 69.080 199.710 ;
        RECT 72.160 199.390 72.480 199.710 ;
        RECT 72.720 199.390 73.040 199.710 ;
        RECT 80.880 199.390 81.200 199.710 ;
        RECT 81.440 199.390 81.760 199.710 ;
        RECT 84.840 199.390 85.160 199.710 ;
        RECT 85.400 199.390 85.720 199.710 ;
        RECT 93.400 199.390 93.720 199.710 ;
        RECT 93.960 199.390 94.280 199.710 ;
        RECT 97.360 199.390 97.680 199.710 ;
        RECT 97.920 199.390 98.240 199.710 ;
        RECT 106.080 199.390 106.400 199.710 ;
        RECT 106.640 199.390 106.960 199.710 ;
        RECT 110.040 199.390 110.360 199.710 ;
        RECT 110.600 199.390 110.920 199.710 ;
        RECT 118.600 199.390 118.920 199.710 ;
        RECT 119.160 199.390 119.480 199.710 ;
        RECT 122.560 199.390 122.880 199.710 ;
        RECT 123.120 199.390 123.440 199.710 ;
        RECT 17.800 197.630 18.120 197.950 ;
        RECT 18.360 197.630 18.680 197.950 ;
        RECT 21.760 197.630 22.080 197.950 ;
        RECT 22.320 197.630 22.640 197.950 ;
        RECT 30.480 197.630 30.800 197.950 ;
        RECT 31.040 197.630 31.360 197.950 ;
        RECT 34.440 197.630 34.760 197.950 ;
        RECT 35.000 197.630 35.320 197.950 ;
        RECT 43.000 197.630 43.320 197.950 ;
        RECT 43.560 197.630 43.880 197.950 ;
        RECT 46.960 197.630 47.280 197.950 ;
        RECT 47.520 197.630 47.840 197.950 ;
        RECT 55.680 197.630 56.000 197.950 ;
        RECT 56.240 197.630 56.560 197.950 ;
        RECT 59.640 197.630 59.960 197.950 ;
        RECT 60.200 197.630 60.520 197.950 ;
        RECT 68.200 197.630 68.520 197.950 ;
        RECT 68.760 197.630 69.080 197.950 ;
        RECT 72.160 197.630 72.480 197.950 ;
        RECT 72.720 197.630 73.040 197.950 ;
        RECT 80.880 197.630 81.200 197.950 ;
        RECT 81.440 197.630 81.760 197.950 ;
        RECT 84.840 197.630 85.160 197.950 ;
        RECT 85.400 197.630 85.720 197.950 ;
        RECT 93.400 197.630 93.720 197.950 ;
        RECT 93.960 197.630 94.280 197.950 ;
        RECT 97.360 197.630 97.680 197.950 ;
        RECT 97.920 197.630 98.240 197.950 ;
        RECT 106.080 197.630 106.400 197.950 ;
        RECT 106.640 197.630 106.960 197.950 ;
        RECT 110.040 197.630 110.360 197.950 ;
        RECT 110.600 197.630 110.920 197.950 ;
        RECT 118.600 197.630 118.920 197.950 ;
        RECT 119.160 197.630 119.480 197.950 ;
        RECT 122.560 197.630 122.880 197.950 ;
        RECT 123.120 197.630 123.440 197.950 ;
        RECT 17.800 195.870 18.120 196.190 ;
        RECT 18.360 195.870 18.680 196.190 ;
        RECT 21.760 195.870 22.080 196.190 ;
        RECT 22.320 195.870 22.640 196.190 ;
        RECT 30.480 195.870 30.800 196.190 ;
        RECT 31.040 195.870 31.360 196.190 ;
        RECT 34.440 195.870 34.760 196.190 ;
        RECT 35.000 195.870 35.320 196.190 ;
        RECT 43.000 195.870 43.320 196.190 ;
        RECT 43.560 195.870 43.880 196.190 ;
        RECT 46.960 195.870 47.280 196.190 ;
        RECT 47.520 195.870 47.840 196.190 ;
        RECT 55.680 195.870 56.000 196.190 ;
        RECT 56.240 195.870 56.560 196.190 ;
        RECT 59.640 195.870 59.960 196.190 ;
        RECT 60.200 195.870 60.520 196.190 ;
        RECT 68.200 195.870 68.520 196.190 ;
        RECT 68.760 195.870 69.080 196.190 ;
        RECT 72.160 195.870 72.480 196.190 ;
        RECT 72.720 195.870 73.040 196.190 ;
        RECT 80.880 195.870 81.200 196.190 ;
        RECT 81.440 195.870 81.760 196.190 ;
        RECT 84.840 195.870 85.160 196.190 ;
        RECT 85.400 195.870 85.720 196.190 ;
        RECT 93.400 195.870 93.720 196.190 ;
        RECT 93.960 195.870 94.280 196.190 ;
        RECT 97.360 195.870 97.680 196.190 ;
        RECT 97.920 195.870 98.240 196.190 ;
        RECT 106.080 195.870 106.400 196.190 ;
        RECT 106.640 195.870 106.960 196.190 ;
        RECT 110.040 195.870 110.360 196.190 ;
        RECT 110.600 195.870 110.920 196.190 ;
        RECT 143.740 201.860 144.060 202.180 ;
        RECT 144.300 201.860 144.620 202.180 ;
        RECT 147.700 201.860 148.020 202.180 ;
        RECT 148.260 201.860 148.580 202.180 ;
        RECT 143.740 200.100 144.060 200.420 ;
        RECT 144.300 200.100 144.620 200.420 ;
        RECT 147.700 200.100 148.020 200.420 ;
        RECT 148.260 200.100 148.580 200.420 ;
        RECT 147.700 199.220 148.020 199.540 ;
        RECT 148.260 199.220 148.580 199.540 ;
        RECT 143.740 196.580 144.060 196.900 ;
        RECT 144.300 196.580 144.620 196.900 ;
        RECT 147.700 196.580 148.020 196.900 ;
        RECT 148.260 196.580 148.580 196.900 ;
        RECT 143.740 194.820 144.060 195.140 ;
        RECT 144.300 194.820 144.620 195.140 ;
        RECT 147.700 194.820 148.020 195.140 ;
        RECT 148.260 194.820 148.580 195.140 ;
        RECT 17.800 192.350 18.120 192.670 ;
        RECT 18.360 192.350 18.680 192.670 ;
        RECT 21.760 192.350 22.080 192.670 ;
        RECT 22.320 192.350 22.640 192.670 ;
        RECT 30.480 192.350 30.800 192.670 ;
        RECT 31.040 192.350 31.360 192.670 ;
        RECT 34.440 192.350 34.760 192.670 ;
        RECT 35.000 192.350 35.320 192.670 ;
        RECT 43.000 192.350 43.320 192.670 ;
        RECT 43.560 192.350 43.880 192.670 ;
        RECT 46.960 192.350 47.280 192.670 ;
        RECT 47.520 192.350 47.840 192.670 ;
        RECT 55.680 192.350 56.000 192.670 ;
        RECT 56.240 192.350 56.560 192.670 ;
        RECT 59.640 192.350 59.960 192.670 ;
        RECT 60.200 192.350 60.520 192.670 ;
        RECT 68.200 192.350 68.520 192.670 ;
        RECT 68.760 192.350 69.080 192.670 ;
        RECT 72.160 192.350 72.480 192.670 ;
        RECT 72.720 192.350 73.040 192.670 ;
        RECT 80.880 192.350 81.200 192.670 ;
        RECT 81.440 192.350 81.760 192.670 ;
        RECT 84.840 192.350 85.160 192.670 ;
        RECT 85.400 192.350 85.720 192.670 ;
        RECT 93.400 192.350 93.720 192.670 ;
        RECT 93.960 192.350 94.280 192.670 ;
        RECT 97.360 192.350 97.680 192.670 ;
        RECT 97.920 192.350 98.240 192.670 ;
        RECT 106.080 192.350 106.400 192.670 ;
        RECT 106.640 192.350 106.960 192.670 ;
        RECT 110.040 192.350 110.360 192.670 ;
        RECT 110.600 192.350 110.920 192.670 ;
        RECT 17.800 191.470 18.120 191.790 ;
        RECT 18.360 191.470 18.680 191.790 ;
        RECT 21.760 191.470 22.080 191.790 ;
        RECT 22.320 191.470 22.640 191.790 ;
        RECT 30.480 191.470 30.800 191.790 ;
        RECT 31.040 191.470 31.360 191.790 ;
        RECT 34.440 191.470 34.760 191.790 ;
        RECT 35.000 191.470 35.320 191.790 ;
        RECT 43.000 191.470 43.320 191.790 ;
        RECT 43.560 191.470 43.880 191.790 ;
        RECT 46.960 191.470 47.280 191.790 ;
        RECT 47.520 191.470 47.840 191.790 ;
        RECT 55.680 191.470 56.000 191.790 ;
        RECT 56.240 191.470 56.560 191.790 ;
        RECT 59.640 191.470 59.960 191.790 ;
        RECT 60.200 191.470 60.520 191.790 ;
        RECT 68.200 191.470 68.520 191.790 ;
        RECT 68.760 191.470 69.080 191.790 ;
        RECT 72.160 191.470 72.480 191.790 ;
        RECT 72.720 191.470 73.040 191.790 ;
        RECT 80.880 191.470 81.200 191.790 ;
        RECT 81.440 191.470 81.760 191.790 ;
        RECT 84.840 191.470 85.160 191.790 ;
        RECT 85.400 191.470 85.720 191.790 ;
        RECT 93.400 191.470 93.720 191.790 ;
        RECT 93.960 191.470 94.280 191.790 ;
        RECT 97.360 191.470 97.680 191.790 ;
        RECT 97.920 191.470 98.240 191.790 ;
        RECT 106.080 191.470 106.400 191.790 ;
        RECT 106.640 191.470 106.960 191.790 ;
        RECT 110.040 191.470 110.360 191.790 ;
        RECT 110.600 191.470 110.920 191.790 ;
        RECT 17.800 188.830 18.120 189.150 ;
        RECT 18.360 188.830 18.680 189.150 ;
        RECT 34.440 188.830 34.760 189.150 ;
        RECT 35.000 188.830 35.320 189.150 ;
        RECT 43.000 188.830 43.320 189.150 ;
        RECT 43.560 188.830 43.880 189.150 ;
        RECT 59.640 188.830 59.960 189.150 ;
        RECT 60.200 188.830 60.520 189.150 ;
        RECT 68.200 188.830 68.520 189.150 ;
        RECT 68.760 188.830 69.080 189.150 ;
        RECT 84.840 188.830 85.160 189.150 ;
        RECT 85.400 188.830 85.720 189.150 ;
        RECT 93.400 188.830 93.720 189.150 ;
        RECT 93.960 188.830 94.280 189.150 ;
        RECT 110.040 188.830 110.360 189.150 ;
        RECT 110.600 188.830 110.920 189.150 ;
        RECT 147.700 191.300 148.020 191.620 ;
        RECT 148.260 191.300 148.580 191.620 ;
        RECT 147.700 190.420 148.020 190.740 ;
        RECT 148.260 190.420 148.580 190.740 ;
        RECT 143.740 189.540 144.060 189.860 ;
        RECT 144.300 189.540 144.620 189.860 ;
        RECT 17.800 187.950 18.120 188.270 ;
        RECT 18.360 187.950 18.680 188.270 ;
        RECT 17.800 185.310 18.120 185.630 ;
        RECT 18.360 185.310 18.680 185.630 ;
        RECT 34.440 187.950 34.760 188.270 ;
        RECT 35.000 187.950 35.320 188.270 ;
        RECT 43.000 187.950 43.320 188.270 ;
        RECT 43.560 187.950 43.880 188.270 ;
        RECT 24.640 185.020 24.960 185.340 ;
        RECT 25.200 185.020 25.520 185.340 ;
        RECT 17.800 184.430 18.120 184.750 ;
        RECT 18.360 184.430 18.680 184.750 ;
        RECT 24.640 184.460 24.960 184.780 ;
        RECT 25.200 184.460 25.520 184.780 ;
        RECT 27.600 185.020 27.920 185.340 ;
        RECT 28.160 185.020 28.480 185.340 ;
        RECT 34.440 185.310 34.760 185.630 ;
        RECT 35.000 185.310 35.320 185.630 ;
        RECT 43.000 185.310 43.320 185.630 ;
        RECT 43.560 185.310 43.880 185.630 ;
        RECT 59.640 187.950 59.960 188.270 ;
        RECT 60.200 187.950 60.520 188.270 ;
        RECT 68.200 187.950 68.520 188.270 ;
        RECT 68.760 187.950 69.080 188.270 ;
        RECT 49.840 185.020 50.160 185.340 ;
        RECT 50.400 185.020 50.720 185.340 ;
        RECT 27.600 184.460 27.920 184.780 ;
        RECT 28.160 184.460 28.480 184.780 ;
        RECT 34.440 184.430 34.760 184.750 ;
        RECT 35.000 184.430 35.320 184.750 ;
        RECT 43.000 184.430 43.320 184.750 ;
        RECT 43.560 184.430 43.880 184.750 ;
        RECT 49.840 184.460 50.160 184.780 ;
        RECT 50.400 184.460 50.720 184.780 ;
        RECT 52.800 185.020 53.120 185.340 ;
        RECT 53.360 185.020 53.680 185.340 ;
        RECT 59.640 185.310 59.960 185.630 ;
        RECT 60.200 185.310 60.520 185.630 ;
        RECT 68.200 185.310 68.520 185.630 ;
        RECT 68.760 185.310 69.080 185.630 ;
        RECT 84.840 187.950 85.160 188.270 ;
        RECT 85.400 187.950 85.720 188.270 ;
        RECT 93.400 187.950 93.720 188.270 ;
        RECT 93.960 187.950 94.280 188.270 ;
        RECT 75.040 185.020 75.360 185.340 ;
        RECT 75.600 185.020 75.920 185.340 ;
        RECT 52.800 184.460 53.120 184.780 ;
        RECT 53.360 184.460 53.680 184.780 ;
        RECT 59.640 184.430 59.960 184.750 ;
        RECT 60.200 184.430 60.520 184.750 ;
        RECT 68.200 184.430 68.520 184.750 ;
        RECT 68.760 184.430 69.080 184.750 ;
        RECT 75.040 184.460 75.360 184.780 ;
        RECT 75.600 184.460 75.920 184.780 ;
        RECT 78.000 185.020 78.320 185.340 ;
        RECT 78.560 185.020 78.880 185.340 ;
        RECT 84.840 185.310 85.160 185.630 ;
        RECT 85.400 185.310 85.720 185.630 ;
        RECT 93.400 185.310 93.720 185.630 ;
        RECT 93.960 185.310 94.280 185.630 ;
        RECT 110.040 187.950 110.360 188.270 ;
        RECT 110.600 187.950 110.920 188.270 ;
        RECT 100.240 185.020 100.560 185.340 ;
        RECT 100.800 185.020 101.120 185.340 ;
        RECT 78.000 184.460 78.320 184.780 ;
        RECT 78.560 184.460 78.880 184.780 ;
        RECT 84.840 184.430 85.160 184.750 ;
        RECT 85.400 184.430 85.720 184.750 ;
        RECT 93.400 184.430 93.720 184.750 ;
        RECT 93.960 184.430 94.280 184.750 ;
        RECT 100.240 184.460 100.560 184.780 ;
        RECT 100.800 184.460 101.120 184.780 ;
        RECT 103.200 185.020 103.520 185.340 ;
        RECT 103.760 185.020 104.080 185.340 ;
        RECT 122.560 186.190 122.880 186.510 ;
        RECT 123.120 186.190 123.440 186.510 ;
        RECT 143.740 186.020 144.060 186.340 ;
        RECT 144.300 186.020 144.620 186.340 ;
        RECT 147.700 186.020 148.020 186.340 ;
        RECT 148.260 186.020 148.580 186.340 ;
        RECT 110.040 185.310 110.360 185.630 ;
        RECT 110.600 185.310 110.920 185.630 ;
        RECT 118.600 185.310 118.920 185.630 ;
        RECT 119.160 185.310 119.480 185.630 ;
        RECT 103.200 184.460 103.520 184.780 ;
        RECT 103.760 184.460 104.080 184.780 ;
        RECT 110.040 184.430 110.360 184.750 ;
        RECT 110.600 184.430 110.920 184.750 ;
        RECT 122.560 184.430 122.880 184.750 ;
        RECT 123.120 184.430 123.440 184.750 ;
        RECT 20.940 182.910 21.260 183.230 ;
        RECT 20.940 182.350 21.260 182.670 ;
        RECT 17.800 181.790 18.120 182.110 ;
        RECT 18.360 181.790 18.680 182.110 ;
        RECT 31.860 182.910 32.180 183.230 ;
        RECT 31.860 182.350 32.180 182.670 ;
        RECT 46.140 182.910 46.460 183.230 ;
        RECT 46.140 182.350 46.460 182.670 ;
        RECT 34.440 181.790 34.760 182.110 ;
        RECT 35.000 181.790 35.320 182.110 ;
        RECT 43.000 181.790 43.320 182.110 ;
        RECT 43.560 181.790 43.880 182.110 ;
        RECT 57.060 182.910 57.380 183.230 ;
        RECT 57.060 182.350 57.380 182.670 ;
        RECT 71.340 182.910 71.660 183.230 ;
        RECT 71.340 182.350 71.660 182.670 ;
        RECT 59.640 181.790 59.960 182.110 ;
        RECT 60.200 181.790 60.520 182.110 ;
        RECT 68.200 181.790 68.520 182.110 ;
        RECT 68.760 181.790 69.080 182.110 ;
        RECT 82.260 182.910 82.580 183.230 ;
        RECT 82.260 182.350 82.580 182.670 ;
        RECT 96.540 182.910 96.860 183.230 ;
        RECT 96.540 182.350 96.860 182.670 ;
        RECT 84.840 181.790 85.160 182.110 ;
        RECT 85.400 181.790 85.720 182.110 ;
        RECT 93.400 181.790 93.720 182.110 ;
        RECT 93.960 181.790 94.280 182.110 ;
        RECT 143.740 184.260 144.060 184.580 ;
        RECT 144.300 184.260 144.620 184.580 ;
        RECT 147.700 184.260 148.020 184.580 ;
        RECT 148.260 184.260 148.580 184.580 ;
        RECT 107.460 182.910 107.780 183.230 ;
        RECT 107.460 182.350 107.780 182.670 ;
        RECT 117.220 182.230 117.540 182.550 ;
        RECT 117.780 182.230 118.100 182.550 ;
        RECT 110.040 181.790 110.360 182.110 ;
        RECT 110.600 181.790 110.920 182.110 ;
        RECT 122.560 181.790 122.880 182.110 ;
        RECT 123.120 181.790 123.440 182.110 ;
        RECT 17.800 180.910 18.120 181.230 ;
        RECT 18.360 180.910 18.680 181.230 ;
        RECT 17.800 178.270 18.120 178.590 ;
        RECT 18.360 178.270 18.680 178.590 ;
        RECT 34.440 180.910 34.760 181.230 ;
        RECT 35.000 180.910 35.320 181.230 ;
        RECT 43.000 180.910 43.320 181.230 ;
        RECT 43.560 180.910 43.880 181.230 ;
        RECT 24.640 177.980 24.960 178.300 ;
        RECT 25.200 177.980 25.520 178.300 ;
        RECT 17.800 177.390 18.120 177.710 ;
        RECT 18.360 177.390 18.680 177.710 ;
        RECT 24.640 177.420 24.960 177.740 ;
        RECT 25.200 177.420 25.520 177.740 ;
        RECT 27.600 177.980 27.920 178.300 ;
        RECT 28.160 177.980 28.480 178.300 ;
        RECT 34.440 178.270 34.760 178.590 ;
        RECT 35.000 178.270 35.320 178.590 ;
        RECT 43.000 178.270 43.320 178.590 ;
        RECT 43.560 178.270 43.880 178.590 ;
        RECT 59.640 180.910 59.960 181.230 ;
        RECT 60.200 180.910 60.520 181.230 ;
        RECT 68.200 180.910 68.520 181.230 ;
        RECT 68.760 180.910 69.080 181.230 ;
        RECT 49.840 177.980 50.160 178.300 ;
        RECT 50.400 177.980 50.720 178.300 ;
        RECT 27.600 177.420 27.920 177.740 ;
        RECT 28.160 177.420 28.480 177.740 ;
        RECT 34.440 177.390 34.760 177.710 ;
        RECT 35.000 177.390 35.320 177.710 ;
        RECT 43.000 177.390 43.320 177.710 ;
        RECT 43.560 177.390 43.880 177.710 ;
        RECT 49.840 177.420 50.160 177.740 ;
        RECT 50.400 177.420 50.720 177.740 ;
        RECT 52.800 177.980 53.120 178.300 ;
        RECT 53.360 177.980 53.680 178.300 ;
        RECT 59.640 178.270 59.960 178.590 ;
        RECT 60.200 178.270 60.520 178.590 ;
        RECT 68.200 178.270 68.520 178.590 ;
        RECT 68.760 178.270 69.080 178.590 ;
        RECT 84.840 180.910 85.160 181.230 ;
        RECT 85.400 180.910 85.720 181.230 ;
        RECT 93.400 180.910 93.720 181.230 ;
        RECT 93.960 180.910 94.280 181.230 ;
        RECT 75.040 177.980 75.360 178.300 ;
        RECT 75.600 177.980 75.920 178.300 ;
        RECT 52.800 177.420 53.120 177.740 ;
        RECT 53.360 177.420 53.680 177.740 ;
        RECT 59.640 177.390 59.960 177.710 ;
        RECT 60.200 177.390 60.520 177.710 ;
        RECT 68.200 177.390 68.520 177.710 ;
        RECT 68.760 177.390 69.080 177.710 ;
        RECT 75.040 177.420 75.360 177.740 ;
        RECT 75.600 177.420 75.920 177.740 ;
        RECT 78.000 177.980 78.320 178.300 ;
        RECT 78.560 177.980 78.880 178.300 ;
        RECT 84.840 178.270 85.160 178.590 ;
        RECT 85.400 178.270 85.720 178.590 ;
        RECT 93.400 178.270 93.720 178.590 ;
        RECT 93.960 178.270 94.280 178.590 ;
        RECT 110.040 180.910 110.360 181.230 ;
        RECT 110.600 180.910 110.920 181.230 ;
        RECT 122.560 180.910 122.880 181.230 ;
        RECT 123.120 180.910 123.440 181.230 ;
        RECT 100.240 177.980 100.560 178.300 ;
        RECT 100.800 177.980 101.120 178.300 ;
        RECT 78.000 177.420 78.320 177.740 ;
        RECT 78.560 177.420 78.880 177.740 ;
        RECT 84.840 177.390 85.160 177.710 ;
        RECT 85.400 177.390 85.720 177.710 ;
        RECT 93.400 177.390 93.720 177.710 ;
        RECT 93.960 177.390 94.280 177.710 ;
        RECT 100.240 177.420 100.560 177.740 ;
        RECT 100.800 177.420 101.120 177.740 ;
        RECT 103.200 177.980 103.520 178.300 ;
        RECT 103.760 177.980 104.080 178.300 ;
        RECT 143.740 180.740 144.060 181.060 ;
        RECT 144.300 180.740 144.620 181.060 ;
        RECT 147.700 180.740 148.020 181.060 ;
        RECT 148.260 180.740 148.580 181.060 ;
        RECT 110.040 178.270 110.360 178.590 ;
        RECT 110.600 178.270 110.920 178.590 ;
        RECT 122.560 178.270 122.880 178.590 ;
        RECT 123.120 178.270 123.440 178.590 ;
        RECT 103.200 177.420 103.520 177.740 ;
        RECT 103.760 177.420 104.080 177.740 ;
        RECT 110.040 177.390 110.360 177.710 ;
        RECT 110.600 177.390 110.920 177.710 ;
        RECT 122.560 177.390 122.880 177.710 ;
        RECT 123.120 177.390 123.440 177.710 ;
        RECT 20.065 175.870 20.385 176.190 ;
        RECT 20.065 175.310 20.385 175.630 ;
        RECT 17.800 174.750 18.120 175.070 ;
        RECT 18.360 174.750 18.680 175.070 ;
        RECT 32.735 175.870 33.055 176.190 ;
        RECT 32.735 175.310 33.055 175.630 ;
        RECT 45.265 175.870 45.585 176.190 ;
        RECT 45.265 175.310 45.585 175.630 ;
        RECT 34.440 174.750 34.760 175.070 ;
        RECT 35.000 174.750 35.320 175.070 ;
        RECT 43.000 174.750 43.320 175.070 ;
        RECT 43.560 174.750 43.880 175.070 ;
        RECT 57.935 175.870 58.255 176.190 ;
        RECT 57.935 175.310 58.255 175.630 ;
        RECT 70.465 175.870 70.785 176.190 ;
        RECT 70.465 175.310 70.785 175.630 ;
        RECT 59.640 174.750 59.960 175.070 ;
        RECT 60.200 174.750 60.520 175.070 ;
        RECT 68.200 174.750 68.520 175.070 ;
        RECT 68.760 174.750 69.080 175.070 ;
        RECT 83.135 175.870 83.455 176.190 ;
        RECT 83.135 175.310 83.455 175.630 ;
        RECT 95.665 175.870 95.985 176.190 ;
        RECT 95.665 175.310 95.985 175.630 ;
        RECT 84.840 174.750 85.160 175.070 ;
        RECT 85.400 174.750 85.720 175.070 ;
        RECT 93.400 174.750 93.720 175.070 ;
        RECT 93.960 174.750 94.280 175.070 ;
        RECT 124.720 176.950 125.040 177.270 ;
        RECT 125.280 176.950 125.600 177.270 ;
        RECT 143.740 177.220 144.060 177.540 ;
        RECT 144.300 177.220 144.620 177.540 ;
        RECT 147.700 177.220 148.020 177.540 ;
        RECT 148.260 177.220 148.580 177.540 ;
        RECT 108.335 175.870 108.655 176.190 ;
        RECT 108.335 175.310 108.655 175.630 ;
        RECT 143.740 175.460 144.060 175.780 ;
        RECT 144.300 175.460 144.620 175.780 ;
        RECT 147.700 175.460 148.020 175.780 ;
        RECT 148.260 175.460 148.580 175.780 ;
        RECT 110.040 174.750 110.360 175.070 ;
        RECT 110.600 174.750 110.920 175.070 ;
        RECT 122.560 174.750 122.880 175.070 ;
        RECT 123.120 174.750 123.440 175.070 ;
        RECT 147.700 174.580 148.020 174.900 ;
        RECT 148.260 174.580 148.580 174.900 ;
        RECT 17.800 173.870 18.120 174.190 ;
        RECT 18.360 173.870 18.680 174.190 ;
        RECT 17.800 171.230 18.120 171.550 ;
        RECT 18.360 171.230 18.680 171.550 ;
        RECT 34.440 173.870 34.760 174.190 ;
        RECT 35.000 173.870 35.320 174.190 ;
        RECT 43.000 173.870 43.320 174.190 ;
        RECT 43.560 173.870 43.880 174.190 ;
        RECT 24.640 170.940 24.960 171.260 ;
        RECT 25.200 170.940 25.520 171.260 ;
        RECT 17.800 170.350 18.120 170.670 ;
        RECT 18.360 170.350 18.680 170.670 ;
        RECT 24.640 170.380 24.960 170.700 ;
        RECT 25.200 170.380 25.520 170.700 ;
        RECT 27.600 170.940 27.920 171.260 ;
        RECT 28.160 170.940 28.480 171.260 ;
        RECT 34.440 171.230 34.760 171.550 ;
        RECT 35.000 171.230 35.320 171.550 ;
        RECT 43.000 171.230 43.320 171.550 ;
        RECT 43.560 171.230 43.880 171.550 ;
        RECT 59.640 173.870 59.960 174.190 ;
        RECT 60.200 173.870 60.520 174.190 ;
        RECT 68.200 173.870 68.520 174.190 ;
        RECT 68.760 173.870 69.080 174.190 ;
        RECT 49.840 170.940 50.160 171.260 ;
        RECT 50.400 170.940 50.720 171.260 ;
        RECT 27.600 170.380 27.920 170.700 ;
        RECT 28.160 170.380 28.480 170.700 ;
        RECT 34.440 170.350 34.760 170.670 ;
        RECT 35.000 170.350 35.320 170.670 ;
        RECT 43.000 170.350 43.320 170.670 ;
        RECT 43.560 170.350 43.880 170.670 ;
        RECT 49.840 170.380 50.160 170.700 ;
        RECT 50.400 170.380 50.720 170.700 ;
        RECT 52.800 170.940 53.120 171.260 ;
        RECT 53.360 170.940 53.680 171.260 ;
        RECT 59.640 171.230 59.960 171.550 ;
        RECT 60.200 171.230 60.520 171.550 ;
        RECT 68.200 171.230 68.520 171.550 ;
        RECT 68.760 171.230 69.080 171.550 ;
        RECT 84.840 173.870 85.160 174.190 ;
        RECT 85.400 173.870 85.720 174.190 ;
        RECT 93.400 173.870 93.720 174.190 ;
        RECT 93.960 173.870 94.280 174.190 ;
        RECT 75.040 170.940 75.360 171.260 ;
        RECT 75.600 170.940 75.920 171.260 ;
        RECT 52.800 170.380 53.120 170.700 ;
        RECT 53.360 170.380 53.680 170.700 ;
        RECT 59.640 170.350 59.960 170.670 ;
        RECT 60.200 170.350 60.520 170.670 ;
        RECT 68.200 170.350 68.520 170.670 ;
        RECT 68.760 170.350 69.080 170.670 ;
        RECT 75.040 170.380 75.360 170.700 ;
        RECT 75.600 170.380 75.920 170.700 ;
        RECT 78.000 170.940 78.320 171.260 ;
        RECT 78.560 170.940 78.880 171.260 ;
        RECT 84.840 171.230 85.160 171.550 ;
        RECT 85.400 171.230 85.720 171.550 ;
        RECT 93.400 171.230 93.720 171.550 ;
        RECT 93.960 171.230 94.280 171.550 ;
        RECT 110.040 173.870 110.360 174.190 ;
        RECT 110.600 173.870 110.920 174.190 ;
        RECT 122.560 173.870 122.880 174.190 ;
        RECT 123.120 173.870 123.440 174.190 ;
        RECT 100.240 170.940 100.560 171.260 ;
        RECT 100.800 170.940 101.120 171.260 ;
        RECT 78.000 170.380 78.320 170.700 ;
        RECT 78.560 170.380 78.880 170.700 ;
        RECT 84.840 170.350 85.160 170.670 ;
        RECT 85.400 170.350 85.720 170.670 ;
        RECT 93.400 170.350 93.720 170.670 ;
        RECT 93.960 170.350 94.280 170.670 ;
        RECT 100.240 170.380 100.560 170.700 ;
        RECT 100.800 170.380 101.120 170.700 ;
        RECT 103.200 170.940 103.520 171.260 ;
        RECT 103.760 170.940 104.080 171.260 ;
        RECT 118.600 172.990 118.920 173.310 ;
        RECT 119.160 172.990 119.480 173.310 ;
        RECT 118.600 172.110 118.920 172.430 ;
        RECT 119.160 172.110 119.480 172.430 ;
        RECT 122.560 172.110 122.880 172.430 ;
        RECT 123.120 172.110 123.440 172.430 ;
        RECT 143.740 171.940 144.060 172.260 ;
        RECT 144.300 171.940 144.620 172.260 ;
        RECT 147.700 171.940 148.020 172.260 ;
        RECT 148.260 171.940 148.580 172.260 ;
        RECT 110.040 171.230 110.360 171.550 ;
        RECT 110.600 171.230 110.920 171.550 ;
        RECT 103.200 170.380 103.520 170.700 ;
        RECT 103.760 170.380 104.080 170.700 ;
        RECT 110.040 170.350 110.360 170.670 ;
        RECT 110.600 170.350 110.920 170.670 ;
        RECT 19.265 168.830 19.585 169.150 ;
        RECT 15.720 168.110 16.040 168.430 ;
        RECT 16.280 168.110 16.600 168.430 ;
        RECT 19.265 168.270 19.585 168.590 ;
        RECT 17.800 167.710 18.120 168.030 ;
        RECT 18.360 167.710 18.680 168.030 ;
        RECT 33.535 168.830 33.855 169.150 ;
        RECT 33.535 168.270 33.855 168.590 ;
        RECT 44.465 168.830 44.785 169.150 ;
        RECT 36.520 168.110 36.840 168.430 ;
        RECT 37.080 168.110 37.400 168.430 ;
        RECT 40.920 168.110 41.240 168.430 ;
        RECT 41.480 168.110 41.800 168.430 ;
        RECT 44.465 168.270 44.785 168.590 ;
        RECT 34.440 167.710 34.760 168.030 ;
        RECT 35.000 167.710 35.320 168.030 ;
        RECT 43.000 167.710 43.320 168.030 ;
        RECT 43.560 167.710 43.880 168.030 ;
        RECT 58.735 168.830 59.055 169.150 ;
        RECT 58.735 168.270 59.055 168.590 ;
        RECT 69.665 168.830 69.985 169.150 ;
        RECT 61.720 168.110 62.040 168.430 ;
        RECT 62.280 168.110 62.600 168.430 ;
        RECT 66.120 168.110 66.440 168.430 ;
        RECT 66.680 168.110 67.000 168.430 ;
        RECT 69.665 168.270 69.985 168.590 ;
        RECT 59.640 167.710 59.960 168.030 ;
        RECT 60.200 167.710 60.520 168.030 ;
        RECT 68.200 167.710 68.520 168.030 ;
        RECT 68.760 167.710 69.080 168.030 ;
        RECT 83.935 168.830 84.255 169.150 ;
        RECT 83.935 168.270 84.255 168.590 ;
        RECT 94.865 168.830 95.185 169.150 ;
        RECT 86.920 168.110 87.240 168.430 ;
        RECT 87.480 168.110 87.800 168.430 ;
        RECT 91.320 168.110 91.640 168.430 ;
        RECT 91.880 168.110 92.200 168.430 ;
        RECT 94.865 168.270 95.185 168.590 ;
        RECT 84.840 167.710 85.160 168.030 ;
        RECT 85.400 167.710 85.720 168.030 ;
        RECT 93.400 167.710 93.720 168.030 ;
        RECT 93.960 167.710 94.280 168.030 ;
        RECT 109.135 168.830 109.455 169.150 ;
        RECT 109.135 168.270 109.455 168.590 ;
        RECT 112.120 168.110 112.440 168.430 ;
        RECT 112.680 168.110 113.000 168.430 ;
        RECT 110.040 167.710 110.360 168.030 ;
        RECT 110.600 167.710 110.920 168.030 ;
        RECT 17.800 166.830 18.120 167.150 ;
        RECT 18.360 166.830 18.680 167.150 ;
        RECT 17.800 164.190 18.120 164.510 ;
        RECT 18.360 164.190 18.680 164.510 ;
        RECT 34.440 166.830 34.760 167.150 ;
        RECT 35.000 166.830 35.320 167.150 ;
        RECT 43.000 166.830 43.320 167.150 ;
        RECT 43.560 166.830 43.880 167.150 ;
        RECT 24.640 163.900 24.960 164.220 ;
        RECT 25.200 163.900 25.520 164.220 ;
        RECT 17.800 163.310 18.120 163.630 ;
        RECT 18.360 163.310 18.680 163.630 ;
        RECT 24.640 163.340 24.960 163.660 ;
        RECT 25.200 163.340 25.520 163.660 ;
        RECT 27.600 163.900 27.920 164.220 ;
        RECT 28.160 163.900 28.480 164.220 ;
        RECT 34.440 164.190 34.760 164.510 ;
        RECT 35.000 164.190 35.320 164.510 ;
        RECT 43.000 164.190 43.320 164.510 ;
        RECT 43.560 164.190 43.880 164.510 ;
        RECT 59.640 166.830 59.960 167.150 ;
        RECT 60.200 166.830 60.520 167.150 ;
        RECT 68.200 166.830 68.520 167.150 ;
        RECT 68.760 166.830 69.080 167.150 ;
        RECT 49.840 163.900 50.160 164.220 ;
        RECT 50.400 163.900 50.720 164.220 ;
        RECT 27.600 163.340 27.920 163.660 ;
        RECT 28.160 163.340 28.480 163.660 ;
        RECT 34.440 163.310 34.760 163.630 ;
        RECT 35.000 163.310 35.320 163.630 ;
        RECT 43.000 163.310 43.320 163.630 ;
        RECT 43.560 163.310 43.880 163.630 ;
        RECT 49.840 163.340 50.160 163.660 ;
        RECT 50.400 163.340 50.720 163.660 ;
        RECT 52.800 163.900 53.120 164.220 ;
        RECT 53.360 163.900 53.680 164.220 ;
        RECT 59.640 164.190 59.960 164.510 ;
        RECT 60.200 164.190 60.520 164.510 ;
        RECT 68.200 164.190 68.520 164.510 ;
        RECT 68.760 164.190 69.080 164.510 ;
        RECT 84.840 166.830 85.160 167.150 ;
        RECT 85.400 166.830 85.720 167.150 ;
        RECT 93.400 166.830 93.720 167.150 ;
        RECT 93.960 166.830 94.280 167.150 ;
        RECT 75.040 163.900 75.360 164.220 ;
        RECT 75.600 163.900 75.920 164.220 ;
        RECT 52.800 163.340 53.120 163.660 ;
        RECT 53.360 163.340 53.680 163.660 ;
        RECT 59.640 163.310 59.960 163.630 ;
        RECT 60.200 163.310 60.520 163.630 ;
        RECT 68.200 163.310 68.520 163.630 ;
        RECT 68.760 163.310 69.080 163.630 ;
        RECT 75.040 163.340 75.360 163.660 ;
        RECT 75.600 163.340 75.920 163.660 ;
        RECT 78.000 163.900 78.320 164.220 ;
        RECT 78.560 163.900 78.880 164.220 ;
        RECT 84.840 164.190 85.160 164.510 ;
        RECT 85.400 164.190 85.720 164.510 ;
        RECT 93.400 164.190 93.720 164.510 ;
        RECT 93.960 164.190 94.280 164.510 ;
        RECT 110.040 166.830 110.360 167.150 ;
        RECT 110.600 166.830 110.920 167.150 ;
        RECT 100.240 163.900 100.560 164.220 ;
        RECT 100.800 163.900 101.120 164.220 ;
        RECT 78.000 163.340 78.320 163.660 ;
        RECT 78.560 163.340 78.880 163.660 ;
        RECT 84.840 163.310 85.160 163.630 ;
        RECT 85.400 163.310 85.720 163.630 ;
        RECT 93.400 163.310 93.720 163.630 ;
        RECT 93.960 163.310 94.280 163.630 ;
        RECT 100.240 163.340 100.560 163.660 ;
        RECT 100.800 163.340 101.120 163.660 ;
        RECT 103.200 163.900 103.520 164.220 ;
        RECT 103.760 163.900 104.080 164.220 ;
        RECT 110.040 164.190 110.360 164.510 ;
        RECT 110.600 164.190 110.920 164.510 ;
        RECT 103.200 163.340 103.520 163.660 ;
        RECT 103.760 163.340 104.080 163.660 ;
        RECT 110.040 163.310 110.360 163.630 ;
        RECT 110.600 163.310 110.920 163.630 ;
        RECT 17.800 160.670 18.120 160.990 ;
        RECT 18.360 160.670 18.680 160.990 ;
        RECT 34.440 160.670 34.760 160.990 ;
        RECT 35.000 160.670 35.320 160.990 ;
        RECT 43.000 160.670 43.320 160.990 ;
        RECT 43.560 160.670 43.880 160.990 ;
        RECT 59.640 160.670 59.960 160.990 ;
        RECT 60.200 160.670 60.520 160.990 ;
        RECT 68.200 160.670 68.520 160.990 ;
        RECT 68.760 160.670 69.080 160.990 ;
        RECT 84.840 160.670 85.160 160.990 ;
        RECT 85.400 160.670 85.720 160.990 ;
        RECT 93.400 160.670 93.720 160.990 ;
        RECT 93.960 160.670 94.280 160.990 ;
        RECT 110.040 160.670 110.360 160.990 ;
        RECT 110.600 160.670 110.920 160.990 ;
        RECT 143.740 170.180 144.060 170.500 ;
        RECT 144.300 170.180 144.620 170.500 ;
        RECT 147.700 170.180 148.020 170.500 ;
        RECT 148.260 170.180 148.580 170.500 ;
        RECT 118.600 169.470 118.920 169.790 ;
        RECT 119.160 169.470 119.480 169.790 ;
        RECT 122.560 169.470 122.880 169.790 ;
        RECT 123.120 169.470 123.440 169.790 ;
        RECT 118.600 168.590 118.920 168.910 ;
        RECT 119.160 168.590 119.480 168.910 ;
        RECT 122.560 168.590 122.880 168.910 ;
        RECT 123.120 168.590 123.440 168.910 ;
        RECT 17.800 155.390 18.120 155.710 ;
        RECT 18.360 155.390 18.680 155.710 ;
        RECT 21.760 155.390 22.080 155.710 ;
        RECT 22.320 155.390 22.640 155.710 ;
        RECT 30.480 155.390 30.800 155.710 ;
        RECT 31.040 155.390 31.360 155.710 ;
        RECT 34.440 155.390 34.760 155.710 ;
        RECT 35.000 155.390 35.320 155.710 ;
        RECT 43.000 155.390 43.320 155.710 ;
        RECT 43.560 155.390 43.880 155.710 ;
        RECT 46.960 155.390 47.280 155.710 ;
        RECT 47.520 155.390 47.840 155.710 ;
        RECT 55.680 155.390 56.000 155.710 ;
        RECT 56.240 155.390 56.560 155.710 ;
        RECT 59.640 155.390 59.960 155.710 ;
        RECT 60.200 155.390 60.520 155.710 ;
        RECT 68.200 155.390 68.520 155.710 ;
        RECT 68.760 155.390 69.080 155.710 ;
        RECT 72.160 155.390 72.480 155.710 ;
        RECT 72.720 155.390 73.040 155.710 ;
        RECT 80.880 155.390 81.200 155.710 ;
        RECT 81.440 155.390 81.760 155.710 ;
        RECT 84.840 155.390 85.160 155.710 ;
        RECT 85.400 155.390 85.720 155.710 ;
        RECT 93.400 155.390 93.720 155.710 ;
        RECT 93.960 155.390 94.280 155.710 ;
        RECT 97.360 155.390 97.680 155.710 ;
        RECT 97.920 155.390 98.240 155.710 ;
        RECT 106.080 155.390 106.400 155.710 ;
        RECT 106.640 155.390 106.960 155.710 ;
        RECT 110.040 155.390 110.360 155.710 ;
        RECT 110.600 155.390 110.920 155.710 ;
        RECT 118.600 165.950 118.920 166.270 ;
        RECT 119.160 165.950 119.480 166.270 ;
        RECT 122.560 165.950 122.880 166.270 ;
        RECT 123.120 165.950 123.440 166.270 ;
        RECT 122.560 165.070 122.880 165.390 ;
        RECT 123.120 165.070 123.440 165.390 ;
        RECT 147.700 166.660 148.020 166.980 ;
        RECT 148.260 166.660 148.580 166.980 ;
        RECT 147.700 165.780 148.020 166.100 ;
        RECT 148.260 165.780 148.580 166.100 ;
        RECT 143.740 164.900 144.060 165.220 ;
        RECT 144.300 164.900 144.620 165.220 ;
        RECT 122.560 162.430 122.880 162.750 ;
        RECT 123.120 162.430 123.440 162.750 ;
        RECT 122.560 161.550 122.880 161.870 ;
        RECT 123.120 161.550 123.440 161.870 ;
        RECT 143.740 161.380 144.060 161.700 ;
        RECT 144.300 161.380 144.620 161.700 ;
        RECT 147.700 161.380 148.020 161.700 ;
        RECT 148.260 161.380 148.580 161.700 ;
        RECT 143.740 159.620 144.060 159.940 ;
        RECT 144.300 159.620 144.620 159.940 ;
        RECT 147.700 159.620 148.020 159.940 ;
        RECT 148.260 159.620 148.580 159.940 ;
        RECT 122.560 158.910 122.880 159.230 ;
        RECT 123.120 158.910 123.440 159.230 ;
        RECT 122.560 158.030 122.880 158.350 ;
        RECT 123.120 158.030 123.440 158.350 ;
        RECT 124.720 157.590 125.040 157.910 ;
        RECT 125.280 157.590 125.600 157.910 ;
        RECT 143.740 156.100 144.060 156.420 ;
        RECT 144.300 156.100 144.620 156.420 ;
        RECT 147.700 156.100 148.020 156.420 ;
        RECT 148.260 156.100 148.580 156.420 ;
        RECT 122.560 155.390 122.880 155.710 ;
        RECT 123.120 155.390 123.440 155.710 ;
        RECT 122.560 154.510 122.880 154.830 ;
        RECT 123.120 154.510 123.440 154.830 ;
        RECT 118.600 153.630 118.920 153.950 ;
        RECT 119.160 153.630 119.480 153.950 ;
        RECT 143.740 152.580 144.060 152.900 ;
        RECT 144.300 152.580 144.620 152.900 ;
        RECT 147.700 152.580 148.020 152.900 ;
        RECT 148.260 152.580 148.580 152.900 ;
        RECT 116.440 150.550 116.760 150.870 ;
        RECT 117.000 150.550 117.320 150.870 ;
        RECT 143.740 150.820 144.060 151.140 ;
        RECT 144.300 150.820 144.620 151.140 ;
        RECT 147.700 150.820 148.020 151.140 ;
        RECT 148.260 150.820 148.580 151.140 ;
        RECT 17.800 150.110 18.120 150.430 ;
        RECT 18.360 150.110 18.680 150.430 ;
        RECT 21.760 150.110 22.080 150.430 ;
        RECT 22.320 150.110 22.640 150.430 ;
        RECT 30.480 150.110 30.800 150.430 ;
        RECT 31.040 150.110 31.360 150.430 ;
        RECT 34.440 150.110 34.760 150.430 ;
        RECT 35.000 150.110 35.320 150.430 ;
        RECT 43.000 150.110 43.320 150.430 ;
        RECT 43.560 150.110 43.880 150.430 ;
        RECT 46.960 150.110 47.280 150.430 ;
        RECT 47.520 150.110 47.840 150.430 ;
        RECT 55.680 150.110 56.000 150.430 ;
        RECT 56.240 150.110 56.560 150.430 ;
        RECT 59.640 150.110 59.960 150.430 ;
        RECT 60.200 150.110 60.520 150.430 ;
        RECT 68.200 150.110 68.520 150.430 ;
        RECT 68.760 150.110 69.080 150.430 ;
        RECT 72.160 150.110 72.480 150.430 ;
        RECT 72.720 150.110 73.040 150.430 ;
        RECT 80.880 150.110 81.200 150.430 ;
        RECT 81.440 150.110 81.760 150.430 ;
        RECT 84.840 150.110 85.160 150.430 ;
        RECT 85.400 150.110 85.720 150.430 ;
        RECT 93.400 150.110 93.720 150.430 ;
        RECT 93.960 150.110 94.280 150.430 ;
        RECT 97.360 150.110 97.680 150.430 ;
        RECT 97.920 150.110 98.240 150.430 ;
        RECT 106.080 150.110 106.400 150.430 ;
        RECT 106.640 150.110 106.960 150.430 ;
        RECT 110.040 150.110 110.360 150.430 ;
        RECT 110.600 150.110 110.920 150.430 ;
        RECT 147.700 149.940 148.020 150.260 ;
        RECT 148.260 149.940 148.580 150.260 ;
        RECT 17.800 148.350 18.120 148.670 ;
        RECT 18.360 148.350 18.680 148.670 ;
        RECT 21.760 148.350 22.080 148.670 ;
        RECT 22.320 148.350 22.640 148.670 ;
        RECT 30.480 148.350 30.800 148.670 ;
        RECT 31.040 148.350 31.360 148.670 ;
        RECT 34.440 148.350 34.760 148.670 ;
        RECT 35.000 148.350 35.320 148.670 ;
        RECT 43.000 148.350 43.320 148.670 ;
        RECT 43.560 148.350 43.880 148.670 ;
        RECT 46.960 148.350 47.280 148.670 ;
        RECT 47.520 148.350 47.840 148.670 ;
        RECT 55.680 148.350 56.000 148.670 ;
        RECT 56.240 148.350 56.560 148.670 ;
        RECT 59.640 148.350 59.960 148.670 ;
        RECT 60.200 148.350 60.520 148.670 ;
        RECT 68.200 148.350 68.520 148.670 ;
        RECT 68.760 148.350 69.080 148.670 ;
        RECT 72.160 148.350 72.480 148.670 ;
        RECT 72.720 148.350 73.040 148.670 ;
        RECT 80.880 148.350 81.200 148.670 ;
        RECT 81.440 148.350 81.760 148.670 ;
        RECT 84.840 148.350 85.160 148.670 ;
        RECT 85.400 148.350 85.720 148.670 ;
        RECT 93.400 148.350 93.720 148.670 ;
        RECT 93.960 148.350 94.280 148.670 ;
        RECT 97.360 148.350 97.680 148.670 ;
        RECT 97.920 148.350 98.240 148.670 ;
        RECT 106.080 148.350 106.400 148.670 ;
        RECT 106.640 148.350 106.960 148.670 ;
        RECT 110.040 148.350 110.360 148.670 ;
        RECT 110.600 148.350 110.920 148.670 ;
        RECT 21.760 147.470 22.080 147.790 ;
        RECT 22.320 147.470 22.640 147.790 ;
        RECT 30.480 147.470 30.800 147.790 ;
        RECT 31.040 147.470 31.360 147.790 ;
        RECT 46.960 147.470 47.280 147.790 ;
        RECT 47.520 147.470 47.840 147.790 ;
        RECT 55.680 147.470 56.000 147.790 ;
        RECT 56.240 147.470 56.560 147.790 ;
        RECT 72.160 147.470 72.480 147.790 ;
        RECT 72.720 147.470 73.040 147.790 ;
        RECT 80.880 147.470 81.200 147.790 ;
        RECT 81.440 147.470 81.760 147.790 ;
        RECT 97.360 147.470 97.680 147.790 ;
        RECT 97.920 147.470 98.240 147.790 ;
        RECT 106.080 147.470 106.400 147.790 ;
        RECT 106.640 147.470 106.960 147.790 ;
        RECT 143.740 147.300 144.060 147.620 ;
        RECT 144.300 147.300 144.620 147.620 ;
        RECT 147.700 147.300 148.020 147.620 ;
        RECT 148.260 147.300 148.580 147.620 ;
        RECT 17.800 146.590 18.120 146.910 ;
        RECT 18.360 146.590 18.680 146.910 ;
        RECT 34.440 146.590 34.760 146.910 ;
        RECT 35.000 146.590 35.320 146.910 ;
        RECT 43.000 146.590 43.320 146.910 ;
        RECT 43.560 146.590 43.880 146.910 ;
        RECT 59.640 146.590 59.960 146.910 ;
        RECT 60.200 146.590 60.520 146.910 ;
        RECT 68.200 146.590 68.520 146.910 ;
        RECT 68.760 146.590 69.080 146.910 ;
        RECT 84.840 146.590 85.160 146.910 ;
        RECT 85.400 146.590 85.720 146.910 ;
        RECT 93.400 146.590 93.720 146.910 ;
        RECT 93.960 146.590 94.280 146.910 ;
        RECT 110.040 146.590 110.360 146.910 ;
        RECT 110.600 146.590 110.920 146.910 ;
        RECT 17.800 145.710 18.120 146.030 ;
        RECT 18.360 145.710 18.680 146.030 ;
        RECT 34.440 145.710 34.760 146.030 ;
        RECT 35.000 145.710 35.320 146.030 ;
        RECT 43.000 145.710 43.320 146.030 ;
        RECT 43.560 145.710 43.880 146.030 ;
        RECT 59.640 145.710 59.960 146.030 ;
        RECT 60.200 145.710 60.520 146.030 ;
        RECT 68.200 145.710 68.520 146.030 ;
        RECT 68.760 145.710 69.080 146.030 ;
        RECT 84.840 145.710 85.160 146.030 ;
        RECT 85.400 145.710 85.720 146.030 ;
        RECT 93.400 145.710 93.720 146.030 ;
        RECT 93.960 145.710 94.280 146.030 ;
        RECT 110.040 145.710 110.360 146.030 ;
        RECT 110.600 145.710 110.920 146.030 ;
        RECT 143.740 145.540 144.060 145.860 ;
        RECT 144.300 145.540 144.620 145.860 ;
        RECT 147.700 145.540 148.020 145.860 ;
        RECT 148.260 145.540 148.580 145.860 ;
        RECT 17.800 143.070 18.120 143.390 ;
        RECT 18.360 143.070 18.680 143.390 ;
        RECT 34.440 143.070 34.760 143.390 ;
        RECT 35.000 143.070 35.320 143.390 ;
        RECT 21.760 142.190 22.080 142.510 ;
        RECT 22.320 142.190 22.640 142.510 ;
        RECT 30.480 142.190 30.800 142.510 ;
        RECT 31.040 142.190 31.360 142.510 ;
        RECT 43.000 143.070 43.320 143.390 ;
        RECT 43.560 143.070 43.880 143.390 ;
        RECT 59.640 143.070 59.960 143.390 ;
        RECT 60.200 143.070 60.520 143.390 ;
        RECT 46.960 142.190 47.280 142.510 ;
        RECT 47.520 142.190 47.840 142.510 ;
        RECT 55.680 142.190 56.000 142.510 ;
        RECT 56.240 142.190 56.560 142.510 ;
        RECT 68.200 143.070 68.520 143.390 ;
        RECT 68.760 143.070 69.080 143.390 ;
        RECT 84.840 143.070 85.160 143.390 ;
        RECT 85.400 143.070 85.720 143.390 ;
        RECT 72.160 142.190 72.480 142.510 ;
        RECT 72.720 142.190 73.040 142.510 ;
        RECT 80.880 142.190 81.200 142.510 ;
        RECT 81.440 142.190 81.760 142.510 ;
        RECT 93.400 143.070 93.720 143.390 ;
        RECT 93.960 143.070 94.280 143.390 ;
        RECT 110.040 143.070 110.360 143.390 ;
        RECT 110.600 143.070 110.920 143.390 ;
        RECT 97.360 142.190 97.680 142.510 ;
        RECT 97.920 142.190 98.240 142.510 ;
        RECT 106.080 142.190 106.400 142.510 ;
        RECT 106.640 142.190 106.960 142.510 ;
        RECT 122.560 142.190 122.880 142.510 ;
        RECT 123.120 142.190 123.440 142.510 ;
        RECT 118.600 141.310 118.920 141.630 ;
        RECT 119.160 141.310 119.480 141.630 ;
        RECT 17.800 140.430 18.120 140.750 ;
        RECT 18.360 140.430 18.680 140.750 ;
        RECT 21.760 140.430 22.080 140.750 ;
        RECT 22.320 140.430 22.640 140.750 ;
        RECT 30.480 140.430 30.800 140.750 ;
        RECT 31.040 140.430 31.360 140.750 ;
        RECT 34.440 140.430 34.760 140.750 ;
        RECT 35.000 140.430 35.320 140.750 ;
        RECT 43.000 140.430 43.320 140.750 ;
        RECT 43.560 140.430 43.880 140.750 ;
        RECT 46.960 140.430 47.280 140.750 ;
        RECT 47.520 140.430 47.840 140.750 ;
        RECT 55.680 140.430 56.000 140.750 ;
        RECT 56.240 140.430 56.560 140.750 ;
        RECT 59.640 140.430 59.960 140.750 ;
        RECT 60.200 140.430 60.520 140.750 ;
        RECT 68.200 140.430 68.520 140.750 ;
        RECT 68.760 140.430 69.080 140.750 ;
        RECT 72.160 140.430 72.480 140.750 ;
        RECT 72.720 140.430 73.040 140.750 ;
        RECT 80.880 140.430 81.200 140.750 ;
        RECT 81.440 140.430 81.760 140.750 ;
        RECT 84.840 140.430 85.160 140.750 ;
        RECT 85.400 140.430 85.720 140.750 ;
        RECT 93.400 140.430 93.720 140.750 ;
        RECT 93.960 140.430 94.280 140.750 ;
        RECT 97.360 140.430 97.680 140.750 ;
        RECT 97.920 140.430 98.240 140.750 ;
        RECT 106.080 140.430 106.400 140.750 ;
        RECT 106.640 140.430 106.960 140.750 ;
        RECT 110.040 140.430 110.360 140.750 ;
        RECT 110.600 140.430 110.920 140.750 ;
        RECT 118.600 140.430 118.920 140.750 ;
        RECT 119.160 140.430 119.480 140.750 ;
        RECT 122.560 140.430 122.880 140.750 ;
        RECT 123.120 140.430 123.440 140.750 ;
        RECT 17.800 139.550 18.120 139.870 ;
        RECT 18.360 139.550 18.680 139.870 ;
        RECT 21.760 139.550 22.080 139.870 ;
        RECT 22.320 139.550 22.640 139.870 ;
        RECT 30.480 139.550 30.800 139.870 ;
        RECT 31.040 139.550 31.360 139.870 ;
        RECT 34.440 139.550 34.760 139.870 ;
        RECT 35.000 139.550 35.320 139.870 ;
        RECT 43.000 139.550 43.320 139.870 ;
        RECT 43.560 139.550 43.880 139.870 ;
        RECT 46.960 139.550 47.280 139.870 ;
        RECT 47.520 139.550 47.840 139.870 ;
        RECT 55.680 139.550 56.000 139.870 ;
        RECT 56.240 139.550 56.560 139.870 ;
        RECT 59.640 139.550 59.960 139.870 ;
        RECT 60.200 139.550 60.520 139.870 ;
        RECT 68.200 139.550 68.520 139.870 ;
        RECT 68.760 139.550 69.080 139.870 ;
        RECT 72.160 139.550 72.480 139.870 ;
        RECT 72.720 139.550 73.040 139.870 ;
        RECT 80.880 139.550 81.200 139.870 ;
        RECT 81.440 139.550 81.760 139.870 ;
        RECT 84.840 139.550 85.160 139.870 ;
        RECT 85.400 139.550 85.720 139.870 ;
        RECT 93.400 139.550 93.720 139.870 ;
        RECT 93.960 139.550 94.280 139.870 ;
        RECT 97.360 139.550 97.680 139.870 ;
        RECT 97.920 139.550 98.240 139.870 ;
        RECT 106.080 139.550 106.400 139.870 ;
        RECT 106.640 139.550 106.960 139.870 ;
        RECT 110.040 139.550 110.360 139.870 ;
        RECT 110.600 139.550 110.920 139.870 ;
        RECT 118.600 139.550 118.920 139.870 ;
        RECT 119.160 139.550 119.480 139.870 ;
        RECT 122.560 139.550 122.880 139.870 ;
        RECT 123.120 139.550 123.440 139.870 ;
        RECT 147.700 142.020 148.020 142.340 ;
        RECT 148.260 142.020 148.580 142.340 ;
        RECT 147.700 141.140 148.020 141.460 ;
        RECT 148.260 141.140 148.580 141.460 ;
        RECT 143.740 140.260 144.060 140.580 ;
        RECT 144.300 140.260 144.620 140.580 ;
        RECT 143.740 136.740 144.060 137.060 ;
        RECT 144.300 136.740 144.620 137.060 ;
        RECT 147.700 136.740 148.020 137.060 ;
        RECT 148.260 136.740 148.580 137.060 ;
        RECT 96.540 135.660 96.860 135.980 ;
        RECT 96.540 135.100 96.860 135.420 ;
        RECT 82.260 134.690 82.580 135.010 ;
        RECT 143.740 134.980 144.060 135.300 ;
        RECT 144.300 134.980 144.620 135.300 ;
        RECT 147.700 134.980 148.020 135.300 ;
        RECT 148.260 134.980 148.580 135.300 ;
        RECT 82.260 134.130 82.580 134.450 ;
        RECT 71.340 133.720 71.660 134.040 ;
        RECT 71.340 133.160 71.660 133.480 ;
        RECT 57.060 132.750 57.380 133.070 ;
        RECT 57.060 132.190 57.380 132.510 ;
        RECT 46.140 131.780 46.460 132.100 ;
        RECT 46.140 131.220 46.460 131.540 ;
        RECT 143.740 131.460 144.060 131.780 ;
        RECT 144.300 131.460 144.620 131.780 ;
        RECT 147.700 131.460 148.020 131.780 ;
        RECT 148.260 131.460 148.580 131.780 ;
        RECT 31.860 130.810 32.180 131.130 ;
        RECT 31.860 130.250 32.180 130.570 ;
        RECT 20.940 129.840 21.260 130.160 ;
        RECT 20.940 129.280 21.260 129.600 ;
        RECT 45.265 128.870 45.585 129.190 ;
        RECT 45.265 128.310 45.585 128.630 ;
        RECT 32.730 127.900 33.050 128.220 ;
        RECT 143.740 127.940 144.060 128.260 ;
        RECT 144.300 127.940 144.620 128.260 ;
        RECT 147.700 127.940 148.020 128.260 ;
        RECT 148.260 127.940 148.580 128.260 ;
        RECT 32.730 127.340 33.050 127.660 ;
        RECT 20.065 126.930 20.385 127.250 ;
        RECT 20.065 126.370 20.385 126.690 ;
        RECT 94.865 125.960 95.185 126.280 ;
        RECT 143.740 126.180 144.060 126.500 ;
        RECT 144.300 126.180 144.620 126.500 ;
        RECT 147.700 126.180 148.020 126.500 ;
        RECT 148.260 126.180 148.580 126.500 ;
        RECT 94.865 125.400 95.185 125.720 ;
        RECT 83.930 124.990 84.250 125.310 ;
        RECT 147.700 125.300 148.020 125.620 ;
        RECT 148.260 125.300 148.580 125.620 ;
        RECT 83.930 124.430 84.250 124.750 ;
        RECT 69.665 124.020 69.985 124.340 ;
        RECT 58.730 123.050 59.050 123.370 ;
        RECT 69.665 123.460 69.985 123.780 ;
        RECT 58.730 122.490 59.050 122.810 ;
        RECT 44.465 122.080 44.785 122.400 ;
        RECT 143.740 122.660 144.060 122.980 ;
        RECT 144.300 122.660 144.620 122.980 ;
        RECT 147.700 122.660 148.020 122.980 ;
        RECT 148.260 122.660 148.580 122.980 ;
        RECT 44.465 121.520 44.785 121.840 ;
        RECT 33.530 121.110 33.850 121.430 ;
        RECT 143.740 120.900 144.060 121.220 ;
        RECT 144.300 120.900 144.620 121.220 ;
        RECT 147.700 120.900 148.020 121.220 ;
        RECT 148.260 120.900 148.580 121.220 ;
        RECT 33.530 120.550 33.850 120.870 ;
        RECT 19.265 120.140 19.585 120.460 ;
        RECT 19.265 119.580 19.585 119.900 ;
        RECT 40.890 119.170 41.210 119.490 ;
        RECT 40.890 118.610 41.210 118.930 ;
        RECT 36.490 118.200 36.810 118.520 ;
        RECT 36.490 117.640 36.810 117.960 ;
        RECT 15.690 117.230 16.010 117.550 ;
        RECT 116.410 117.500 116.730 117.820 ;
        RECT 15.690 116.670 16.010 116.990 ;
        RECT 116.410 116.940 116.730 117.260 ;
        RECT 117.810 117.500 118.130 117.820 ;
        RECT 117.810 116.940 118.130 117.260 ;
        RECT 57.800 115.010 58.120 115.330 ;
        RECT 58.360 115.010 58.680 115.330 ;
        RECT 116.440 115.010 116.760 115.330 ;
        RECT 117.000 115.010 117.320 115.330 ;
        RECT 147.700 117.380 148.020 117.700 ;
        RECT 148.260 117.380 148.580 117.700 ;
        RECT 147.700 116.500 148.020 116.820 ;
        RECT 148.260 116.500 148.580 116.820 ;
        RECT 143.740 115.620 144.060 115.940 ;
        RECT 144.300 115.620 144.620 115.940 ;
        RECT 57.770 111.130 58.090 111.450 ;
        RECT 57.770 110.570 58.090 110.890 ;
        RECT 83.060 113.070 83.380 113.390 ;
        RECT 83.620 113.070 83.940 113.390 ;
        RECT 117.840 113.070 118.160 113.390 ;
        RECT 118.400 113.070 118.720 113.390 ;
        RECT 143.740 112.100 144.060 112.420 ;
        RECT 144.300 112.100 144.620 112.420 ;
        RECT 147.700 112.100 148.020 112.420 ;
        RECT 148.260 112.100 148.580 112.420 ;
        RECT 83.030 111.130 83.350 111.450 ;
        RECT 83.030 110.570 83.350 110.890 ;
        RECT 23.470 109.430 23.790 109.750 ;
        RECT 23.470 108.870 23.790 109.190 ;
        RECT 117.330 109.430 117.650 109.750 ;
        RECT 117.330 108.870 117.650 109.190 ;
        RECT 22.070 106.370 22.390 106.690 ;
        RECT 22.070 105.810 22.390 106.130 ;
        RECT 26.270 106.370 26.590 106.690 ;
        RECT 26.270 105.810 26.590 106.130 ;
        RECT 44.470 106.370 44.790 106.690 ;
        RECT 44.470 105.810 44.790 106.130 ;
        RECT 48.670 106.370 48.990 106.690 ;
        RECT 48.670 105.810 48.990 106.130 ;
        RECT 92.130 106.370 92.450 106.690 ;
        RECT 92.130 105.810 92.450 106.130 ;
        RECT 96.330 106.370 96.650 106.690 ;
        RECT 96.330 105.810 96.650 106.130 ;
        RECT 114.530 106.370 114.850 106.690 ;
        RECT 114.530 105.810 114.850 106.130 ;
        RECT 118.730 106.370 119.050 106.690 ;
        RECT 118.730 105.810 119.050 106.130 ;
        RECT 19.270 103.310 19.590 103.630 ;
        RECT 19.270 102.750 19.590 103.070 ;
        RECT 20.670 103.310 20.990 103.630 ;
        RECT 20.670 102.750 20.990 103.070 ;
        RECT 27.670 103.310 27.990 103.630 ;
        RECT 27.670 102.750 27.990 103.070 ;
        RECT 29.070 103.310 29.390 103.630 ;
        RECT 29.070 102.750 29.390 103.070 ;
        RECT 41.670 103.310 41.990 103.630 ;
        RECT 41.670 102.750 41.990 103.070 ;
        RECT 43.070 103.310 43.390 103.630 ;
        RECT 43.070 102.750 43.390 103.070 ;
        RECT 50.070 103.310 50.390 103.630 ;
        RECT 50.070 102.750 50.390 103.070 ;
        RECT 51.470 103.310 51.790 103.630 ;
        RECT 51.470 102.750 51.790 103.070 ;
        RECT 89.330 103.310 89.650 103.630 ;
        RECT 89.330 102.750 89.650 103.070 ;
        RECT 90.730 103.310 91.050 103.630 ;
        RECT 90.730 102.750 91.050 103.070 ;
        RECT 97.730 103.310 98.050 103.630 ;
        RECT 97.730 102.750 98.050 103.070 ;
        RECT 99.130 103.310 99.450 103.630 ;
        RECT 99.130 102.750 99.450 103.070 ;
        RECT 111.730 103.310 112.050 103.630 ;
        RECT 111.730 102.750 112.050 103.070 ;
        RECT 113.130 103.310 113.450 103.630 ;
        RECT 113.130 102.750 113.450 103.070 ;
        RECT 120.130 103.310 120.450 103.630 ;
        RECT 120.130 102.750 120.450 103.070 ;
        RECT 121.530 103.310 121.850 103.630 ;
        RECT 121.530 102.750 121.850 103.070 ;
        RECT 12.270 101.280 12.590 101.600 ;
        RECT 12.270 100.720 12.590 101.040 ;
        RECT 143.740 110.340 144.060 110.660 ;
        RECT 144.300 110.340 144.620 110.660 ;
        RECT 147.700 110.340 148.020 110.660 ;
        RECT 148.260 110.340 148.580 110.660 ;
        RECT 143.740 106.820 144.060 107.140 ;
        RECT 144.300 106.820 144.620 107.140 ;
        RECT 147.700 106.820 148.020 107.140 ;
        RECT 148.260 106.820 148.580 107.140 ;
        RECT 143.740 103.300 144.060 103.620 ;
        RECT 144.300 103.300 144.620 103.620 ;
        RECT 147.700 103.300 148.020 103.620 ;
        RECT 148.260 103.300 148.580 103.620 ;
        RECT 128.530 101.280 128.850 101.600 ;
        RECT 143.740 101.540 144.060 101.860 ;
        RECT 144.300 101.540 144.620 101.860 ;
        RECT 147.700 101.540 148.020 101.860 ;
        RECT 148.260 101.540 148.580 101.860 ;
        RECT 128.530 100.720 128.850 101.040 ;
        RECT 24.870 100.250 25.190 100.570 ;
        RECT 24.870 99.690 25.190 100.010 ;
        RECT 45.870 100.250 46.190 100.570 ;
        RECT 45.870 99.690 46.190 100.010 ;
        RECT 94.930 100.250 95.250 100.570 ;
        RECT 94.930 99.690 95.250 100.010 ;
        RECT 115.930 100.250 116.250 100.570 ;
        RECT 115.930 99.690 116.250 100.010 ;
        RECT 13.670 97.190 13.990 97.510 ;
        RECT 13.670 96.630 13.990 96.950 ;
        RECT 15.070 97.190 15.390 97.510 ;
        RECT 15.070 96.630 15.390 96.950 ;
        RECT 16.470 97.190 16.790 97.510 ;
        RECT 16.470 96.630 16.790 96.950 ;
        RECT 17.870 97.190 18.190 97.510 ;
        RECT 17.870 96.630 18.190 96.950 ;
        RECT 30.470 97.190 30.790 97.510 ;
        RECT 30.470 96.630 30.790 96.950 ;
        RECT 31.870 97.190 32.190 97.510 ;
        RECT 31.870 96.630 32.190 96.950 ;
        RECT 33.270 97.190 33.590 97.510 ;
        RECT 33.270 96.630 33.590 96.950 ;
        RECT 34.670 97.190 34.990 97.510 ;
        RECT 34.670 96.630 34.990 96.950 ;
        RECT 36.070 97.190 36.390 97.510 ;
        RECT 36.070 96.630 36.390 96.950 ;
        RECT 37.470 97.190 37.790 97.510 ;
        RECT 37.470 96.630 37.790 96.950 ;
        RECT 38.870 97.190 39.190 97.510 ;
        RECT 38.870 96.630 39.190 96.950 ;
        RECT 40.270 97.190 40.590 97.510 ;
        RECT 40.270 96.630 40.590 96.950 ;
        RECT 52.870 97.190 53.190 97.510 ;
        RECT 52.870 96.630 53.190 96.950 ;
        RECT 54.270 97.190 54.590 97.510 ;
        RECT 54.270 96.630 54.590 96.950 ;
        RECT 55.670 97.190 55.990 97.510 ;
        RECT 55.670 96.630 55.990 96.950 ;
        RECT 57.070 97.190 57.390 97.510 ;
        RECT 57.070 96.630 57.390 96.950 ;
        RECT 83.730 97.190 84.050 97.510 ;
        RECT 83.730 96.630 84.050 96.950 ;
        RECT 85.130 97.190 85.450 97.510 ;
        RECT 85.130 96.630 85.450 96.950 ;
        RECT 86.530 97.190 86.850 97.510 ;
        RECT 86.530 96.630 86.850 96.950 ;
        RECT 87.930 97.190 88.250 97.510 ;
        RECT 87.930 96.630 88.250 96.950 ;
        RECT 100.530 97.190 100.850 97.510 ;
        RECT 100.530 96.630 100.850 96.950 ;
        RECT 101.930 97.190 102.250 97.510 ;
        RECT 101.930 96.630 102.250 96.950 ;
        RECT 103.330 97.190 103.650 97.510 ;
        RECT 103.330 96.630 103.650 96.950 ;
        RECT 104.730 97.190 105.050 97.510 ;
        RECT 104.730 96.630 105.050 96.950 ;
        RECT 106.130 97.190 106.450 97.510 ;
        RECT 106.130 96.630 106.450 96.950 ;
        RECT 107.530 97.190 107.850 97.510 ;
        RECT 107.530 96.630 107.850 96.950 ;
        RECT 108.930 97.190 109.250 97.510 ;
        RECT 108.930 96.630 109.250 96.950 ;
        RECT 110.330 97.190 110.650 97.510 ;
        RECT 110.330 96.630 110.650 96.950 ;
        RECT 122.930 97.190 123.250 97.510 ;
        RECT 122.930 96.630 123.250 96.950 ;
        RECT 124.330 97.190 124.650 97.510 ;
        RECT 124.330 96.630 124.650 96.950 ;
        RECT 125.730 97.190 126.050 97.510 ;
        RECT 125.730 96.630 126.050 96.950 ;
        RECT 127.130 97.190 127.450 97.510 ;
        RECT 127.130 96.630 127.450 96.950 ;
        RECT 47.270 94.130 47.590 94.450 ;
        RECT 47.270 93.570 47.590 93.890 ;
        RECT 93.530 94.130 93.850 94.450 ;
        RECT 93.530 93.570 93.850 93.890 ;
        RECT 23.470 92.030 23.790 92.350 ;
        RECT 23.470 91.470 23.790 91.790 ;
        RECT 117.330 92.030 117.650 92.350 ;
        RECT 117.330 91.470 117.650 91.790 ;
        RECT 22.070 88.970 22.390 89.290 ;
        RECT 22.070 88.410 22.390 88.730 ;
        RECT 26.270 88.970 26.590 89.290 ;
        RECT 26.270 88.410 26.590 88.730 ;
        RECT 44.470 88.970 44.790 89.290 ;
        RECT 44.470 88.410 44.790 88.730 ;
        RECT 48.670 88.970 48.990 89.290 ;
        RECT 48.670 88.410 48.990 88.730 ;
        RECT 92.130 88.970 92.450 89.290 ;
        RECT 92.130 88.410 92.450 88.730 ;
        RECT 96.330 88.970 96.650 89.290 ;
        RECT 96.330 88.410 96.650 88.730 ;
        RECT 114.530 88.970 114.850 89.290 ;
        RECT 114.530 88.410 114.850 88.730 ;
        RECT 118.730 88.970 119.050 89.290 ;
        RECT 118.730 88.410 119.050 88.730 ;
        RECT 19.270 85.910 19.590 86.230 ;
        RECT 19.270 85.350 19.590 85.670 ;
        RECT 20.670 85.910 20.990 86.230 ;
        RECT 20.670 85.350 20.990 85.670 ;
        RECT 27.670 85.910 27.990 86.230 ;
        RECT 27.670 85.350 27.990 85.670 ;
        RECT 29.070 85.910 29.390 86.230 ;
        RECT 29.070 85.350 29.390 85.670 ;
        RECT 41.670 85.910 41.990 86.230 ;
        RECT 41.670 85.350 41.990 85.670 ;
        RECT 43.070 85.910 43.390 86.230 ;
        RECT 43.070 85.350 43.390 85.670 ;
        RECT 50.070 85.910 50.390 86.230 ;
        RECT 50.070 85.350 50.390 85.670 ;
        RECT 51.470 85.910 51.790 86.230 ;
        RECT 51.470 85.350 51.790 85.670 ;
        RECT 89.330 85.910 89.650 86.230 ;
        RECT 89.330 85.350 89.650 85.670 ;
        RECT 90.730 85.910 91.050 86.230 ;
        RECT 90.730 85.350 91.050 85.670 ;
        RECT 97.730 85.910 98.050 86.230 ;
        RECT 97.730 85.350 98.050 85.670 ;
        RECT 99.130 85.910 99.450 86.230 ;
        RECT 99.130 85.350 99.450 85.670 ;
        RECT 111.730 85.910 112.050 86.230 ;
        RECT 111.730 85.350 112.050 85.670 ;
        RECT 113.130 85.910 113.450 86.230 ;
        RECT 113.130 85.350 113.450 85.670 ;
        RECT 120.130 85.910 120.450 86.230 ;
        RECT 120.130 85.350 120.450 85.670 ;
        RECT 121.530 85.910 121.850 86.230 ;
        RECT 121.530 85.350 121.850 85.670 ;
        RECT 12.270 83.880 12.590 84.200 ;
        RECT 12.270 83.320 12.590 83.640 ;
        RECT 147.700 100.660 148.020 100.980 ;
        RECT 148.260 100.660 148.580 100.980 ;
        RECT 143.740 98.020 144.060 98.340 ;
        RECT 144.300 98.020 144.620 98.340 ;
        RECT 147.700 98.020 148.020 98.340 ;
        RECT 148.260 98.020 148.580 98.340 ;
        RECT 143.740 96.260 144.060 96.580 ;
        RECT 144.300 96.260 144.620 96.580 ;
        RECT 147.700 96.260 148.020 96.580 ;
        RECT 148.260 96.260 148.580 96.580 ;
        RECT 147.700 92.740 148.020 93.060 ;
        RECT 148.260 92.740 148.580 93.060 ;
        RECT 147.700 91.860 148.020 92.180 ;
        RECT 148.260 91.860 148.580 92.180 ;
        RECT 143.740 90.980 144.060 91.300 ;
        RECT 144.300 90.980 144.620 91.300 ;
        RECT 143.740 87.460 144.060 87.780 ;
        RECT 144.300 87.460 144.620 87.780 ;
        RECT 147.700 87.460 148.020 87.780 ;
        RECT 148.260 87.460 148.580 87.780 ;
        RECT 143.740 85.700 144.060 86.020 ;
        RECT 144.300 85.700 144.620 86.020 ;
        RECT 147.700 85.700 148.020 86.020 ;
        RECT 148.260 85.700 148.580 86.020 ;
        RECT 128.530 83.880 128.850 84.200 ;
        RECT 128.530 83.320 128.850 83.640 ;
        RECT 24.870 82.850 25.190 83.170 ;
        RECT 24.870 82.290 25.190 82.610 ;
        RECT 45.870 82.850 46.190 83.170 ;
        RECT 45.870 82.290 46.190 82.610 ;
        RECT 94.930 82.850 95.250 83.170 ;
        RECT 94.930 82.290 95.250 82.610 ;
        RECT 115.930 82.850 116.250 83.170 ;
        RECT 115.930 82.290 116.250 82.610 ;
        RECT 13.670 79.790 13.990 80.110 ;
        RECT 13.670 79.230 13.990 79.550 ;
        RECT 15.070 79.790 15.390 80.110 ;
        RECT 15.070 79.230 15.390 79.550 ;
        RECT 16.470 79.790 16.790 80.110 ;
        RECT 16.470 79.230 16.790 79.550 ;
        RECT 17.870 79.790 18.190 80.110 ;
        RECT 17.870 79.230 18.190 79.550 ;
        RECT 30.470 79.790 30.790 80.110 ;
        RECT 30.470 79.230 30.790 79.550 ;
        RECT 31.870 79.790 32.190 80.110 ;
        RECT 31.870 79.230 32.190 79.550 ;
        RECT 33.270 79.790 33.590 80.110 ;
        RECT 33.270 79.230 33.590 79.550 ;
        RECT 34.670 79.790 34.990 80.110 ;
        RECT 34.670 79.230 34.990 79.550 ;
        RECT 36.070 79.790 36.390 80.110 ;
        RECT 36.070 79.230 36.390 79.550 ;
        RECT 37.470 79.790 37.790 80.110 ;
        RECT 37.470 79.230 37.790 79.550 ;
        RECT 38.870 79.790 39.190 80.110 ;
        RECT 38.870 79.230 39.190 79.550 ;
        RECT 40.270 79.790 40.590 80.110 ;
        RECT 40.270 79.230 40.590 79.550 ;
        RECT 52.870 79.790 53.190 80.110 ;
        RECT 52.870 79.230 53.190 79.550 ;
        RECT 54.270 79.790 54.590 80.110 ;
        RECT 54.270 79.230 54.590 79.550 ;
        RECT 55.670 79.790 55.990 80.110 ;
        RECT 55.670 79.230 55.990 79.550 ;
        RECT 57.070 79.790 57.390 80.110 ;
        RECT 57.070 79.230 57.390 79.550 ;
        RECT 83.730 79.790 84.050 80.110 ;
        RECT 83.730 79.230 84.050 79.550 ;
        RECT 85.130 79.790 85.450 80.110 ;
        RECT 85.130 79.230 85.450 79.550 ;
        RECT 86.530 79.790 86.850 80.110 ;
        RECT 86.530 79.230 86.850 79.550 ;
        RECT 87.930 79.790 88.250 80.110 ;
        RECT 87.930 79.230 88.250 79.550 ;
        RECT 100.530 79.790 100.850 80.110 ;
        RECT 100.530 79.230 100.850 79.550 ;
        RECT 101.930 79.790 102.250 80.110 ;
        RECT 101.930 79.230 102.250 79.550 ;
        RECT 103.330 79.790 103.650 80.110 ;
        RECT 103.330 79.230 103.650 79.550 ;
        RECT 104.730 79.790 105.050 80.110 ;
        RECT 104.730 79.230 105.050 79.550 ;
        RECT 106.130 79.790 106.450 80.110 ;
        RECT 106.130 79.230 106.450 79.550 ;
        RECT 107.530 79.790 107.850 80.110 ;
        RECT 107.530 79.230 107.850 79.550 ;
        RECT 108.930 79.790 109.250 80.110 ;
        RECT 108.930 79.230 109.250 79.550 ;
        RECT 110.330 79.790 110.650 80.110 ;
        RECT 110.330 79.230 110.650 79.550 ;
        RECT 122.930 79.790 123.250 80.110 ;
        RECT 122.930 79.230 123.250 79.550 ;
        RECT 124.330 79.790 124.650 80.110 ;
        RECT 124.330 79.230 124.650 79.550 ;
        RECT 125.730 79.790 126.050 80.110 ;
        RECT 125.730 79.230 126.050 79.550 ;
        RECT 127.130 79.790 127.450 80.110 ;
        RECT 127.130 79.230 127.450 79.550 ;
        RECT 47.270 76.730 47.590 77.050 ;
        RECT 47.270 76.170 47.590 76.490 ;
        RECT 93.530 76.730 93.850 77.050 ;
        RECT 93.530 76.170 93.850 76.490 ;
        RECT 23.470 74.630 23.790 74.950 ;
        RECT 23.470 74.070 23.790 74.390 ;
        RECT 117.330 74.630 117.650 74.950 ;
        RECT 117.330 74.070 117.650 74.390 ;
        RECT 22.070 71.570 22.390 71.890 ;
        RECT 22.070 71.010 22.390 71.330 ;
        RECT 26.270 71.570 26.590 71.890 ;
        RECT 26.270 71.010 26.590 71.330 ;
        RECT 44.470 71.570 44.790 71.890 ;
        RECT 44.470 71.010 44.790 71.330 ;
        RECT 48.670 71.570 48.990 71.890 ;
        RECT 48.670 71.010 48.990 71.330 ;
        RECT 92.130 71.570 92.450 71.890 ;
        RECT 92.130 71.010 92.450 71.330 ;
        RECT 96.330 71.570 96.650 71.890 ;
        RECT 96.330 71.010 96.650 71.330 ;
        RECT 114.530 71.570 114.850 71.890 ;
        RECT 114.530 71.010 114.850 71.330 ;
        RECT 118.730 71.570 119.050 71.890 ;
        RECT 118.730 71.010 119.050 71.330 ;
        RECT 19.270 68.510 19.590 68.830 ;
        RECT 19.270 67.950 19.590 68.270 ;
        RECT 20.670 68.510 20.990 68.830 ;
        RECT 20.670 67.950 20.990 68.270 ;
        RECT 27.670 68.510 27.990 68.830 ;
        RECT 27.670 67.950 27.990 68.270 ;
        RECT 29.070 68.510 29.390 68.830 ;
        RECT 29.070 67.950 29.390 68.270 ;
        RECT 41.670 68.510 41.990 68.830 ;
        RECT 41.670 67.950 41.990 68.270 ;
        RECT 43.070 68.510 43.390 68.830 ;
        RECT 43.070 67.950 43.390 68.270 ;
        RECT 50.070 68.510 50.390 68.830 ;
        RECT 50.070 67.950 50.390 68.270 ;
        RECT 51.470 68.510 51.790 68.830 ;
        RECT 51.470 67.950 51.790 68.270 ;
        RECT 89.330 68.510 89.650 68.830 ;
        RECT 89.330 67.950 89.650 68.270 ;
        RECT 90.730 68.510 91.050 68.830 ;
        RECT 90.730 67.950 91.050 68.270 ;
        RECT 97.730 68.510 98.050 68.830 ;
        RECT 97.730 67.950 98.050 68.270 ;
        RECT 99.130 68.510 99.450 68.830 ;
        RECT 99.130 67.950 99.450 68.270 ;
        RECT 111.730 68.510 112.050 68.830 ;
        RECT 111.730 67.950 112.050 68.270 ;
        RECT 113.130 68.510 113.450 68.830 ;
        RECT 113.130 67.950 113.450 68.270 ;
        RECT 120.130 68.510 120.450 68.830 ;
        RECT 120.130 67.950 120.450 68.270 ;
        RECT 121.530 68.510 121.850 68.830 ;
        RECT 121.530 67.950 121.850 68.270 ;
        RECT 12.270 66.480 12.590 66.800 ;
        RECT 12.270 65.920 12.590 66.240 ;
        RECT 143.740 82.180 144.060 82.500 ;
        RECT 144.300 82.180 144.620 82.500 ;
        RECT 147.700 82.180 148.020 82.500 ;
        RECT 148.260 82.180 148.580 82.500 ;
        RECT 143.740 78.660 144.060 78.980 ;
        RECT 144.300 78.660 144.620 78.980 ;
        RECT 147.700 78.660 148.020 78.980 ;
        RECT 148.260 78.660 148.580 78.980 ;
        RECT 143.740 76.900 144.060 77.220 ;
        RECT 144.300 76.900 144.620 77.220 ;
        RECT 147.700 76.900 148.020 77.220 ;
        RECT 148.260 76.900 148.580 77.220 ;
        RECT 147.700 76.020 148.020 76.340 ;
        RECT 148.260 76.020 148.580 76.340 ;
        RECT 143.740 73.380 144.060 73.700 ;
        RECT 144.300 73.380 144.620 73.700 ;
        RECT 147.700 73.380 148.020 73.700 ;
        RECT 148.260 73.380 148.580 73.700 ;
        RECT 143.740 71.620 144.060 71.940 ;
        RECT 144.300 71.620 144.620 71.940 ;
        RECT 147.700 71.620 148.020 71.940 ;
        RECT 148.260 71.620 148.580 71.940 ;
        RECT 128.530 66.480 128.850 66.800 ;
        RECT 128.530 65.920 128.850 66.240 ;
        RECT 24.870 65.450 25.190 65.770 ;
        RECT 24.870 64.890 25.190 65.210 ;
        RECT 45.870 65.450 46.190 65.770 ;
        RECT 45.870 64.890 46.190 65.210 ;
        RECT 94.930 65.450 95.250 65.770 ;
        RECT 94.930 64.890 95.250 65.210 ;
        RECT 115.930 65.450 116.250 65.770 ;
        RECT 115.930 64.890 116.250 65.210 ;
        RECT 13.670 62.390 13.990 62.710 ;
        RECT 13.670 61.830 13.990 62.150 ;
        RECT 15.070 62.390 15.390 62.710 ;
        RECT 15.070 61.830 15.390 62.150 ;
        RECT 16.470 62.390 16.790 62.710 ;
        RECT 16.470 61.830 16.790 62.150 ;
        RECT 17.870 62.390 18.190 62.710 ;
        RECT 17.870 61.830 18.190 62.150 ;
        RECT 30.470 62.390 30.790 62.710 ;
        RECT 30.470 61.830 30.790 62.150 ;
        RECT 31.870 62.390 32.190 62.710 ;
        RECT 31.870 61.830 32.190 62.150 ;
        RECT 33.270 62.390 33.590 62.710 ;
        RECT 33.270 61.830 33.590 62.150 ;
        RECT 34.670 62.390 34.990 62.710 ;
        RECT 34.670 61.830 34.990 62.150 ;
        RECT 36.070 62.390 36.390 62.710 ;
        RECT 36.070 61.830 36.390 62.150 ;
        RECT 37.470 62.390 37.790 62.710 ;
        RECT 37.470 61.830 37.790 62.150 ;
        RECT 38.870 62.390 39.190 62.710 ;
        RECT 38.870 61.830 39.190 62.150 ;
        RECT 40.270 62.390 40.590 62.710 ;
        RECT 40.270 61.830 40.590 62.150 ;
        RECT 52.870 62.390 53.190 62.710 ;
        RECT 52.870 61.830 53.190 62.150 ;
        RECT 54.270 62.390 54.590 62.710 ;
        RECT 54.270 61.830 54.590 62.150 ;
        RECT 55.670 62.390 55.990 62.710 ;
        RECT 55.670 61.830 55.990 62.150 ;
        RECT 57.070 62.390 57.390 62.710 ;
        RECT 57.070 61.830 57.390 62.150 ;
        RECT 83.730 62.390 84.050 62.710 ;
        RECT 83.730 61.830 84.050 62.150 ;
        RECT 85.130 62.390 85.450 62.710 ;
        RECT 85.130 61.830 85.450 62.150 ;
        RECT 86.530 62.390 86.850 62.710 ;
        RECT 86.530 61.830 86.850 62.150 ;
        RECT 87.930 62.390 88.250 62.710 ;
        RECT 87.930 61.830 88.250 62.150 ;
        RECT 100.530 62.390 100.850 62.710 ;
        RECT 100.530 61.830 100.850 62.150 ;
        RECT 101.930 62.390 102.250 62.710 ;
        RECT 101.930 61.830 102.250 62.150 ;
        RECT 103.330 62.390 103.650 62.710 ;
        RECT 103.330 61.830 103.650 62.150 ;
        RECT 104.730 62.390 105.050 62.710 ;
        RECT 104.730 61.830 105.050 62.150 ;
        RECT 106.130 62.390 106.450 62.710 ;
        RECT 106.130 61.830 106.450 62.150 ;
        RECT 107.530 62.390 107.850 62.710 ;
        RECT 107.530 61.830 107.850 62.150 ;
        RECT 108.930 62.390 109.250 62.710 ;
        RECT 108.930 61.830 109.250 62.150 ;
        RECT 110.330 62.390 110.650 62.710 ;
        RECT 110.330 61.830 110.650 62.150 ;
        RECT 122.930 62.390 123.250 62.710 ;
        RECT 122.930 61.830 123.250 62.150 ;
        RECT 124.330 62.390 124.650 62.710 ;
        RECT 124.330 61.830 124.650 62.150 ;
        RECT 125.730 62.390 126.050 62.710 ;
        RECT 125.730 61.830 126.050 62.150 ;
        RECT 127.130 62.390 127.450 62.710 ;
        RECT 127.130 61.830 127.450 62.150 ;
        RECT 47.270 59.330 47.590 59.650 ;
        RECT 47.270 58.770 47.590 59.090 ;
        RECT 93.530 59.330 93.850 59.650 ;
        RECT 93.530 58.770 93.850 59.090 ;
        RECT 23.470 57.230 23.790 57.550 ;
        RECT 23.470 56.670 23.790 56.990 ;
        RECT 117.330 57.230 117.650 57.550 ;
        RECT 117.330 56.670 117.650 56.990 ;
        RECT 22.070 54.170 22.390 54.490 ;
        RECT 22.070 53.610 22.390 53.930 ;
        RECT 26.270 54.170 26.590 54.490 ;
        RECT 26.270 53.610 26.590 53.930 ;
        RECT 44.470 54.170 44.790 54.490 ;
        RECT 44.470 53.610 44.790 53.930 ;
        RECT 48.670 54.170 48.990 54.490 ;
        RECT 48.670 53.610 48.990 53.930 ;
        RECT 92.130 54.170 92.450 54.490 ;
        RECT 92.130 53.610 92.450 53.930 ;
        RECT 96.330 54.170 96.650 54.490 ;
        RECT 96.330 53.610 96.650 53.930 ;
        RECT 114.530 54.170 114.850 54.490 ;
        RECT 114.530 53.610 114.850 53.930 ;
        RECT 118.730 54.170 119.050 54.490 ;
        RECT 118.730 53.610 119.050 53.930 ;
        RECT 19.270 51.110 19.590 51.430 ;
        RECT 19.270 50.550 19.590 50.870 ;
        RECT 20.670 51.110 20.990 51.430 ;
        RECT 20.670 50.550 20.990 50.870 ;
        RECT 27.670 51.110 27.990 51.430 ;
        RECT 27.670 50.550 27.990 50.870 ;
        RECT 29.070 51.110 29.390 51.430 ;
        RECT 29.070 50.550 29.390 50.870 ;
        RECT 41.670 51.110 41.990 51.430 ;
        RECT 41.670 50.550 41.990 50.870 ;
        RECT 43.070 51.110 43.390 51.430 ;
        RECT 43.070 50.550 43.390 50.870 ;
        RECT 50.070 51.110 50.390 51.430 ;
        RECT 50.070 50.550 50.390 50.870 ;
        RECT 51.470 51.110 51.790 51.430 ;
        RECT 51.470 50.550 51.790 50.870 ;
        RECT 89.330 51.110 89.650 51.430 ;
        RECT 89.330 50.550 89.650 50.870 ;
        RECT 90.730 51.110 91.050 51.430 ;
        RECT 90.730 50.550 91.050 50.870 ;
        RECT 97.730 51.110 98.050 51.430 ;
        RECT 97.730 50.550 98.050 50.870 ;
        RECT 99.130 51.110 99.450 51.430 ;
        RECT 99.130 50.550 99.450 50.870 ;
        RECT 111.730 51.110 112.050 51.430 ;
        RECT 111.730 50.550 112.050 50.870 ;
        RECT 113.130 51.110 113.450 51.430 ;
        RECT 113.130 50.550 113.450 50.870 ;
        RECT 120.130 51.110 120.450 51.430 ;
        RECT 120.130 50.550 120.450 50.870 ;
        RECT 121.530 51.110 121.850 51.430 ;
        RECT 121.530 50.550 121.850 50.870 ;
        RECT 12.270 49.080 12.590 49.400 ;
        RECT 12.270 48.520 12.590 48.840 ;
        RECT 147.700 68.100 148.020 68.420 ;
        RECT 148.260 68.100 148.580 68.420 ;
        RECT 147.700 67.220 148.020 67.540 ;
        RECT 148.260 67.220 148.580 67.540 ;
        RECT 143.740 66.340 144.060 66.660 ;
        RECT 144.300 66.340 144.620 66.660 ;
        RECT 143.740 62.820 144.060 63.140 ;
        RECT 144.300 62.820 144.620 63.140 ;
        RECT 147.700 62.820 148.020 63.140 ;
        RECT 148.260 62.820 148.580 63.140 ;
        RECT 143.740 61.060 144.060 61.380 ;
        RECT 144.300 61.060 144.620 61.380 ;
        RECT 147.700 61.060 148.020 61.380 ;
        RECT 148.260 61.060 148.580 61.380 ;
        RECT 143.740 57.540 144.060 57.860 ;
        RECT 144.300 57.540 144.620 57.860 ;
        RECT 147.700 57.540 148.020 57.860 ;
        RECT 148.260 57.540 148.580 57.860 ;
        RECT 143.740 54.020 144.060 54.340 ;
        RECT 144.300 54.020 144.620 54.340 ;
        RECT 147.700 54.020 148.020 54.340 ;
        RECT 148.260 54.020 148.580 54.340 ;
        RECT 143.740 52.260 144.060 52.580 ;
        RECT 144.300 52.260 144.620 52.580 ;
        RECT 147.700 52.260 148.020 52.580 ;
        RECT 148.260 52.260 148.580 52.580 ;
        RECT 147.700 51.380 148.020 51.700 ;
        RECT 148.260 51.380 148.580 51.700 ;
        RECT 128.530 49.080 128.850 49.400 ;
        RECT 128.530 48.520 128.850 48.840 ;
        RECT 143.740 48.740 144.060 49.060 ;
        RECT 144.300 48.740 144.620 49.060 ;
        RECT 147.700 48.740 148.020 49.060 ;
        RECT 148.260 48.740 148.580 49.060 ;
        RECT 24.870 48.050 25.190 48.370 ;
        RECT 24.870 47.490 25.190 47.810 ;
        RECT 45.870 48.050 46.190 48.370 ;
        RECT 45.870 47.490 46.190 47.810 ;
        RECT 94.930 48.050 95.250 48.370 ;
        RECT 94.930 47.490 95.250 47.810 ;
        RECT 115.930 48.050 116.250 48.370 ;
        RECT 115.930 47.490 116.250 47.810 ;
        RECT 13.670 44.990 13.990 45.310 ;
        RECT 13.670 44.430 13.990 44.750 ;
        RECT 15.070 44.990 15.390 45.310 ;
        RECT 15.070 44.430 15.390 44.750 ;
        RECT 16.470 44.990 16.790 45.310 ;
        RECT 16.470 44.430 16.790 44.750 ;
        RECT 17.870 44.990 18.190 45.310 ;
        RECT 17.870 44.430 18.190 44.750 ;
        RECT 30.470 44.990 30.790 45.310 ;
        RECT 30.470 44.430 30.790 44.750 ;
        RECT 31.870 44.990 32.190 45.310 ;
        RECT 31.870 44.430 32.190 44.750 ;
        RECT 33.270 44.990 33.590 45.310 ;
        RECT 33.270 44.430 33.590 44.750 ;
        RECT 34.670 44.990 34.990 45.310 ;
        RECT 34.670 44.430 34.990 44.750 ;
        RECT 36.070 44.990 36.390 45.310 ;
        RECT 36.070 44.430 36.390 44.750 ;
        RECT 37.470 44.990 37.790 45.310 ;
        RECT 37.470 44.430 37.790 44.750 ;
        RECT 38.870 44.990 39.190 45.310 ;
        RECT 38.870 44.430 39.190 44.750 ;
        RECT 40.270 44.990 40.590 45.310 ;
        RECT 40.270 44.430 40.590 44.750 ;
        RECT 52.870 44.990 53.190 45.310 ;
        RECT 52.870 44.430 53.190 44.750 ;
        RECT 54.270 44.990 54.590 45.310 ;
        RECT 54.270 44.430 54.590 44.750 ;
        RECT 55.670 44.990 55.990 45.310 ;
        RECT 55.670 44.430 55.990 44.750 ;
        RECT 57.070 44.990 57.390 45.310 ;
        RECT 57.070 44.430 57.390 44.750 ;
        RECT 83.730 44.990 84.050 45.310 ;
        RECT 83.730 44.430 84.050 44.750 ;
        RECT 85.130 44.990 85.450 45.310 ;
        RECT 85.130 44.430 85.450 44.750 ;
        RECT 86.530 44.990 86.850 45.310 ;
        RECT 86.530 44.430 86.850 44.750 ;
        RECT 87.930 44.990 88.250 45.310 ;
        RECT 87.930 44.430 88.250 44.750 ;
        RECT 100.530 44.990 100.850 45.310 ;
        RECT 100.530 44.430 100.850 44.750 ;
        RECT 101.930 44.990 102.250 45.310 ;
        RECT 101.930 44.430 102.250 44.750 ;
        RECT 103.330 44.990 103.650 45.310 ;
        RECT 103.330 44.430 103.650 44.750 ;
        RECT 104.730 44.990 105.050 45.310 ;
        RECT 104.730 44.430 105.050 44.750 ;
        RECT 106.130 44.990 106.450 45.310 ;
        RECT 106.130 44.430 106.450 44.750 ;
        RECT 107.530 44.990 107.850 45.310 ;
        RECT 107.530 44.430 107.850 44.750 ;
        RECT 108.930 44.990 109.250 45.310 ;
        RECT 108.930 44.430 109.250 44.750 ;
        RECT 110.330 44.990 110.650 45.310 ;
        RECT 110.330 44.430 110.650 44.750 ;
        RECT 122.930 44.990 123.250 45.310 ;
        RECT 122.930 44.430 123.250 44.750 ;
        RECT 124.330 44.990 124.650 45.310 ;
        RECT 124.330 44.430 124.650 44.750 ;
        RECT 125.730 44.990 126.050 45.310 ;
        RECT 125.730 44.430 126.050 44.750 ;
        RECT 127.130 44.990 127.450 45.310 ;
        RECT 127.130 44.430 127.450 44.750 ;
        RECT 47.270 41.930 47.590 42.250 ;
        RECT 47.270 41.370 47.590 41.690 ;
        RECT 93.530 41.930 93.850 42.250 ;
        RECT 93.530 41.370 93.850 41.690 ;
        RECT 143.740 46.980 144.060 47.300 ;
        RECT 144.300 46.980 144.620 47.300 ;
        RECT 147.700 46.980 148.020 47.300 ;
        RECT 148.260 46.980 148.580 47.300 ;
        RECT 147.700 43.460 148.020 43.780 ;
        RECT 148.260 43.460 148.580 43.780 ;
        RECT 147.700 42.580 148.020 42.900 ;
        RECT 148.260 42.580 148.580 42.900 ;
        RECT 143.740 41.700 144.060 42.020 ;
        RECT 144.300 41.700 144.620 42.020 ;
        RECT 47.080 38.580 48.160 38.935 ;
        RECT 14.320 37.700 15.400 38.055 ;
        RECT 47.080 36.820 48.160 37.175 ;
        RECT 14.320 35.940 15.400 36.295 ;
        RECT 47.080 35.060 48.160 35.415 ;
        RECT 93.160 38.580 94.240 38.935 ;
        RECT 143.740 38.180 144.060 38.500 ;
        RECT 144.300 38.180 144.620 38.500 ;
        RECT 147.700 38.180 148.020 38.500 ;
        RECT 148.260 38.180 148.580 38.500 ;
        RECT 125.920 37.700 127.000 38.055 ;
        RECT 93.160 36.820 94.240 37.175 ;
        RECT 143.740 36.420 144.060 36.740 ;
        RECT 144.300 36.420 144.620 36.740 ;
        RECT 147.700 36.420 148.020 36.740 ;
        RECT 148.260 36.420 148.580 36.740 ;
        RECT 125.920 35.940 127.000 36.295 ;
        RECT 93.160 35.060 94.240 35.415 ;
        RECT 14.320 34.185 15.400 34.535 ;
        RECT 125.920 34.185 127.000 34.535 ;
        RECT 47.080 33.300 48.160 33.655 ;
        RECT 14.320 32.420 15.400 32.775 ;
        RECT 93.160 33.300 94.240 33.655 ;
        RECT 54.780 32.040 55.100 32.360 ;
        RECT 55.340 32.040 55.660 32.360 ;
        RECT 58.740 32.040 59.060 32.360 ;
        RECT 59.300 32.040 59.620 32.360 ;
        RECT 81.700 32.040 82.020 32.360 ;
        RECT 82.260 32.040 82.580 32.360 ;
        RECT 85.660 32.040 85.980 32.360 ;
        RECT 86.220 32.040 86.540 32.360 ;
        RECT 47.080 31.540 48.160 31.895 ;
        RECT 143.740 32.900 144.060 33.220 ;
        RECT 144.300 32.900 144.620 33.220 ;
        RECT 147.700 32.900 148.020 33.220 ;
        RECT 148.260 32.900 148.580 33.220 ;
        RECT 125.920 32.420 127.000 32.775 ;
        RECT 93.160 31.540 94.240 31.895 ;
        RECT 14.320 30.660 15.400 31.015 ;
        RECT 54.780 31.160 55.100 31.480 ;
        RECT 55.340 31.160 55.660 31.480 ;
        RECT 58.740 31.160 59.060 31.480 ;
        RECT 59.300 31.160 59.620 31.480 ;
        RECT 81.700 31.160 82.020 31.480 ;
        RECT 82.260 31.160 82.580 31.480 ;
        RECT 85.660 31.160 85.980 31.480 ;
        RECT 86.220 31.160 86.540 31.480 ;
        RECT 61.660 30.240 61.980 30.560 ;
        RECT 62.220 30.240 62.540 30.560 ;
        RECT 78.780 30.240 79.100 30.560 ;
        RECT 79.340 30.240 79.660 30.560 ;
        RECT 47.080 29.780 48.160 30.135 ;
        RECT 125.920 30.660 127.000 31.015 ;
        RECT 93.160 29.780 94.240 30.135 ;
        RECT 54.780 29.400 55.100 29.720 ;
        RECT 55.340 29.400 55.660 29.720 ;
        RECT 58.740 29.400 59.060 29.720 ;
        RECT 59.300 29.400 59.620 29.720 ;
        RECT 81.700 29.400 82.020 29.720 ;
        RECT 82.260 29.400 82.580 29.720 ;
        RECT 85.660 29.400 85.980 29.720 ;
        RECT 86.220 29.400 86.540 29.720 ;
        RECT 143.740 29.380 144.060 29.700 ;
        RECT 144.300 29.380 144.620 29.700 ;
        RECT 147.700 29.380 148.020 29.700 ;
        RECT 148.260 29.380 148.580 29.700 ;
        RECT 14.320 28.905 15.400 29.255 ;
        RECT 125.920 28.905 127.000 29.255 ;
        RECT 54.780 28.520 55.100 28.840 ;
        RECT 55.340 28.520 55.660 28.840 ;
        RECT 58.740 28.520 59.060 28.840 ;
        RECT 59.300 28.520 59.620 28.840 ;
        RECT 81.700 28.520 82.020 28.840 ;
        RECT 82.260 28.520 82.580 28.840 ;
        RECT 85.660 28.520 85.980 28.840 ;
        RECT 86.220 28.520 86.540 28.840 ;
        RECT 47.080 28.020 48.160 28.375 ;
        RECT 93.160 28.020 94.240 28.375 ;
        RECT 14.320 27.140 15.400 27.495 ;
        RECT 54.780 27.640 55.100 27.960 ;
        RECT 55.340 27.640 55.660 27.960 ;
        RECT 58.740 27.640 59.060 27.960 ;
        RECT 59.300 27.640 59.620 27.960 ;
        RECT 81.700 27.640 82.020 27.960 ;
        RECT 82.260 27.640 82.580 27.960 ;
        RECT 85.660 27.640 85.980 27.960 ;
        RECT 86.220 27.640 86.540 27.960 ;
        RECT 47.080 26.260 48.160 26.615 ;
        RECT 143.740 27.620 144.060 27.940 ;
        RECT 144.300 27.620 144.620 27.940 ;
        RECT 147.700 27.620 148.020 27.940 ;
        RECT 148.260 27.620 148.580 27.940 ;
        RECT 125.920 27.140 127.000 27.495 ;
        RECT 93.160 26.260 94.240 26.615 ;
        RECT 14.320 25.380 15.400 25.735 ;
        RECT 54.780 25.880 55.100 26.200 ;
        RECT 55.340 25.880 55.660 26.200 ;
        RECT 58.740 25.880 59.060 26.200 ;
        RECT 59.300 25.880 59.620 26.200 ;
        RECT 74.500 25.880 74.820 26.200 ;
        RECT 75.060 25.880 75.380 26.200 ;
        RECT 81.700 25.880 82.020 26.200 ;
        RECT 82.260 25.880 82.580 26.200 ;
        RECT 85.660 25.880 85.980 26.200 ;
        RECT 86.220 25.880 86.540 26.200 ;
        RECT 54.780 25.000 55.100 25.320 ;
        RECT 55.340 25.000 55.660 25.320 ;
        RECT 47.080 24.500 48.160 24.855 ;
        RECT 14.320 23.625 15.400 23.975 ;
        RECT 52.620 23.240 52.940 23.560 ;
        RECT 53.180 23.240 53.500 23.560 ;
        RECT 47.080 22.740 48.160 23.095 ;
        RECT 14.320 21.860 15.400 22.215 ;
        RECT 58.740 22.360 59.060 22.680 ;
        RECT 59.300 22.360 59.620 22.680 ;
        RECT 47.080 20.980 48.160 21.335 ;
        RECT 14.320 20.100 15.400 20.455 ;
        RECT 47.080 19.220 48.160 19.575 ;
        RECT 52.620 19.280 52.940 19.600 ;
        RECT 53.180 19.280 53.500 19.600 ;
        RECT 14.320 18.345 15.400 18.695 ;
        RECT 47.080 17.460 48.160 17.815 ;
        RECT 14.320 16.580 15.400 16.935 ;
        RECT 47.080 15.700 48.160 16.055 ;
        RECT 14.320 14.820 15.400 15.175 ;
        RECT 47.080 13.940 48.160 14.295 ;
        RECT 14.320 13.065 15.400 13.415 ;
        RECT 54.780 18.840 55.100 19.160 ;
        RECT 55.340 18.840 55.660 19.160 ;
        RECT 58.740 18.840 59.060 19.160 ;
        RECT 59.300 18.840 59.620 19.160 ;
        RECT 54.780 17.960 55.100 18.280 ;
        RECT 55.340 17.960 55.660 18.280 ;
        RECT 58.740 17.960 59.060 18.280 ;
        RECT 59.300 17.960 59.620 18.280 ;
        RECT 85.660 25.000 85.980 25.320 ;
        RECT 86.220 25.000 86.540 25.320 ;
        RECT 65.860 18.840 66.180 19.160 ;
        RECT 66.420 18.840 66.740 19.160 ;
        RECT 74.500 18.840 74.820 19.160 ;
        RECT 75.060 18.840 75.380 19.160 ;
        RECT 147.700 26.740 148.020 27.060 ;
        RECT 148.260 26.740 148.580 27.060 ;
        RECT 125.920 25.380 127.000 25.735 ;
        RECT 93.160 24.500 94.240 24.855 ;
        RECT 143.740 24.100 144.060 24.420 ;
        RECT 144.300 24.100 144.620 24.420 ;
        RECT 147.700 24.100 148.020 24.420 ;
        RECT 148.260 24.100 148.580 24.420 ;
        RECT 125.920 23.625 127.000 23.975 ;
        RECT 87.820 23.240 88.140 23.560 ;
        RECT 88.380 23.240 88.700 23.560 ;
        RECT 93.160 22.740 94.240 23.095 ;
        RECT 81.700 22.360 82.020 22.680 ;
        RECT 82.260 22.360 82.580 22.680 ;
        RECT 143.740 22.340 144.060 22.660 ;
        RECT 144.300 22.340 144.620 22.660 ;
        RECT 147.700 22.340 148.020 22.660 ;
        RECT 148.260 22.340 148.580 22.660 ;
        RECT 125.920 21.860 127.000 22.215 ;
        RECT 93.160 20.980 94.240 21.335 ;
        RECT 81.700 18.840 82.020 19.160 ;
        RECT 82.260 18.840 82.580 19.160 ;
        RECT 85.660 18.840 85.980 19.160 ;
        RECT 86.220 18.840 86.540 19.160 ;
        RECT 81.700 17.960 82.020 18.280 ;
        RECT 82.260 17.960 82.580 18.280 ;
        RECT 85.660 17.960 85.980 18.280 ;
        RECT 86.220 17.960 86.540 18.280 ;
        RECT 54.780 15.320 55.100 15.640 ;
        RECT 55.340 15.320 55.660 15.640 ;
        RECT 58.740 15.320 59.060 15.640 ;
        RECT 59.300 15.320 59.620 15.640 ;
        RECT 81.700 15.320 82.020 15.640 ;
        RECT 82.260 15.320 82.580 15.640 ;
        RECT 85.660 15.320 85.980 15.640 ;
        RECT 86.220 15.320 86.540 15.640 ;
        RECT 54.780 14.440 55.100 14.760 ;
        RECT 55.340 14.440 55.660 14.760 ;
        RECT 58.740 14.440 59.060 14.760 ;
        RECT 59.300 14.440 59.620 14.760 ;
        RECT 65.860 14.400 66.180 14.720 ;
        RECT 66.420 14.400 66.740 14.720 ;
        RECT 74.580 14.400 74.900 14.720 ;
        RECT 75.140 14.400 75.460 14.720 ;
        RECT 81.700 14.440 82.020 14.760 ;
        RECT 82.260 14.440 82.580 14.760 ;
        RECT 85.660 14.440 85.980 14.760 ;
        RECT 86.220 14.440 86.540 14.760 ;
        RECT 54.780 13.560 55.100 13.880 ;
        RECT 55.340 13.560 55.660 13.880 ;
        RECT 58.740 13.560 59.060 13.880 ;
        RECT 59.300 13.560 59.620 13.880 ;
        RECT 81.700 13.560 82.020 13.880 ;
        RECT 82.260 13.560 82.580 13.880 ;
        RECT 85.660 13.560 85.980 13.880 ;
        RECT 86.220 13.560 86.540 13.880 ;
        RECT 48.300 13.050 48.620 13.370 ;
        RECT 48.860 13.050 49.180 13.370 ;
        RECT 87.820 19.280 88.140 19.600 ;
        RECT 88.380 19.280 88.700 19.600 ;
        RECT 147.700 21.460 148.020 21.780 ;
        RECT 148.260 21.460 148.580 21.780 ;
        RECT 125.920 20.100 127.000 20.455 ;
        RECT 93.160 19.220 94.240 19.575 ;
        RECT 143.740 18.820 144.060 19.140 ;
        RECT 144.300 18.820 144.620 19.140 ;
        RECT 147.700 18.820 148.020 19.140 ;
        RECT 148.260 18.820 148.580 19.140 ;
        RECT 125.920 18.345 127.000 18.695 ;
        RECT 93.160 17.460 94.240 17.815 ;
        RECT 143.740 17.060 144.060 17.380 ;
        RECT 144.300 17.060 144.620 17.380 ;
        RECT 147.700 17.060 148.020 17.380 ;
        RECT 148.260 17.060 148.580 17.380 ;
        RECT 125.920 16.580 127.000 16.935 ;
        RECT 93.160 15.700 94.240 16.055 ;
        RECT 143.740 15.300 144.060 15.620 ;
        RECT 144.300 15.300 144.620 15.620 ;
        RECT 147.700 15.300 148.020 15.620 ;
        RECT 148.260 15.300 148.580 15.620 ;
        RECT 125.920 14.820 127.000 15.175 ;
        RECT 93.160 13.940 94.240 14.295 ;
        RECT 143.740 14.420 144.060 14.740 ;
        RECT 144.300 14.420 144.620 14.740 ;
        RECT 92.140 13.050 92.460 13.370 ;
        RECT 92.700 13.050 93.020 13.370 ;
        RECT 125.920 13.065 127.000 13.415 ;
        RECT 143.740 11.780 144.060 12.100 ;
        RECT 144.300 11.780 144.620 12.100 ;
        RECT 147.700 11.780 148.020 12.100 ;
        RECT 148.260 11.780 148.580 12.100 ;
        RECT 58.740 10.260 59.060 10.580 ;
        RECT 59.300 10.260 59.620 10.580 ;
        RECT 58.740 9.700 59.060 10.020 ;
        RECT 59.300 9.700 59.620 10.020 ;
        RECT 81.700 10.260 82.020 10.580 ;
        RECT 82.260 10.260 82.580 10.580 ;
        RECT 81.700 9.700 82.020 10.020 ;
        RECT 82.260 9.700 82.580 10.020 ;
        RECT 143.740 10.020 144.060 10.340 ;
        RECT 144.300 10.020 144.620 10.340 ;
        RECT 147.700 10.020 148.020 10.340 ;
        RECT 148.260 10.020 148.580 10.340 ;
        RECT 143.740 9.140 144.060 9.460 ;
        RECT 144.300 9.140 144.620 9.460 ;
        RECT 147.700 9.140 148.020 9.460 ;
        RECT 148.260 9.140 148.580 9.460 ;
        RECT 54.780 6.660 55.100 6.980 ;
        RECT 55.340 6.660 55.660 6.980 ;
        RECT 54.780 6.100 55.100 6.420 ;
        RECT 55.340 6.100 55.660 6.420 ;
        RECT 85.660 6.660 85.980 6.980 ;
        RECT 86.220 6.660 86.540 6.980 ;
        RECT 143.740 6.500 144.060 6.820 ;
        RECT 144.300 6.500 144.620 6.820 ;
        RECT 147.700 6.500 148.020 6.820 ;
        RECT 148.260 6.500 148.580 6.820 ;
        RECT 85.660 6.100 85.980 6.420 ;
        RECT 86.220 6.100 86.540 6.420 ;
        RECT 143.740 4.740 144.060 5.060 ;
        RECT 144.300 4.740 144.620 5.060 ;
        RECT 147.700 4.740 148.020 5.060 ;
        RECT 148.260 4.740 148.580 5.060 ;
        RECT 61.660 4.030 61.980 4.350 ;
        RECT 62.220 4.030 62.540 4.350 ;
        RECT 78.780 4.030 79.100 4.350 ;
        RECT 79.340 4.030 79.660 4.350 ;
        RECT 143.740 3.860 144.060 4.180 ;
        RECT 144.300 3.860 144.620 4.180 ;
        RECT 147.700 3.860 148.020 4.180 ;
        RECT 148.260 3.860 148.580 4.180 ;
        RECT 143.740 2.980 144.060 3.300 ;
        RECT 144.300 2.980 144.620 3.300 ;
        RECT 147.700 2.980 148.020 3.300 ;
        RECT 148.260 2.980 148.580 3.300 ;
      LAYER met3 ;
        RECT 15.660 168.080 16.660 168.460 ;
        RECT 15.660 116.610 16.040 168.080 ;
        RECT 17.740 139.230 18.740 214.990 ;
        RECT 19.235 119.520 19.615 169.210 ;
        RECT 20.035 126.310 20.415 176.250 ;
        RECT 20.910 129.220 21.290 183.290 ;
        RECT 21.700 139.230 22.700 218.590 ;
        RECT 24.580 163.280 25.580 222.190 ;
        RECT 27.540 163.280 28.540 222.190 ;
        RECT 30.420 139.230 31.420 218.590 ;
        RECT 31.830 130.190 32.210 183.290 ;
        RECT 32.705 175.250 33.085 176.250 ;
        RECT 32.700 127.280 33.080 175.250 ;
        RECT 33.505 168.210 33.885 169.210 ;
        RECT 33.500 120.490 33.880 168.210 ;
        RECT 34.380 139.230 35.380 214.990 ;
        RECT 36.460 168.080 37.460 168.460 ;
        RECT 40.860 168.080 41.860 168.460 ;
        RECT 36.460 117.580 36.840 168.080 ;
        RECT 40.860 118.550 41.240 168.080 ;
        RECT 42.940 139.230 43.940 214.990 ;
        RECT 44.435 121.460 44.815 169.210 ;
        RECT 45.235 128.250 45.615 176.250 ;
        RECT 46.110 131.160 46.490 183.290 ;
        RECT 46.900 139.230 47.900 218.590 ;
        RECT 49.780 163.280 50.780 222.190 ;
        RECT 52.740 163.280 53.740 222.190 ;
        RECT 55.620 139.230 56.620 218.590 ;
        RECT 57.030 132.130 57.410 183.290 ;
        RECT 57.905 175.250 58.285 176.250 ;
        RECT 58.705 168.210 59.085 169.210 ;
        RECT 58.700 122.430 59.080 168.210 ;
        RECT 59.580 139.230 60.580 214.990 ;
        RECT 61.660 168.080 62.660 168.460 ;
        RECT 66.060 168.080 67.060 168.460 ;
        RECT 68.140 139.230 69.140 214.990 ;
        RECT 70.435 175.250 70.815 176.250 ;
        RECT 69.635 123.400 70.015 169.210 ;
        RECT 71.310 133.100 71.690 183.290 ;
        RECT 72.100 139.230 73.100 218.590 ;
        RECT 74.980 163.280 75.980 222.190 ;
        RECT 77.940 163.280 78.940 222.190 ;
        RECT 80.820 139.230 81.820 218.590 ;
        RECT 82.230 134.070 82.610 183.290 ;
        RECT 83.105 175.250 83.485 176.250 ;
        RECT 83.905 168.210 84.285 169.210 ;
        RECT 83.900 124.370 84.280 168.210 ;
        RECT 84.780 139.230 85.780 214.990 ;
        RECT 86.860 168.080 87.860 168.460 ;
        RECT 91.260 168.080 92.260 168.460 ;
        RECT 93.340 139.230 94.340 214.990 ;
        RECT 95.635 175.250 96.015 176.250 ;
        RECT 94.835 125.340 95.215 169.210 ;
        RECT 96.510 135.040 96.890 183.290 ;
        RECT 97.300 139.230 98.300 218.590 ;
        RECT 100.180 163.280 101.180 222.190 ;
        RECT 103.140 163.280 104.140 222.190 ;
        RECT 106.020 139.230 107.020 218.590 ;
        RECT 107.430 182.290 107.810 183.290 ;
        RECT 108.305 175.250 108.685 176.250 ;
        RECT 109.100 168.210 109.485 169.210 ;
        RECT 109.980 139.230 110.980 214.990 ;
        RECT 117.160 182.200 118.160 182.580 ;
        RECT 112.060 168.080 113.060 168.460 ;
        RECT 116.380 150.520 117.380 150.900 ;
        RECT 116.380 116.880 116.760 150.520 ;
        RECT 117.780 116.880 118.160 182.200 ;
        RECT 118.540 139.230 119.540 214.990 ;
        RECT 122.500 177.740 123.500 218.590 ;
        RECT 122.500 177.360 124.320 177.740 ;
        RECT 122.500 158.380 123.500 177.360 ;
        RECT 123.940 177.300 124.320 177.360 ;
        RECT 123.940 176.920 125.660 177.300 ;
        RECT 122.500 158.000 124.320 158.380 ;
        RECT 122.500 139.230 123.500 158.000 ;
        RECT 123.940 157.940 124.320 158.000 ;
        RECT 123.940 157.560 125.660 157.940 ;
        RECT 57.740 114.980 127.350 115.360 ;
        RECT 57.740 113.040 127.350 113.420 ;
        RECT 57.740 110.510 58.120 111.510 ;
        RECT 12.240 40.610 12.620 110.510 ;
        RECT 12.940 110.130 58.120 110.510 ;
        RECT 12.940 93.190 13.320 110.130 ;
        RECT 13.640 93.510 14.020 109.810 ;
        RECT 14.340 93.190 14.720 110.130 ;
        RECT 15.040 93.510 15.420 109.810 ;
        RECT 15.740 93.190 16.120 110.130 ;
        RECT 16.440 93.510 16.820 109.810 ;
        RECT 17.140 93.190 17.520 110.130 ;
        RECT 17.840 93.510 18.220 109.810 ;
        RECT 18.540 93.190 18.920 110.130 ;
        RECT 19.240 93.510 19.620 109.810 ;
        RECT 19.940 93.190 20.320 110.130 ;
        RECT 20.640 93.510 21.020 109.810 ;
        RECT 21.340 93.190 21.720 110.130 ;
        RECT 22.040 93.510 22.420 109.810 ;
        RECT 22.740 93.190 23.120 110.130 ;
        RECT 23.440 93.510 23.820 109.810 ;
        RECT 24.140 93.190 24.520 110.130 ;
        RECT 24.840 93.510 25.220 109.810 ;
        RECT 25.540 93.190 25.920 110.130 ;
        RECT 26.240 93.510 26.620 109.810 ;
        RECT 26.940 93.190 27.320 110.130 ;
        RECT 27.640 93.510 28.020 109.810 ;
        RECT 28.340 93.190 28.720 110.130 ;
        RECT 29.040 93.510 29.420 109.810 ;
        RECT 29.740 93.190 30.120 110.130 ;
        RECT 30.440 93.510 30.820 109.810 ;
        RECT 31.140 93.190 31.520 110.130 ;
        RECT 31.840 93.510 32.220 109.810 ;
        RECT 32.540 93.190 32.920 110.130 ;
        RECT 33.240 93.510 33.620 109.810 ;
        RECT 33.940 93.190 34.320 110.130 ;
        RECT 34.640 93.510 35.020 109.810 ;
        RECT 35.340 93.190 35.720 110.130 ;
        RECT 36.040 93.510 36.420 109.810 ;
        RECT 36.740 93.190 37.120 110.130 ;
        RECT 37.440 93.510 37.820 109.810 ;
        RECT 38.140 93.190 38.520 110.130 ;
        RECT 38.840 93.510 39.220 109.810 ;
        RECT 39.540 93.190 39.920 110.130 ;
        RECT 40.240 93.510 40.620 109.810 ;
        RECT 40.940 93.190 41.320 110.130 ;
        RECT 41.640 93.510 42.020 109.810 ;
        RECT 42.340 93.190 42.720 110.130 ;
        RECT 43.040 93.510 43.420 109.810 ;
        RECT 43.740 93.190 44.120 110.130 ;
        RECT 44.440 93.510 44.820 109.810 ;
        RECT 45.140 93.190 45.520 110.130 ;
        RECT 45.840 93.510 46.220 109.810 ;
        RECT 46.540 93.190 46.920 110.130 ;
        RECT 47.240 93.510 47.620 109.810 ;
        RECT 47.940 93.190 48.320 110.130 ;
        RECT 48.640 93.510 49.020 109.810 ;
        RECT 49.340 93.190 49.720 110.130 ;
        RECT 50.040 93.510 50.420 109.810 ;
        RECT 50.740 93.190 51.120 110.130 ;
        RECT 51.440 93.510 51.820 109.810 ;
        RECT 52.140 93.190 52.520 110.130 ;
        RECT 52.840 93.510 53.220 109.810 ;
        RECT 53.540 93.190 53.920 110.130 ;
        RECT 54.240 93.510 54.620 109.810 ;
        RECT 54.940 93.190 55.320 110.130 ;
        RECT 55.640 93.510 56.020 109.810 ;
        RECT 56.340 93.190 56.720 110.130 ;
        RECT 57.040 93.510 57.420 109.810 ;
        RECT 57.740 93.190 58.120 110.130 ;
        RECT 12.940 92.730 58.120 93.190 ;
        RECT 12.940 75.790 13.320 92.730 ;
        RECT 13.640 76.110 14.020 92.410 ;
        RECT 14.340 75.790 14.720 92.730 ;
        RECT 15.040 76.110 15.420 92.410 ;
        RECT 15.740 75.790 16.120 92.730 ;
        RECT 16.440 76.110 16.820 92.410 ;
        RECT 17.140 75.790 17.520 92.730 ;
        RECT 17.840 76.110 18.220 92.410 ;
        RECT 18.540 75.790 18.920 92.730 ;
        RECT 19.240 76.110 19.620 92.410 ;
        RECT 19.940 75.790 20.320 92.730 ;
        RECT 20.640 76.110 21.020 92.410 ;
        RECT 21.340 75.790 21.720 92.730 ;
        RECT 22.040 76.110 22.420 92.410 ;
        RECT 22.740 75.790 23.120 92.730 ;
        RECT 23.440 76.110 23.820 92.410 ;
        RECT 24.140 75.790 24.520 92.730 ;
        RECT 24.840 76.110 25.220 92.410 ;
        RECT 25.540 75.790 25.920 92.730 ;
        RECT 26.240 76.110 26.620 92.410 ;
        RECT 26.940 75.790 27.320 92.730 ;
        RECT 27.640 76.110 28.020 92.410 ;
        RECT 28.340 75.790 28.720 92.730 ;
        RECT 29.040 76.110 29.420 92.410 ;
        RECT 29.740 75.790 30.120 92.730 ;
        RECT 30.440 76.110 30.820 92.410 ;
        RECT 31.140 75.790 31.520 92.730 ;
        RECT 31.840 76.110 32.220 92.410 ;
        RECT 32.540 75.790 32.920 92.730 ;
        RECT 33.240 76.110 33.620 92.410 ;
        RECT 33.940 75.790 34.320 92.730 ;
        RECT 34.640 76.110 35.020 92.410 ;
        RECT 35.340 75.790 35.720 92.730 ;
        RECT 36.040 76.110 36.420 92.410 ;
        RECT 36.740 75.790 37.120 92.730 ;
        RECT 37.440 76.110 37.820 92.410 ;
        RECT 38.140 75.790 38.520 92.730 ;
        RECT 38.840 76.110 39.220 92.410 ;
        RECT 39.540 75.790 39.920 92.730 ;
        RECT 40.240 76.110 40.620 92.410 ;
        RECT 40.940 75.790 41.320 92.730 ;
        RECT 41.640 76.110 42.020 92.410 ;
        RECT 42.340 75.790 42.720 92.730 ;
        RECT 43.040 76.110 43.420 92.410 ;
        RECT 43.740 75.790 44.120 92.730 ;
        RECT 44.440 76.110 44.820 92.410 ;
        RECT 45.140 75.790 45.520 92.730 ;
        RECT 45.840 76.110 46.220 92.410 ;
        RECT 46.540 75.790 46.920 92.730 ;
        RECT 47.240 76.110 47.620 92.410 ;
        RECT 47.940 75.790 48.320 92.730 ;
        RECT 48.640 76.110 49.020 92.410 ;
        RECT 49.340 75.790 49.720 92.730 ;
        RECT 50.040 76.110 50.420 92.410 ;
        RECT 50.740 75.790 51.120 92.730 ;
        RECT 51.440 76.110 51.820 92.410 ;
        RECT 52.140 75.790 52.520 92.730 ;
        RECT 52.840 76.110 53.220 92.410 ;
        RECT 53.540 75.790 53.920 92.730 ;
        RECT 54.240 76.110 54.620 92.410 ;
        RECT 54.940 75.790 55.320 92.730 ;
        RECT 55.640 76.110 56.020 92.410 ;
        RECT 56.340 75.790 56.720 92.730 ;
        RECT 57.040 76.110 57.420 92.410 ;
        RECT 57.740 75.790 58.120 92.730 ;
        RECT 12.940 75.330 58.120 75.790 ;
        RECT 12.940 58.390 13.320 75.330 ;
        RECT 13.640 58.710 14.020 75.010 ;
        RECT 14.340 58.390 14.720 75.330 ;
        RECT 15.040 58.710 15.420 75.010 ;
        RECT 15.740 58.390 16.120 75.330 ;
        RECT 16.440 58.710 16.820 75.010 ;
        RECT 17.140 58.390 17.520 75.330 ;
        RECT 17.840 58.710 18.220 75.010 ;
        RECT 18.540 58.390 18.920 75.330 ;
        RECT 19.240 58.710 19.620 75.010 ;
        RECT 19.940 58.390 20.320 75.330 ;
        RECT 20.640 58.710 21.020 75.010 ;
        RECT 21.340 58.390 21.720 75.330 ;
        RECT 22.040 58.710 22.420 75.010 ;
        RECT 22.740 58.390 23.120 75.330 ;
        RECT 23.440 58.710 23.820 75.010 ;
        RECT 24.140 58.390 24.520 75.330 ;
        RECT 24.840 58.710 25.220 75.010 ;
        RECT 25.540 58.390 25.920 75.330 ;
        RECT 26.240 58.710 26.620 75.010 ;
        RECT 26.940 58.390 27.320 75.330 ;
        RECT 27.640 58.710 28.020 75.010 ;
        RECT 28.340 58.390 28.720 75.330 ;
        RECT 29.040 58.710 29.420 75.010 ;
        RECT 29.740 58.390 30.120 75.330 ;
        RECT 30.440 58.710 30.820 75.010 ;
        RECT 31.140 58.390 31.520 75.330 ;
        RECT 31.840 58.710 32.220 75.010 ;
        RECT 32.540 58.390 32.920 75.330 ;
        RECT 33.240 58.710 33.620 75.010 ;
        RECT 33.940 58.390 34.320 75.330 ;
        RECT 34.640 58.710 35.020 75.010 ;
        RECT 35.340 58.390 35.720 75.330 ;
        RECT 36.040 58.710 36.420 75.010 ;
        RECT 36.740 58.390 37.120 75.330 ;
        RECT 37.440 58.710 37.820 75.010 ;
        RECT 38.140 58.390 38.520 75.330 ;
        RECT 38.840 58.710 39.220 75.010 ;
        RECT 39.540 58.390 39.920 75.330 ;
        RECT 40.240 58.710 40.620 75.010 ;
        RECT 40.940 58.390 41.320 75.330 ;
        RECT 41.640 58.710 42.020 75.010 ;
        RECT 42.340 58.390 42.720 75.330 ;
        RECT 43.040 58.710 43.420 75.010 ;
        RECT 43.740 58.390 44.120 75.330 ;
        RECT 44.440 58.710 44.820 75.010 ;
        RECT 45.140 58.390 45.520 75.330 ;
        RECT 45.840 58.710 46.220 75.010 ;
        RECT 46.540 58.390 46.920 75.330 ;
        RECT 47.240 58.710 47.620 75.010 ;
        RECT 47.940 58.390 48.320 75.330 ;
        RECT 48.640 58.710 49.020 75.010 ;
        RECT 49.340 58.390 49.720 75.330 ;
        RECT 50.040 58.710 50.420 75.010 ;
        RECT 50.740 58.390 51.120 75.330 ;
        RECT 51.440 58.710 51.820 75.010 ;
        RECT 52.140 58.390 52.520 75.330 ;
        RECT 52.840 58.710 53.220 75.010 ;
        RECT 53.540 58.390 53.920 75.330 ;
        RECT 54.240 58.710 54.620 75.010 ;
        RECT 54.940 58.390 55.320 75.330 ;
        RECT 55.640 58.710 56.020 75.010 ;
        RECT 56.340 58.390 56.720 75.330 ;
        RECT 57.040 58.710 57.420 75.010 ;
        RECT 57.740 58.390 58.120 75.330 ;
        RECT 12.940 57.930 58.120 58.390 ;
        RECT 12.940 40.990 13.320 57.930 ;
        RECT 13.640 41.310 14.020 57.610 ;
        RECT 14.340 40.990 14.720 57.930 ;
        RECT 15.040 41.310 15.420 57.610 ;
        RECT 15.740 40.990 16.120 57.930 ;
        RECT 16.440 41.310 16.820 57.610 ;
        RECT 17.140 40.990 17.520 57.930 ;
        RECT 17.840 41.310 18.220 57.610 ;
        RECT 18.540 40.990 18.920 57.930 ;
        RECT 19.240 41.310 19.620 57.610 ;
        RECT 19.940 40.990 20.320 57.930 ;
        RECT 20.640 41.310 21.020 57.610 ;
        RECT 21.340 40.990 21.720 57.930 ;
        RECT 22.040 41.310 22.420 57.610 ;
        RECT 22.740 40.990 23.120 57.930 ;
        RECT 23.440 41.310 23.820 57.610 ;
        RECT 24.140 40.990 24.520 57.930 ;
        RECT 24.840 41.310 25.220 57.610 ;
        RECT 25.540 40.990 25.920 57.930 ;
        RECT 26.240 41.310 26.620 57.610 ;
        RECT 26.940 40.990 27.320 57.930 ;
        RECT 27.640 41.310 28.020 57.610 ;
        RECT 28.340 40.990 28.720 57.930 ;
        RECT 29.040 41.310 29.420 57.610 ;
        RECT 29.740 40.990 30.120 57.930 ;
        RECT 30.440 41.310 30.820 57.610 ;
        RECT 31.140 40.990 31.520 57.930 ;
        RECT 31.840 41.310 32.220 57.610 ;
        RECT 32.540 40.990 32.920 57.930 ;
        RECT 33.240 41.310 33.620 57.610 ;
        RECT 33.940 40.990 34.320 57.930 ;
        RECT 34.640 41.310 35.020 57.610 ;
        RECT 35.340 40.990 35.720 57.930 ;
        RECT 36.040 41.310 36.420 57.610 ;
        RECT 36.740 40.990 37.120 57.930 ;
        RECT 37.440 41.310 37.820 57.610 ;
        RECT 38.140 40.990 38.520 57.930 ;
        RECT 38.840 41.310 39.220 57.610 ;
        RECT 39.540 40.990 39.920 57.930 ;
        RECT 40.240 41.310 40.620 57.610 ;
        RECT 40.940 40.990 41.320 57.930 ;
        RECT 41.640 41.310 42.020 57.610 ;
        RECT 42.340 40.990 42.720 57.930 ;
        RECT 43.040 41.310 43.420 57.610 ;
        RECT 43.740 40.990 44.120 57.930 ;
        RECT 44.440 41.310 44.820 57.610 ;
        RECT 45.140 40.990 45.520 57.930 ;
        RECT 45.840 41.310 46.220 57.610 ;
        RECT 46.540 40.990 46.920 57.930 ;
        RECT 47.240 41.310 47.620 57.610 ;
        RECT 47.940 40.990 48.320 57.930 ;
        RECT 48.640 41.310 49.020 57.610 ;
        RECT 49.340 40.990 49.720 57.930 ;
        RECT 50.040 41.310 50.420 57.610 ;
        RECT 50.740 40.990 51.120 57.930 ;
        RECT 51.440 41.310 51.820 57.610 ;
        RECT 52.140 40.990 52.520 57.930 ;
        RECT 52.840 41.310 53.220 57.610 ;
        RECT 53.540 40.990 53.920 57.930 ;
        RECT 54.240 41.310 54.620 57.610 ;
        RECT 54.940 40.990 55.320 57.930 ;
        RECT 55.640 41.310 56.020 57.610 ;
        RECT 56.340 40.990 56.720 57.930 ;
        RECT 57.040 41.310 57.420 57.610 ;
        RECT 57.740 40.990 58.120 57.930 ;
        RECT 83.000 110.510 83.380 111.510 ;
        RECT 83.000 110.130 128.180 110.510 ;
        RECT 83.000 93.190 83.380 110.130 ;
        RECT 83.700 93.510 84.080 109.810 ;
        RECT 84.400 93.190 84.780 110.130 ;
        RECT 85.100 93.510 85.480 109.810 ;
        RECT 85.800 93.190 86.180 110.130 ;
        RECT 86.500 93.510 86.880 109.810 ;
        RECT 87.200 93.190 87.580 110.130 ;
        RECT 87.900 93.510 88.280 109.810 ;
        RECT 88.600 93.190 88.980 110.130 ;
        RECT 89.300 93.510 89.680 109.810 ;
        RECT 90.000 93.190 90.380 110.130 ;
        RECT 90.700 93.510 91.080 109.810 ;
        RECT 91.400 93.190 91.780 110.130 ;
        RECT 92.100 93.510 92.480 109.810 ;
        RECT 92.800 93.190 93.180 110.130 ;
        RECT 93.500 93.510 93.880 109.810 ;
        RECT 94.200 93.190 94.580 110.130 ;
        RECT 94.900 93.510 95.280 109.810 ;
        RECT 95.600 93.190 95.980 110.130 ;
        RECT 96.300 93.510 96.680 109.810 ;
        RECT 97.000 93.190 97.380 110.130 ;
        RECT 97.700 93.510 98.080 109.810 ;
        RECT 98.400 93.190 98.780 110.130 ;
        RECT 99.100 93.510 99.480 109.810 ;
        RECT 99.800 93.190 100.180 110.130 ;
        RECT 100.500 93.510 100.880 109.810 ;
        RECT 101.200 93.190 101.580 110.130 ;
        RECT 101.900 93.510 102.280 109.810 ;
        RECT 102.600 93.190 102.980 110.130 ;
        RECT 103.300 93.510 103.680 109.810 ;
        RECT 104.000 93.190 104.380 110.130 ;
        RECT 104.700 93.510 105.080 109.810 ;
        RECT 105.400 93.190 105.780 110.130 ;
        RECT 106.100 93.510 106.480 109.810 ;
        RECT 106.800 93.190 107.180 110.130 ;
        RECT 107.500 93.510 107.880 109.810 ;
        RECT 108.200 93.190 108.580 110.130 ;
        RECT 108.900 93.510 109.280 109.810 ;
        RECT 109.600 93.190 109.980 110.130 ;
        RECT 110.300 93.510 110.680 109.810 ;
        RECT 111.000 93.190 111.380 110.130 ;
        RECT 111.700 93.510 112.080 109.810 ;
        RECT 112.400 93.190 112.780 110.130 ;
        RECT 113.100 93.510 113.480 109.810 ;
        RECT 113.800 93.190 114.180 110.130 ;
        RECT 114.500 93.510 114.880 109.810 ;
        RECT 115.200 93.190 115.580 110.130 ;
        RECT 115.900 93.510 116.280 109.810 ;
        RECT 116.600 93.190 116.980 110.130 ;
        RECT 117.300 93.510 117.680 109.810 ;
        RECT 118.000 93.190 118.380 110.130 ;
        RECT 118.700 93.510 119.080 109.810 ;
        RECT 119.400 93.190 119.780 110.130 ;
        RECT 120.100 93.510 120.480 109.810 ;
        RECT 120.800 93.190 121.180 110.130 ;
        RECT 121.500 93.510 121.880 109.810 ;
        RECT 122.200 93.190 122.580 110.130 ;
        RECT 122.900 93.510 123.280 109.810 ;
        RECT 123.600 93.190 123.980 110.130 ;
        RECT 124.300 93.510 124.680 109.810 ;
        RECT 125.000 93.190 125.380 110.130 ;
        RECT 125.700 93.510 126.080 109.810 ;
        RECT 126.400 93.190 126.780 110.130 ;
        RECT 127.100 93.510 127.480 109.810 ;
        RECT 127.800 93.190 128.180 110.130 ;
        RECT 83.000 92.730 128.180 93.190 ;
        RECT 83.000 75.790 83.380 92.730 ;
        RECT 83.700 76.110 84.080 92.410 ;
        RECT 84.400 75.790 84.780 92.730 ;
        RECT 85.100 76.110 85.480 92.410 ;
        RECT 85.800 75.790 86.180 92.730 ;
        RECT 86.500 76.110 86.880 92.410 ;
        RECT 87.200 75.790 87.580 92.730 ;
        RECT 87.900 76.110 88.280 92.410 ;
        RECT 88.600 75.790 88.980 92.730 ;
        RECT 89.300 76.110 89.680 92.410 ;
        RECT 90.000 75.790 90.380 92.730 ;
        RECT 90.700 76.110 91.080 92.410 ;
        RECT 91.400 75.790 91.780 92.730 ;
        RECT 92.100 76.110 92.480 92.410 ;
        RECT 92.800 75.790 93.180 92.730 ;
        RECT 93.500 76.110 93.880 92.410 ;
        RECT 94.200 75.790 94.580 92.730 ;
        RECT 94.900 76.110 95.280 92.410 ;
        RECT 95.600 75.790 95.980 92.730 ;
        RECT 96.300 76.110 96.680 92.410 ;
        RECT 97.000 75.790 97.380 92.730 ;
        RECT 97.700 76.110 98.080 92.410 ;
        RECT 98.400 75.790 98.780 92.730 ;
        RECT 99.100 76.110 99.480 92.410 ;
        RECT 99.800 75.790 100.180 92.730 ;
        RECT 100.500 76.110 100.880 92.410 ;
        RECT 101.200 75.790 101.580 92.730 ;
        RECT 101.900 76.110 102.280 92.410 ;
        RECT 102.600 75.790 102.980 92.730 ;
        RECT 103.300 76.110 103.680 92.410 ;
        RECT 104.000 75.790 104.380 92.730 ;
        RECT 104.700 76.110 105.080 92.410 ;
        RECT 105.400 75.790 105.780 92.730 ;
        RECT 106.100 76.110 106.480 92.410 ;
        RECT 106.800 75.790 107.180 92.730 ;
        RECT 107.500 76.110 107.880 92.410 ;
        RECT 108.200 75.790 108.580 92.730 ;
        RECT 108.900 76.110 109.280 92.410 ;
        RECT 109.600 75.790 109.980 92.730 ;
        RECT 110.300 76.110 110.680 92.410 ;
        RECT 111.000 75.790 111.380 92.730 ;
        RECT 111.700 76.110 112.080 92.410 ;
        RECT 112.400 75.790 112.780 92.730 ;
        RECT 113.100 76.110 113.480 92.410 ;
        RECT 113.800 75.790 114.180 92.730 ;
        RECT 114.500 76.110 114.880 92.410 ;
        RECT 115.200 75.790 115.580 92.730 ;
        RECT 115.900 76.110 116.280 92.410 ;
        RECT 116.600 75.790 116.980 92.730 ;
        RECT 117.300 76.110 117.680 92.410 ;
        RECT 118.000 75.790 118.380 92.730 ;
        RECT 118.700 76.110 119.080 92.410 ;
        RECT 119.400 75.790 119.780 92.730 ;
        RECT 120.100 76.110 120.480 92.410 ;
        RECT 120.800 75.790 121.180 92.730 ;
        RECT 121.500 76.110 121.880 92.410 ;
        RECT 122.200 75.790 122.580 92.730 ;
        RECT 122.900 76.110 123.280 92.410 ;
        RECT 123.600 75.790 123.980 92.730 ;
        RECT 124.300 76.110 124.680 92.410 ;
        RECT 125.000 75.790 125.380 92.730 ;
        RECT 125.700 76.110 126.080 92.410 ;
        RECT 126.400 75.790 126.780 92.730 ;
        RECT 127.100 76.110 127.480 92.410 ;
        RECT 127.800 75.790 128.180 92.730 ;
        RECT 83.000 75.330 128.180 75.790 ;
        RECT 83.000 58.390 83.380 75.330 ;
        RECT 83.700 58.710 84.080 75.010 ;
        RECT 84.400 58.390 84.780 75.330 ;
        RECT 85.100 58.710 85.480 75.010 ;
        RECT 85.800 58.390 86.180 75.330 ;
        RECT 86.500 58.710 86.880 75.010 ;
        RECT 87.200 58.390 87.580 75.330 ;
        RECT 87.900 58.710 88.280 75.010 ;
        RECT 88.600 58.390 88.980 75.330 ;
        RECT 89.300 58.710 89.680 75.010 ;
        RECT 90.000 58.390 90.380 75.330 ;
        RECT 90.700 58.710 91.080 75.010 ;
        RECT 91.400 58.390 91.780 75.330 ;
        RECT 92.100 58.710 92.480 75.010 ;
        RECT 92.800 58.390 93.180 75.330 ;
        RECT 93.500 58.710 93.880 75.010 ;
        RECT 94.200 58.390 94.580 75.330 ;
        RECT 94.900 58.710 95.280 75.010 ;
        RECT 95.600 58.390 95.980 75.330 ;
        RECT 96.300 58.710 96.680 75.010 ;
        RECT 97.000 58.390 97.380 75.330 ;
        RECT 97.700 58.710 98.080 75.010 ;
        RECT 98.400 58.390 98.780 75.330 ;
        RECT 99.100 58.710 99.480 75.010 ;
        RECT 99.800 58.390 100.180 75.330 ;
        RECT 100.500 58.710 100.880 75.010 ;
        RECT 101.200 58.390 101.580 75.330 ;
        RECT 101.900 58.710 102.280 75.010 ;
        RECT 102.600 58.390 102.980 75.330 ;
        RECT 103.300 58.710 103.680 75.010 ;
        RECT 104.000 58.390 104.380 75.330 ;
        RECT 104.700 58.710 105.080 75.010 ;
        RECT 105.400 58.390 105.780 75.330 ;
        RECT 106.100 58.710 106.480 75.010 ;
        RECT 106.800 58.390 107.180 75.330 ;
        RECT 107.500 58.710 107.880 75.010 ;
        RECT 108.200 58.390 108.580 75.330 ;
        RECT 108.900 58.710 109.280 75.010 ;
        RECT 109.600 58.390 109.980 75.330 ;
        RECT 110.300 58.710 110.680 75.010 ;
        RECT 111.000 58.390 111.380 75.330 ;
        RECT 111.700 58.710 112.080 75.010 ;
        RECT 112.400 58.390 112.780 75.330 ;
        RECT 113.100 58.710 113.480 75.010 ;
        RECT 113.800 58.390 114.180 75.330 ;
        RECT 114.500 58.710 114.880 75.010 ;
        RECT 115.200 58.390 115.580 75.330 ;
        RECT 115.900 58.710 116.280 75.010 ;
        RECT 116.600 58.390 116.980 75.330 ;
        RECT 117.300 58.710 117.680 75.010 ;
        RECT 118.000 58.390 118.380 75.330 ;
        RECT 118.700 58.710 119.080 75.010 ;
        RECT 119.400 58.390 119.780 75.330 ;
        RECT 120.100 58.710 120.480 75.010 ;
        RECT 120.800 58.390 121.180 75.330 ;
        RECT 121.500 58.710 121.880 75.010 ;
        RECT 122.200 58.390 122.580 75.330 ;
        RECT 122.900 58.710 123.280 75.010 ;
        RECT 123.600 58.390 123.980 75.330 ;
        RECT 124.300 58.710 124.680 75.010 ;
        RECT 125.000 58.390 125.380 75.330 ;
        RECT 125.700 58.710 126.080 75.010 ;
        RECT 126.400 58.390 126.780 75.330 ;
        RECT 127.100 58.710 127.480 75.010 ;
        RECT 127.800 58.390 128.180 75.330 ;
        RECT 83.000 57.930 128.180 58.390 ;
        RECT 83.000 40.990 83.380 57.930 ;
        RECT 83.700 41.310 84.080 57.610 ;
        RECT 84.400 40.990 84.780 57.930 ;
        RECT 85.100 41.310 85.480 57.610 ;
        RECT 85.800 40.990 86.180 57.930 ;
        RECT 86.500 41.310 86.880 57.610 ;
        RECT 87.200 40.990 87.580 57.930 ;
        RECT 87.900 41.310 88.280 57.610 ;
        RECT 88.600 40.990 88.980 57.930 ;
        RECT 89.300 41.310 89.680 57.610 ;
        RECT 90.000 40.990 90.380 57.930 ;
        RECT 90.700 41.310 91.080 57.610 ;
        RECT 91.400 40.990 91.780 57.930 ;
        RECT 92.100 41.310 92.480 57.610 ;
        RECT 92.800 40.990 93.180 57.930 ;
        RECT 93.500 41.310 93.880 57.610 ;
        RECT 94.200 40.990 94.580 57.930 ;
        RECT 94.900 41.310 95.280 57.610 ;
        RECT 95.600 40.990 95.980 57.930 ;
        RECT 96.300 41.310 96.680 57.610 ;
        RECT 97.000 40.990 97.380 57.930 ;
        RECT 97.700 41.310 98.080 57.610 ;
        RECT 98.400 40.990 98.780 57.930 ;
        RECT 99.100 41.310 99.480 57.610 ;
        RECT 99.800 40.990 100.180 57.930 ;
        RECT 100.500 41.310 100.880 57.610 ;
        RECT 101.200 40.990 101.580 57.930 ;
        RECT 101.900 41.310 102.280 57.610 ;
        RECT 102.600 40.990 102.980 57.930 ;
        RECT 103.300 41.310 103.680 57.610 ;
        RECT 104.000 40.990 104.380 57.930 ;
        RECT 104.700 41.310 105.080 57.610 ;
        RECT 105.400 40.990 105.780 57.930 ;
        RECT 106.100 41.310 106.480 57.610 ;
        RECT 106.800 40.990 107.180 57.930 ;
        RECT 107.500 41.310 107.880 57.610 ;
        RECT 108.200 40.990 108.580 57.930 ;
        RECT 108.900 41.310 109.280 57.610 ;
        RECT 109.600 40.990 109.980 57.930 ;
        RECT 110.300 41.310 110.680 57.610 ;
        RECT 111.000 40.990 111.380 57.930 ;
        RECT 111.700 41.310 112.080 57.610 ;
        RECT 112.400 40.990 112.780 57.930 ;
        RECT 113.100 41.310 113.480 57.610 ;
        RECT 113.800 40.990 114.180 57.930 ;
        RECT 114.500 41.310 114.880 57.610 ;
        RECT 115.200 40.990 115.580 57.930 ;
        RECT 115.900 41.310 116.280 57.610 ;
        RECT 116.600 40.990 116.980 57.930 ;
        RECT 117.300 41.310 117.680 57.610 ;
        RECT 118.000 40.990 118.380 57.930 ;
        RECT 118.700 41.310 119.080 57.610 ;
        RECT 119.400 40.990 119.780 57.930 ;
        RECT 120.100 41.310 120.480 57.610 ;
        RECT 120.800 40.990 121.180 57.930 ;
        RECT 121.500 41.310 121.880 57.610 ;
        RECT 122.200 40.990 122.580 57.930 ;
        RECT 122.900 41.310 123.280 57.610 ;
        RECT 123.600 40.990 123.980 57.930 ;
        RECT 124.300 41.310 124.680 57.610 ;
        RECT 125.000 40.990 125.380 57.930 ;
        RECT 125.700 41.310 126.080 57.610 ;
        RECT 126.400 40.990 126.780 57.930 ;
        RECT 127.100 41.310 127.480 57.610 ;
        RECT 127.800 40.990 128.180 57.930 ;
        RECT 12.940 40.610 65.440 40.990 ;
        RECT 13.600 38.920 49.240 38.980 ;
        RECT 13.600 38.540 49.980 38.920 ;
        RECT 13.600 37.660 48.520 38.100 ;
        RECT 13.600 36.340 13.960 37.660 ;
        RECT 48.880 37.220 49.240 38.540 ;
        RECT 14.320 36.780 49.240 37.220 ;
        RECT 13.600 35.900 47.800 36.340 ;
        RECT 48.160 35.900 48.520 36.340 ;
        RECT 13.600 34.580 13.960 35.900 ;
        RECT 48.880 35.460 49.240 36.780 ;
        RECT 14.320 35.020 15.040 35.460 ;
        RECT 15.400 35.020 49.240 35.460 ;
        RECT 13.600 34.520 49.240 34.580 ;
        RECT 12.860 34.140 49.240 34.520 ;
        RECT 12.860 29.240 13.240 34.140 ;
        RECT 13.600 33.640 49.240 33.700 ;
        RECT 49.600 33.640 49.980 38.540 ;
        RECT 13.600 33.260 49.980 33.640 ;
        RECT 13.600 32.380 48.520 32.820 ;
        RECT 13.600 31.060 13.960 32.380 ;
        RECT 48.880 31.940 49.240 33.260 ;
        RECT 14.320 31.500 49.240 31.940 ;
        RECT 13.600 30.620 47.800 31.060 ;
        RECT 48.160 30.620 48.520 31.060 ;
        RECT 13.600 29.300 13.960 30.620 ;
        RECT 48.880 30.180 49.240 31.500 ;
        RECT 14.320 29.740 15.040 30.180 ;
        RECT 15.400 29.740 49.240 30.180 ;
        RECT 13.600 29.240 49.240 29.300 ;
        RECT 12.860 28.860 49.240 29.240 ;
        RECT 12.860 23.960 13.240 28.860 ;
        RECT 13.600 28.360 49.240 28.420 ;
        RECT 49.600 28.360 49.980 33.260 ;
        RECT 13.600 27.980 49.980 28.360 ;
        RECT 13.600 27.100 48.520 27.540 ;
        RECT 13.600 25.780 13.960 27.100 ;
        RECT 48.880 26.660 49.240 27.980 ;
        RECT 14.320 26.220 49.240 26.660 ;
        RECT 13.600 25.340 47.800 25.780 ;
        RECT 48.160 25.340 48.520 25.780 ;
        RECT 13.600 24.020 13.960 25.340 ;
        RECT 48.880 24.900 49.240 26.220 ;
        RECT 14.320 24.460 15.040 24.900 ;
        RECT 15.400 24.460 49.240 24.900 ;
        RECT 13.600 23.960 49.240 24.020 ;
        RECT 12.860 23.580 49.240 23.960 ;
        RECT 49.600 23.590 49.980 27.980 ;
        RECT 12.860 18.680 13.240 23.580 ;
        RECT 49.600 23.210 53.560 23.590 ;
        RECT 13.600 23.080 49.240 23.140 ;
        RECT 49.600 23.080 49.980 23.210 ;
        RECT 13.600 22.700 49.980 23.080 ;
        RECT 13.600 21.820 48.520 22.260 ;
        RECT 13.600 20.500 13.960 21.820 ;
        RECT 48.880 21.380 49.240 22.700 ;
        RECT 14.320 20.940 49.240 21.380 ;
        RECT 13.600 20.060 47.800 20.500 ;
        RECT 48.160 20.060 48.520 20.500 ;
        RECT 13.600 18.740 13.960 20.060 ;
        RECT 48.880 19.620 49.240 20.940 ;
        RECT 14.320 19.180 15.040 19.620 ;
        RECT 15.400 19.180 49.240 19.620 ;
        RECT 13.600 18.680 49.240 18.740 ;
        RECT 12.860 18.300 49.240 18.680 ;
        RECT 12.860 13.400 13.240 18.300 ;
        RECT 13.600 17.800 49.240 17.860 ;
        RECT 49.600 17.800 49.980 22.700 ;
        RECT 52.560 19.250 54.280 19.630 ;
        RECT 53.900 19.190 54.280 19.250 ;
        RECT 54.720 19.190 55.720 39.640 ;
        RECT 53.900 18.810 55.720 19.190 ;
        RECT 13.600 17.420 49.980 17.800 ;
        RECT 13.600 16.540 48.520 16.980 ;
        RECT 13.600 15.220 13.960 16.540 ;
        RECT 48.880 16.100 49.240 17.420 ;
        RECT 14.320 15.660 49.240 16.100 ;
        RECT 13.600 14.780 47.800 15.220 ;
        RECT 48.160 14.780 48.520 15.220 ;
        RECT 13.600 13.460 13.960 14.780 ;
        RECT 48.880 14.340 49.240 15.660 ;
        RECT 14.320 13.900 15.040 14.340 ;
        RECT 15.400 13.900 49.240 14.340 ;
        RECT 13.600 13.400 49.240 13.460 ;
        RECT 12.860 13.020 49.240 13.400 ;
        RECT 54.720 6.040 55.720 18.810 ;
        RECT 58.680 9.640 59.680 39.640 ;
        RECT 61.600 30.210 62.600 30.590 ;
        RECT 61.910 4.380 62.290 30.210 ;
        RECT 65.060 19.190 65.440 40.610 ;
        RECT 75.880 40.610 128.180 40.990 ;
        RECT 128.500 40.610 128.880 110.510 ;
        RECT 67.240 25.850 75.440 26.230 ;
        RECT 67.240 19.190 67.620 25.850 ;
        RECT 75.880 19.190 76.260 40.610 ;
        RECT 78.720 30.210 79.720 30.590 ;
        RECT 65.060 18.810 67.620 19.190 ;
        RECT 74.440 18.810 76.260 19.190 ;
        RECT 65.800 14.370 66.800 14.750 ;
        RECT 74.520 14.370 75.520 14.750 ;
        RECT 79.030 4.380 79.410 30.210 ;
        RECT 81.640 9.640 82.640 39.640 ;
        RECT 85.600 19.190 86.600 39.640 ;
        RECT 92.080 38.920 127.720 38.980 ;
        RECT 91.340 38.540 127.720 38.920 ;
        RECT 91.340 33.640 91.720 38.540 ;
        RECT 92.080 37.220 92.440 38.540 ;
        RECT 92.800 37.660 127.720 38.100 ;
        RECT 92.080 36.780 127.000 37.220 ;
        RECT 92.080 35.460 92.440 36.780 ;
        RECT 127.360 36.340 127.720 37.660 ;
        RECT 92.800 35.900 93.160 36.340 ;
        RECT 93.520 35.900 127.720 36.340 ;
        RECT 92.080 35.020 125.920 35.460 ;
        RECT 126.280 35.020 127.000 35.460 ;
        RECT 127.360 34.580 127.720 35.900 ;
        RECT 92.080 34.520 127.720 34.580 ;
        RECT 92.080 34.140 128.460 34.520 ;
        RECT 92.080 33.640 127.720 33.700 ;
        RECT 91.340 33.260 127.720 33.640 ;
        RECT 91.340 28.360 91.720 33.260 ;
        RECT 92.080 31.940 92.440 33.260 ;
        RECT 92.800 32.380 127.720 32.820 ;
        RECT 92.080 31.500 127.000 31.940 ;
        RECT 92.080 30.180 92.440 31.500 ;
        RECT 127.360 31.060 127.720 32.380 ;
        RECT 92.800 30.620 93.160 31.060 ;
        RECT 93.520 30.620 127.720 31.060 ;
        RECT 92.080 29.740 125.920 30.180 ;
        RECT 126.280 29.740 127.000 30.180 ;
        RECT 127.360 29.300 127.720 30.620 ;
        RECT 92.080 29.240 127.720 29.300 ;
        RECT 128.080 29.240 128.460 34.140 ;
        RECT 92.080 28.860 128.460 29.240 ;
        RECT 92.080 28.360 127.720 28.420 ;
        RECT 91.340 27.980 127.720 28.360 ;
        RECT 91.340 23.590 91.720 27.980 ;
        RECT 92.080 26.660 92.440 27.980 ;
        RECT 92.800 27.100 127.720 27.540 ;
        RECT 92.080 26.220 127.000 26.660 ;
        RECT 92.080 24.900 92.440 26.220 ;
        RECT 127.360 25.780 127.720 27.100 ;
        RECT 92.800 25.340 93.160 25.780 ;
        RECT 93.520 25.340 127.720 25.780 ;
        RECT 92.080 24.460 125.920 24.900 ;
        RECT 126.280 24.460 127.000 24.900 ;
        RECT 127.360 24.020 127.720 25.340 ;
        RECT 87.760 23.210 91.720 23.590 ;
        RECT 92.080 23.960 127.720 24.020 ;
        RECT 128.080 23.960 128.460 28.860 ;
        RECT 92.080 23.580 128.460 23.960 ;
        RECT 91.340 23.080 91.720 23.210 ;
        RECT 92.080 23.080 127.720 23.140 ;
        RECT 91.340 22.700 127.720 23.080 ;
        RECT 87.040 19.250 88.760 19.630 ;
        RECT 87.040 19.190 87.420 19.250 ;
        RECT 85.600 18.810 87.420 19.190 ;
        RECT 85.600 6.040 86.600 18.810 ;
        RECT 91.340 17.800 91.720 22.700 ;
        RECT 92.080 21.380 92.440 22.700 ;
        RECT 92.800 21.820 127.720 22.260 ;
        RECT 92.080 20.940 127.000 21.380 ;
        RECT 92.080 19.620 92.440 20.940 ;
        RECT 127.360 20.500 127.720 21.820 ;
        RECT 92.800 20.060 93.160 20.500 ;
        RECT 93.520 20.060 127.720 20.500 ;
        RECT 92.080 19.180 125.920 19.620 ;
        RECT 126.280 19.180 127.000 19.620 ;
        RECT 127.360 18.740 127.720 20.060 ;
        RECT 92.080 18.680 127.720 18.740 ;
        RECT 128.080 18.680 128.460 23.580 ;
        RECT 92.080 18.300 128.460 18.680 ;
        RECT 92.080 17.800 127.720 17.860 ;
        RECT 91.340 17.420 127.720 17.800 ;
        RECT 92.080 16.100 92.440 17.420 ;
        RECT 92.800 16.540 127.720 16.980 ;
        RECT 92.080 15.660 127.000 16.100 ;
        RECT 92.080 14.340 92.440 15.660 ;
        RECT 127.360 15.220 127.720 16.540 ;
        RECT 92.800 14.780 93.160 15.220 ;
        RECT 93.520 14.780 127.720 15.220 ;
        RECT 92.080 13.900 125.920 14.340 ;
        RECT 126.280 13.900 127.000 14.340 ;
        RECT 127.360 13.460 127.720 14.780 ;
        RECT 92.080 13.400 127.720 13.460 ;
        RECT 128.080 13.400 128.460 18.300 ;
        RECT 92.080 13.020 128.460 13.400 ;
        RECT 61.600 4.000 62.600 4.380 ;
        RECT 78.720 4.000 79.720 4.380 ;
        RECT 143.680 2.660 144.680 222.660 ;
        RECT 147.640 2.660 148.640 222.660 ;
  END
END tt_um_TT06_SAR_wulffern
END LIBRARY

