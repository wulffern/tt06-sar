* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130B

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
*+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
*+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7]
*+ uo_out[6] ui_in[0] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=240.246 ps=1.2657k w=1.08 l=0.18
R2 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=244.0044 ps=1.27698k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA3.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X49 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X50 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X51 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X52 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X56 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X58 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X63 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X65 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X66 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X67 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X72 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X74 SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X76 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X77 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X78 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X79 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_SAR8B_CV_0.XA6.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X88 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X90 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X95 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X96 ua[1] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X97 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X98 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X99 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X100 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X101 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X106 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X107 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R8 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X108 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R9 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X114 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X115 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X116 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 VGND SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X118 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X119 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X120 SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X121 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X122 SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X124 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X125 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X130 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X131 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X132 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X134 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X135 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X136 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X137 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X146 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X147 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X148 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X149 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X150 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X155 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X158 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X160 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X163 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA4.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X166 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X167 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X169 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X174 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X175 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R13 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X176 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X177 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X178 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X181 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X185 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X186 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X188 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y SUNSAR_CAPT8B_CV_0.XA3.A SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X193 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X194 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X195 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X198 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R14 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X199 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X201 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R15 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X205 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X206 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X207 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 VGND SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X212 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X213 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X214 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X216 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R16 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X221 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X223 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X225 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X228 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X229 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X230 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X232 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X233 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X235 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X236 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X237 SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X239 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X244 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X246 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X253 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X255 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X263 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X266 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X267 ua[0] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X268 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X270 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X275 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R17 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X276 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R18 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X278 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X280 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA5.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R19 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X282 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X284 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X286 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X288 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X292 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X294 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X295 SUNSAR_CAPT8B_CV_0.XA5.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X300 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X307 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X308 VPWR SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA1.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R20 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X309 VGND SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X310 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X311 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X312 SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X313 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X314 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X316 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X318 SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X321 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X322 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XB2.XA3.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X324 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X328 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X333 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R23 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X337 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X338 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X341 ua[1] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X342 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X344 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X346 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X347 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X348 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X349 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X351 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X352 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X359 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X360 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X364 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X365 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X366 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R24 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X368 SUNSAR_SAR8B_CV_0.XA3.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X370 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X371 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X372 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X373 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X374 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X375 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X376 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X377 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X378 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X379 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X381 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X382 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X384 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X385 SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X386 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X387 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R25 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X388 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X389 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X390 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X391 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X393 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X394 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X395 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X400 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X402 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R26 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X404 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R27 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X407 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X410 SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X413 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X414 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 SUNSAR_CAPT8B_CV_0.XA3.A ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X416 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X417 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X418 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X419 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X420 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X421 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X422 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X423 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X424 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X425 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X426 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X427 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X428 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X429 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X433 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X434 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X435 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X436 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X437 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R29 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X440 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X441 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X442 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X443 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R30 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X447 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X449 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X450 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X452 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X453 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X454 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X455 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X457 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R31 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X458 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X459 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X462 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X463 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X465 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X468 SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R32 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X470 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X471 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X472 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X473 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X474 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X477 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X478 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X479 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X480 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X481 VGND SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X482 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X484 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X486 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X489 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X491 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X492 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X493 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X494 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X496 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R34 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X498 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X499 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X500 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X501 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X502 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R35 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X503 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X505 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X506 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X508 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X510 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X511 SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X512 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X513 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X514 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X515 SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X516 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X517 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X519 ua[0] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X520 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X521 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X522 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X525 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X526 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X527 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X528 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X530 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X532 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X533 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R36 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X536 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X537 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X540 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X541 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X544 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X545 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X548 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 ua[1] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X553 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X554 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X557 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X558 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X560 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X561 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X562 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X564 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X565 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X567 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X568 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X570 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X571 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X572 ua[1] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X573 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S SUNSAR_CAPT8B_CV_0.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X574 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X575 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X578 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X579 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X580 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X581 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X582 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X583 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X584 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R37 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X585 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X587 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X588 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X589 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X590 SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R38 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X591 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X592 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X593 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X594 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X595 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X596 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X598 VGND SUNSAR_CAPT8B_CV_0.XA3.A SUNSAR_CAPT8B_CV_0.XA5.XA1.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X600 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X601 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X602 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X603 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X604 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X605 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X606 SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X607 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X609 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X610 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X612 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X613 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X614 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X615 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X616 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X618 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X619 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X620 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X621 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X624 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X626 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X629 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X631 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X634 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X635 SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X636 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X637 SUNSAR_SAR8B_CV_0.XA7.XA6.MP0.D SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X638 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X639 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X640 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R40 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X641 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X642 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R41 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X643 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X644 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X645 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X646 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X647 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R42 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X648 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X649 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X650 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X652 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X653 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X654 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R43 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R44 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X656 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X657 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X658 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X661 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X663 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X664 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X665 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X666 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X667 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X668 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X669 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X670 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X674 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X675 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X676 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y SUNSAR_CAPT8B_CV_0.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X678 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R45 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X680 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X681 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X682 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X683 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X684 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA3.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R46 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X685 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X686 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X687 SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X688 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 SUNSAR_CAPT8B_CV_0.XA5.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X690 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X691 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X693 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X694 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X695 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X696 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X697 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X698 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X699 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X700 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X701 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X703 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X704 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X705 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X706 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X707 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X709 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X710 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 ua[0] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X713 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R48 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X714 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X715 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X716 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X717 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X718 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X719 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X720 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X721 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X722 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X725 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X726 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X727 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X728 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X729 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X730 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X731 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X732 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X733 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X734 ua[0] SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X735 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X737 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R49 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X738 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X740 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X741 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X742 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 SUNSAR_SAR8B_CV_0.XA2.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X745 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X746 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X747 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X749 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X751 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X752 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X753 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X754 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X755 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R51 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X757 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X759 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X760 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X761 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X762 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X763 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X764 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X765 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X766 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X767 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X768 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X770 VGND SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X771 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X773 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X774 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R53 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X775 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X776 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X777 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X778 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X779 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X780 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X782 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X783 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X786 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X787 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X788 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X790 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X791 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X792 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X793 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X794 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X798 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X800 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XA3.A ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X802 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X808 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X809 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X810 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X813 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X814 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X816 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X817 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X818 SUNSAR_SAR8B_CV_0.XA0.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X819 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X820 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X821 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X822 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X823 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X824 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X825 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X828 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R54 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X829 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X830 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X831 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X832 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X833 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R55 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X834 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X835 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X836 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X837 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X838 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X839 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X840 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X842 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X843 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X844 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X845 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X847 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X848 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X849 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X850 SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X852 SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X853 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X854 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X855 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X857 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X858 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X859 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X862 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X863 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X864 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X865 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X866 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X867 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X868 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X869 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X871 VGND SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X872 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X873 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X874 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X875 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X876 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X878 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R57 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X879 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X883 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X884 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X885 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X886 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R58 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X887 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VGND SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X890 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X892 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X893 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X894 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X895 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X896 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X897 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X898 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X899 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R60 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X901 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X902 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X903 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R61 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X905 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X906 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X908 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X909 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X910 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X911 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X912 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X913 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X914 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X915 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X917 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X918 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X920 SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X923 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X924 SUNSAR_SAR8B_CV_0.XA1.XA6.MP0.D SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X925 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X926 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X928 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X929 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X930 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R62 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X931 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X932 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X933 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X934 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X935 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X936 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X937 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X939 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X940 SUNSAR_SAR8B_CV_0.XB1.XA3.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X941 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X942 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X944 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R63 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X945 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X946 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X947 VGND SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X948 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X949 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X950 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X951 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X953 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X954 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X955 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X957 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X959 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X961 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y SUNSAR_CAPT8B_CV_0.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X962 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X963 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X964 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X965 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X967 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X968 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X970 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X971 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X972 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X974 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X975 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X976 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X978 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X980 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X981 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X982 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X984 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X985 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X986 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X987 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X988 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R65 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R66 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X989 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X993 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X994 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X995 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R67 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X997 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X999 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1000 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1001 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1002 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1003 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1004 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1005 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1008 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1010 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1013 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1014 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1015 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1016 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1018 SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1019 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1020 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1021 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1022 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1025 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1028 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 VGND SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1033 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1034 SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1035 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR 0.916737f
C1 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR 2.52813f
C2 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.611221f
C3 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR 0.877293f
C4 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S 0.142644f
C5 a_13842_36828# VPWR 0.392558f
C6 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.868329f
C7 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.4301f
C8 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.CKN 0.190344f
C9 SUNSAR_CAPT8B_CV_0.XA3.Y VPWR 0.845896f
C10 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_12710_42408# 0.111909f
C11 SUNSAR_SAR8B_CV_0.XA1.ENO VPWR 4.43046f
C12 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VPWR 0.263064f
C13 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO 0.144331f
C14 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.401945f
C15 a_8802_26796# VPWR 0.441293f
C16 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C17 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.885278f
C18 SUNSAR_SAR8B_CV_0.D<3> VPWR 4.54507f
C19 a_23922_35948# VPWR 0.388238f
C20 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR 2.52823f
C21 SUNSAR_SAR8B_CV_0.EN a_15210_29612# 0.143511f
C22 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.133602f
C23 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR 0.877293f
C24 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.180155f
C25 SUNSAR_SAR8B_CV_0.SARN VPWR 0.130754f
C26 a_23942_43640# VPWR 0.410001f
C27 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.290432f
C28 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y a_8822_41000# 0.15757f
C29 SUNSAR_SAR8B_CV_0.XA0.ENO VPWR 5.00453f
C30 a_10190_44168# VPWR 0.338694f
C31 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.965002f
C32 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.275206f
C33 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.78158f
C34 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.51035f
C35 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA8.A 0.527529f
C36 SUNSAR_SAR8B_CV_0.EN a_13842_29612# 0.143511f
C37 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARN 0.639272f
C38 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.Y 0.649845f
C39 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.183479f
C40 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.117496f
C41 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR 0.877293f
C42 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S 0.142624f
C43 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.27418f
C44 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.233892f
C45 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y uo_out[1] 0.305934f
C46 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.146492f
C47 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y a_7670_41000# 0.114097f
C48 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_11342_42408# 0.113479f
C49 a_5150_40296# VPWR 0.452721f
C50 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.1913f
C51 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.885118f
C52 a_8822_44168# VPWR 0.339109f
C53 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y a_8822_42760# 0.113305f
C54 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D 0.150367f
C55 a_20250_32076# VPWR 0.42896f
C56 a_20250_28204# VPWR 0.360102f
C57 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.137745f
C58 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.Y 0.744161f
C59 SUNSAR_SAR8B_CV_0.XA20.XA2.CO a_23922_30844# 0.100515f
C60 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.133602f
C61 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR 0.877293f
C62 a_10170_36828# VPWR 0.392843f
C63 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.105092f
C64 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.29345f
C65 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.ENO 1.22625f
C66 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y uo_out[1] 0.248851f
C67 a_3782_40296# VPWR 0.454411f
C68 a_20250_35068# VPWR 0.388548f
C69 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.ENO 0.497337f
C70 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARN 0.487857f
C71 a_5130_26796# VPWR 0.440138f
C72 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y a_17750_42408# 0.100131f
C73 SUNSAR_SAR8B_CV_0.XA5.XA2.A a_15210_30316# 0.127528f
C74 SUNSAR_SAR8B_CV_0.D<4> VPWR 4.52288f
C75 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.474658f
C76 a_20250_35948# VPWR 0.411511f
C77 a_18882_32076# VPWR 0.430937f
C78 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.412143f
C79 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 0.611321f
C80 a_18882_28204# VPWR 0.360178f
C81 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.05725f
C82 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR 0.877293f
C83 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S 0.142644f
C84 a_8802_36828# VPWR 0.392894f
C85 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR 0.394875f
C86 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.136948f
C87 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.22339f
C88 a_9990_3334# VPWR 0.377065f
C89 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR 0.100103f
C90 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.152047f
C91 a_18882_35068# VPWR 0.391042f
C92 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA10.Y 0.303978f
C93 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.51035f
C94 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.321724f
C95 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35068# 0.127528f
C96 a_3762_26796# VPWR 0.441293f
C97 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.779324f
C98 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C99 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D 0.146505f
C100 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR 0.100103f
C101 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.329693f
C102 a_18882_35948# VPWR 0.414005f
C103 SUNSAR_SAR8B_CV_0.EN a_10170_29612# 0.143511f
C104 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR 0.877293f
C105 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.133602f
C106 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR 1.65869f
C107 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.132806f
C108 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.132601f
C109 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.318734f
C110 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.412248f
C111 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR 2.89798f
C112 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.339883f
C113 a_23942_40648# VPWR 0.486201f
C114 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.13078f
C115 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO 0.144331f
C116 a_5150_44168# VPWR 0.338694f
C117 SUNSAR_SAR8B_CV_0.XA4.XA2.A a_13842_30316# 0.129098f
C118 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR 0.100103f
C119 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.51035f
C120 SUNSAR_SAR8B_CV_0.EN a_8802_29612# 0.143511f
C121 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR 0.877293f
C122 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S 0.142624f
C123 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.121229f
C124 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.513782f
C125 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C126 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.132886f
C127 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.63636f
C128 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.124212f
C129 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VPWR 1.74634f
C130 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.720184f
C131 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y a_6302_41000# 0.115667f
C132 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.D<0> 0.362609f
C133 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_7670_42408# 0.111909f
C134 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.84356f
C135 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C136 a_23922_27148# VPWR 0.480439f
C137 a_3782_44168# VPWR 0.339109f
C138 SUNSAR_SAR8B_CV_0.D<5> VPWR 4.53355f
C139 a_15210_32076# VPWR 0.430937f
C140 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA8.A 0.527529f
C141 a_15210_28204# VPWR 0.360102f
C142 a_23942_42760# VPWR 0.3859f
C143 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.133602f
C144 a_5130_36828# VPWR 0.392615f
C145 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.132806f
C146 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.ENO 1.22625f
C147 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.412248f
C148 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR 1.42562f
C149 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y uo_out[2] 0.246827f
C150 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR 0.100103f
C151 SUNSAR_CAPT8B_CV_0.XA5.A a_22790_41880# 0.107417f
C152 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y a_5150_41000# 0.156079f
C153 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_SAR8B_CV_0.D<0> 0.238616f
C154 a_15210_35068# VPWR 0.391042f
C155 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.331639f
C156 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.ENO 0.431783f
C157 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VPWR 0.263064f
C158 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA5.XA1.Y 0.134182f
C159 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.93403f
C160 a_15210_35948# VPWR 0.414005f
C161 a_13842_32076# VPWR 0.430937f
C162 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.205884f
C163 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.611221f
C164 a_13842_28204# VPWR 0.360178f
C165 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S 0.142644f
C166 a_3762_36828# VPWR 0.392706f
C167 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR 4.25329f
C168 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.132886f
C169 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR 0.175406f
C170 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y uo_out[2] 0.305131f
C171 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.154155f
C172 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.718754f
C173 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_6302_42408# 0.113479f
C174 a_20270_40648# VPWR 0.489593f
C175 a_13842_35068# VPWR 0.391042f
C176 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.111519f
C177 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 54.1913f
C178 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO 0.144331f
C179 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C180 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.779346f
C181 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y a_5150_42760# 0.111734f
C182 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D 0.150367f
C183 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.27006f
C184 a_13842_35948# VPWR 0.414005f
C185 SUNSAR_SAR8B_CV_0.EN a_5130_29612# 0.143511f
C186 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.Y 0.744161f
C187 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.133602f
C188 a_23922_34540# VPWR 0.499758f
C189 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.132806f
C190 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.CKN 0.152587f
C191 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.318734f
C192 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_2768# 0.172147f
C193 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR 1.42654f
C194 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.3401f
C195 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VPWR 1.74633f
C196 a_18902_40648# VPWR 0.488227f
C197 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.141203f
C198 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35068# 0.129098f
C199 a_20250_27148# VPWR 0.468331f
C200 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.282334f
C201 SUNSAR_SAR8B_CV_0.XA3.XA2.A a_10170_30316# 0.127528f
C202 SUNSAR_SAR8B_CV_0.D<6> VPWR 4.55788f
C203 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.1913f
C204 SUNSAR_SAR8B_CV_0.EN a_3762_29612# 0.143511f
C205 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.Y 0.649845f
C206 a_20270_42760# VPWR 0.388849f
C207 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.00437f
C208 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR 0.702312f
C209 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.100251f
C210 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.173526f
C211 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C212 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR 0.175406f
C213 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR 2.89805f
C214 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.718746f
C215 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1383f
C216 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.169736f
C217 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VPWR 0.263064f
C218 a_18882_27148# VPWR 0.468818f
C219 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.206053f
C220 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.188275f
C221 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.204048f
C222 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR 0.100103f
C223 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D 0.146505f
C224 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202696f
C225 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233285f
C226 a_10170_32076# VPWR 0.430937f
C227 a_10170_28204# VPWR 0.360102f
C228 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_34540# 0.103065f
C229 a_18902_42760# VPWR 0.388849f
C230 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.133602f
C231 SUNSAR_SAR8B_CV_0.XA7.CEO VPWR 1.08687f
C232 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.ENO 1.22625f
C233 a_16542_4038# VPWR 0.377115f
C234 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO 1.43919f
C235 a_10170_35068# VPWR 0.391042f
C236 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.ENO 0.497337f
C237 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.143714f
C238 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.199718f
C239 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR 0.100103f
C240 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.275206f
C241 SUNSAR_SAR8B_CV_0.XA2.XA2.A a_8802_30316# 0.129098f
C242 a_10170_35948# VPWR 0.414005f
C243 a_8802_32076# VPWR 0.430937f
C244 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 0.611321f
C245 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.205884f
C246 a_8802_28204# VPWR 0.360178f
C247 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.424961f
C248 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR 0.709784f
C249 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.03892f
C250 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C251 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.124212f
C252 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y uo_out[3] 0.309255f
C253 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR 0.100103f
C254 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.718754f
C255 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_2630_42408# 0.111909f
C256 a_15230_40648# VPWR 0.489593f
C257 a_8802_35068# VPWR 0.391042f
C258 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA10.Y 0.303978f
C259 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 6.84356f
C260 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y a_3782_42760# 0.113305f
C261 SUNSAR_SAR8B_CV_0.D<7> VPWR 3.46417f
C262 a_8802_35948# VPWR 0.414005f
C263 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.109554f
C264 SUNSAR_SAR8B_CV_0.XA6.CEO VPWR 2.14133f
C265 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.160605f
C266 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_3728# 0.172147f
C267 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.440597f
C268 SUNSAR_SAR8B_CV_0.XB2.XA4.GN ua[0] 0.63933f
C269 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y uo_out[3] 0.249748f
C270 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR 2.89805f
C271 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y a_3782_41000# 0.15757f
C272 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_SAR8B_CV_0.D<1> 0.238616f
C273 SUNSAR_SAR8B_CV_0.DONE ui_in[0] 0.167919f
C274 a_13862_40648# VPWR 0.488227f
C275 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.13078f
C276 SUNSAR_SAR8B_CV_0.XA7.XA11.Y a_21402_36828# 0.104051f
C277 a_15210_27148# VPWR 0.468331f
C278 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.12241f
C279 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.126354f
C280 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.SARP 0.12276f
C281 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.01993f
C282 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.84356f
C283 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.170798f
C284 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 2.95957f
C285 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.424961f
C286 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.SARP 0.131335f
C287 a_15230_42760# VPWR 0.388849f
C288 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR 0.706981f
C289 SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.D VPWR 0.105276f
C290 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G 0.22339f
C291 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.CKN 0.152587f
C292 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VPWR 1.74633f
C293 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.718746f
C294 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y a_2630_41000# 0.114097f
C295 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.D<1> 0.362008f
C296 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6267f
C297 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35068# 0.127528f
C298 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.142931f
C299 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.424961f
C300 a_13842_27148# VPWR 0.468818f
C301 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN 0.253395f
C302 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.432466f
C303 a_23942_41880# VPWR 0.395951f
C304 a_5130_32076# VPWR 0.430937f
C305 a_5130_28204# VPWR 0.360102f
C306 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.115348f
C307 a_13862_42760# VPWR 0.388849f
C308 SUNSAR_SAR8B_CV_0.XA5.CEO VPWR 1.02322f
C309 SUNSAR_SAR8B_CV_0.XA6.XA6.MP2.D VPWR 0.105892f
C310 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.109479f
C311 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.318734f
C312 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.440597f
C313 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR 0.100103f
C314 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C315 a_5130_35068# VPWR 0.391042f
C316 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.331639f
C317 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.ENO 0.428606f
C318 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C319 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y a_12710_42408# 0.100131f
C320 SUNSAR_SAR8B_CV_0.XA1.XA2.A a_5130_30316# 0.127528f
C321 a_5130_35948# VPWR 0.414005f
C322 a_3762_32076# VPWR 0.430937f
C323 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.02481f
C324 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.205884f
C325 a_3762_28204# VPWR 0.360178f
C326 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.Y 0.649845f
C327 SUNSAR_SAR8B_CV_0.EN ui_in[0] 0.96947f
C328 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR 0.709798f
C329 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP 0.123668f
C330 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.155714f
C331 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR 4.14837f
C332 SUNSAR_SAR8B_CV_0.XA7.XA10.Y a_21402_36300# 0.13402f
C333 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C334 a_9990_4038# VPWR 0.377115f
C335 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.152047f
C336 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.732448f
C337 a_10190_40648# VPWR 0.489635f
C338 a_3762_35068# VPWR 0.391042f
C339 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 27.1383f
C340 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35420# 0.160931f
C341 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.424961f
C342 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.779324f
C343 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.152662f
C344 a_3762_35948# VPWR 0.414005f
C345 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.Y 0.744161f
C346 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.EN 0.200133f
C347 SUNSAR_SAR8B_CV_0.XA4.CEO VPWR 2.15714f
C348 SUNSAR_SAR8B_CV_0.XB1.XA4.GN ua[1] 0.636092f
C349 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_4688# 0.172147f
C350 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR 2.29796f
C351 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.234118f
C352 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.339883f
C353 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VPWR 1.74633f
C354 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y uo_out[4] 0.246316f
C355 a_8822_40648# VPWR 0.488227f
C356 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VPWR 0.263064f
C357 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_20250_35420# 0.133834f
C358 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.141203f
C359 a_10170_27148# VPWR 0.468331f
C360 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.204048f
C361 a_20270_41880# VPWR 0.393193f
C362 SUNSAR_SAR8B_CV_0.XA0.XA2.A a_3762_30316# 0.129098f
C363 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 27.1383f
C364 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR 0.59973f
C365 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR 0.418836f
C366 a_10190_42760# VPWR 0.388849f
C367 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR 0.707016f
C368 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C369 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.680649f
C370 SUNSAR_SAR8B_CV_0.XB2.CKN VPWR 2.29833f
C371 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR 2.8981f
C372 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y uo_out[4] 0.305131f
C373 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.732438f
C374 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.51035f
C375 SUNSAR_SAR8B_CV_0.XA6.XA11.Y a_17730_36828# 0.10248f
C376 a_8802_27148# VPWR 0.468818f
C377 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.331207f
C378 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.432466f
C379 a_18902_41880# VPWR 0.393193f
C380 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.269899f
C381 SUNSAR_SAR8B_CV_0.XA20.XA10.B VPWR 1.11141f
C382 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR 0.311444f
C383 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.155132f
C384 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.D VPWR 0.127851f
C385 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.437765f
C386 a_8822_42760# VPWR 0.388849f
C387 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.148254f
C388 SUNSAR_SAR8B_CV_0.XA3.CEO VPWR 1.02323f
C389 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.156507f
C390 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR 4.154931f
C391 SUNSAR_SAR8B_CV_0.SARP ua[1] 0.946602f
C392 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.318734f
C393 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C394 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR 2.11326f
C395 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.ENO 0.486144f
C396 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35068# 0.129098f
C397 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C398 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.12241f
C399 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.584654f
C400 SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR 0.758315f
C401 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR 2.23433f
C402 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.205884f
C403 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.15291f
C404 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VPWR 1.04342f
C405 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.428385f
C406 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR 0.709829f
C407 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.CK 1.59176f
C408 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.734068f
C409 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.154155f
C410 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR 0.100103f
C411 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.D<2> 0.362022f
C412 a_5150_40648# VPWR 0.489605f
C413 SUNSAR_SAR8B_CV_0.XA6.DONE VPWR 0.236517f
C414 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA10.Y 0.303978f
C415 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6267f
C416 a_20250_30316# VPWR 0.400467f
C417 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_18882_35420# 0.133834f
C418 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 3.85159f
C419 SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR 0.762903f
C420 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR 2.24344f
C421 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.210891f
C422 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.D VPWR 0.128309f
C423 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.63636f
C424 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.177648f
C425 SUNSAR_SAR8B_CV_0.XA2.CEO VPWR 2.15721f
C426 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_5648# 0.172147f
C427 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.401945f
C428 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C429 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR 2.89809f
C430 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.3401f
C431 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_SAR8B_CV_0.D<2> 0.238616f
C432 a_3782_40648# VPWR 0.488227f
C433 SUNSAR_SAR8B_CV_0.XA5.DONE VPWR 0.235812f
C434 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.13078f
C435 SUNSAR_SAR8B_CV_0.XA5.XA11.Y a_16362_36828# 0.104051f
C436 a_18882_30316# VPWR 0.400438f
C437 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35420# 0.160931f
C438 a_5130_27148# VPWR 0.468331f
C439 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.204048f
C440 a_15230_41880# VPWR 0.393193f
C441 SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR 0.762889f
C442 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6267f
C443 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR 2.24344f
C444 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.133184f
C445 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VPWR 1.04916f
C446 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.164715f
C447 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.428385f
C448 a_5150_42760# VPWR 0.388849f
C449 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.140524f
C450 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR 0.706998f
C451 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.155714f
C452 SUNSAR_SAR8B_CV_0.XA6.XA10.Y a_17730_36300# 0.13253f
C453 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C454 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_2928# 0.105547f
C455 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VPWR 1.74633f
C456 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y uo_out[5] 0.305288f
C457 SUNSAR_SAR8B_CV_0.XA4.DONE VPWR 0.236517f
C458 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.51035f
C459 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.142931f
C460 a_3762_27148# VPWR 0.468818f
C461 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.428385f
C462 a_13862_41880# VPWR 0.393193f
C463 SUNSAR_SAR8B_CV_0.XA0.CEIN a_13950_4390# 0.155588f
C464 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.132976f
C465 SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR 0.762903f
C466 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR 2.24344f
C467 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.45988f
C468 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.D VPWR 0.127851f
C469 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.467457f
C470 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.Y 0.744161f
C471 a_3782_42760# VPWR 0.388849f
C472 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.161289f
C473 SUNSAR_SAR8B_CV_0.XA1.CEO VPWR 1.02323f
C474 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.144773f
C475 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.36495f
C476 SUNSAR_SAR8B_CV_0.XB1.CKN VPWR 2.29833f
C477 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.401945f
C478 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR 0.100103f
C479 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y uo_out[5] 0.246118f
C480 SUNSAR_SAR8B_CV_0.DONE VPWR 7.66429f
C481 SUNSAR_SAR8B_CV_0.XA3.DONE VPWR 0.235812f
C482 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.331639f
C483 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.ENO 0.106942f
C484 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.118161f
C485 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.12241f
C486 SUNSAR_CAPT8B_CV_0.XA3.A ui_in[0] 0.170915f
C487 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.SARP 0.236656f
C488 SUNSAR_SAR8B_CV_0.XA0.CEIN a_12582_4390# 0.155588f
C489 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S 0.307018f
C490 SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR 0.762889f
C491 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR 2.24344f
C492 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.205884f
C493 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VPWR 1.03788f
C494 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.Y 0.649845f
C495 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CN1 0.462451f
C496 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.140524f
C497 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR 0.713854f
C498 SUNSAR_SAR8B_CV_0.XA5.XA6.MP2.D VPWR 0.105892f
C499 SUNSAR_SAR8B_CV_0.XA5.XA10.Y a_16362_36300# 0.13402f
C500 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C501 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA6.ENO 0.29162f
C502 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR 2.29796f
C503 a_23942_41000# VPWR 0.387891f
C504 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.DONE 0.34047f
C505 SUNSAR_SAR8B_CV_0.XA2.DONE VPWR 0.236517f
C506 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.51035f
C507 a_15210_30316# VPWR 0.400991f
C508 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35068# 0.127528f
C509 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.428385f
C510 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.13041f
C511 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.432466f
C512 SUNSAR_CAPT8B_CV_0.XA3.A clk 0.187716f
C513 SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR 0.762903f
C514 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR 2.24344f
C515 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.221335f
C516 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.D VPWR 0.128309f
C517 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.233892f
C518 SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR 8.60088f
C519 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.161289f
C520 SUNSAR_SAR8B_CV_0.XA0.CEO VPWR 2.15876f
C521 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.156507f
C522 SUNSAR_SAR8B_CV_0.XA4.XA6.MP2.D VPWR 0.105892f
C523 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y 0.318734f
C524 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR 0.652264f
C525 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_6608# 0.172147f
C526 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C527 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VPWR 1.74633f
C528 SUNSAR_CAPT8B_CV_0.XA5.A SUNSAR_CAPT8B_CV_0.XA3.A 0.480936f
C529 SUNSAR_SAR8B_CV_0.XA1.DONE VPWR 0.235812f
C530 a_13842_30316# VPWR 0.400991f
C531 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.141203f
C532 a_20250_27500# VPWR 0.380285f
C533 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.118161f
C534 a_10190_41880# VPWR 0.393193f
C535 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.43622f
C536 SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR 0.762889f
C537 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR 2.24344f
C538 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.5128f
C539 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VPWR 1.04916f
C540 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.140524f
C541 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CN1 0.462451f
C542 SUNSAR_SAR8B_CV_0.EN VPWR 41.0271f
C543 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<0> 0.131191f
C544 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR 4.14921f
C545 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA1.Y 0.130935f
C546 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_3888# 0.105547f
C547 a_16542_4566# VPWR 0.41043f
C548 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.175492f
C549 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR 2.89805f
C550 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.35822f
C551 SUNSAR_SAR8B_CV_0.XA0.DONE VPWR 0.237772f
C552 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 54.1913f
C553 SUNSAR_SAR8B_CV_0.XA4.XA11.Y a_12690_36828# 0.10248f
C554 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEIN 0.215804f
C555 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35420# 0.160931f
C556 a_18882_27500# VPWR 0.380119f
C557 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.129613f
C558 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S 0.345133f
C559 a_8822_41880# VPWR 0.393193f
C560 SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR 0.766864f
C561 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR 2.24344f
C562 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.D VPWR 0.127851f
C563 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_3334# 0.120003f
C564 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.161289f
C565 a_23942_43112# VPWR 0.390941f
C566 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<0> 0.280677f
C567 a_20250_37180# VPWR 0.466603f
C568 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_ON 2.71492f
C569 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C570 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y uo_out[6] 0.250672f
C571 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_SAR8B_CV_0.D<3> 0.238616f
C572 a_20270_41000# VPWR 0.385556f
C573 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.DONE 0.150219f
C574 a_23922_35420# VPWR 0.413536f
C575 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_15210_35420# 0.133834f
C576 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.118226f
C577 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y a_7670_42408# 0.100131f
C578 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.150581f
C579 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 1.43616f
C580 a_23922_36300# VPWR 0.469729f
C581 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR 4.61168f
C582 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.205884f
C583 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_3334# 0.109848f
C584 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VPWR 1.03788f
C585 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.412248f
C586 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.140524f
C587 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CN1 0.462451f
C588 a_18882_37180# VPWR 0.470629f
C589 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.155714f
C590 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C591 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR 0.652264f
C592 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.152047f
C593 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.44669f
C594 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y uo_out[6] 0.306831f
C595 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR 0.100103f
C596 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.D<3> 0.362008f
C597 a_18902_41000# VPWR 0.385652f
C598 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.51035f
C599 a_10170_30316# VPWR 0.400991f
C600 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.530644f
C601 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.13041f
C602 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 3.99906f
C603 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.432466f
C604 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.221348f
C605 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.D VPWR 0.128309f
C606 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.63636f
C607 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.476106f
C608 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<1> 0.1286f
C609 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR 4.17894f
C610 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.29886f
C611 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.318734f
C612 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C613 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145003f
C614 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR 2.89806f
C615 SUNSAR_SAR8B_CV_0.XA3.XA11.Y a_11322_36828# 0.104051f
C616 a_8802_30316# VPWR 0.400991f
C617 a_15210_27500# VPWR 0.380285f
C618 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.118161f
C619 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C620 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.12241f
C621 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S 0.314697f
C622 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.204048f
C623 a_5150_41880# VPWR 0.393193f
C624 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.793386f
C625 a_20250_32956# VPWR 0.42896f
C626 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_2982# 0.157687f
C627 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VPWR 1.04916f
C628 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARN 0.567675f
C629 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.412248f
C630 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CN1 0.462451f
C631 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VPWR 1.58781f
C632 SUNSAR_SAR8B_CV_0.XA4.XA10.Y a_12690_36300# 0.13253f
C633 SUNSAR_SAR8B_CV_0.SARP VPWR 0.138198f
C634 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43816# 0.129239f
C635 a_9990_4566# VPWR 0.41043f
C636 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_4848# 0.105547f
C637 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VPWR 1.74633f
C638 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.DONE 0.150402f
C639 a_20250_35420# VPWR 0.39359f
C640 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 6.84356f
C641 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.163923f
C642 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.142931f
C643 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_13842_35420# 0.133834f
C644 a_13842_27500# VPWR 0.380119f
C645 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.412248f
C646 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.21768f
C647 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.129613f
C648 a_3782_41880# VPWR 0.393193f
C649 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.149398f
C650 a_20250_36300# VPWR 0.392819f
C651 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.ENO 0.821625f
C652 a_18882_32956# VPWR 0.430937f
C653 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.D VPWR 0.127851f
C654 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARP 0.520264f
C655 a_15210_37180# VPWR 0.470519f
C656 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.156507f
C657 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VPWR 0.428795f
C658 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C659 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C660 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR 0.100103f
C661 a_15230_41000# VPWR 0.385556f
C662 a_18882_35420# VPWR 0.396084f
C663 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35420# 0.160931f
C664 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.398211f
C665 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.118226f
C666 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_23922_29964# 0.151031f
C667 a_18882_36300# VPWR 0.395565f
C668 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.ENO 0.837821f
C669 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.205884f
C670 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C671 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VPWR 1.03788f
C672 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CN1 0.462451f
C673 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<2> 0.129233f
C674 a_13842_37180# VPWR 0.470643f
C675 SUNSAR_SAR8B_CV_0.XA3.XA10.Y a_11322_36300# 0.13402f
C676 a_20250_29612# VPWR 0.395402f
C677 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_2768# 0.172147f
C678 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y uo_out[7] 0.308468f
C679 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA1.Y 0.227108f
C680 a_13862_41000# VPWR 0.385652f
C681 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.351225f
C682 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.292709f
C683 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.1913f
C684 a_5130_30316# VPWR 0.400991f
C685 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.412248f
C686 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.13041f
C687 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.24317f
C688 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.SARP 0.532453f
C689 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S 0.345133f
C690 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_22770_29964# 0.134249f
C691 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR 0.11134f
C692 SUNSAR_CAPT8B_CV_0.XA3.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.138433f
C693 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.ENO 0.888066f
C694 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.221335f
C695 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.D VPWR 0.128309f
C696 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.107674f
C697 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VPWR 1.58781f
C698 a_18882_29612# VPWR 0.394799f
C699 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C700 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y uo_out[7] 0.248878f
C701 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VPWR 1.74633f
C702 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y a_20270_41880# 0.100592f
C703 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.DONE 0.150216f
C704 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.CEO 0.136315f
C705 a_3762_30316# VPWR 0.400991f
C706 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.141203f
C707 a_10170_27500# VPWR 0.380285f
C708 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.118161f
C709 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C710 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.74007f
C711 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.12241f
C712 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.204048f
C713 SUNSAR_CAPT8B_CV_0.XA3.A VPWR 1.18393f
C714 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.ENO 0.837821f
C715 a_15210_32956# VPWR 0.430937f
C716 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.379169p
C717 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_2982# 0.157687f
C718 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VPWR 1.04916f
C719 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.164715f
C720 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.510531f
C721 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.155714f
C722 SUNSAR_SAR8B_CV_0.XA3.XA6.MP2.D VPWR 0.105892f
C723 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43816# 0.127669f
C724 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR 0.515447f
C725 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_5808# 0.105547f
C726 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR 2.89812f
C727 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.D<4> 0.362014f
C728 a_15210_35420# VPWR 0.396084f
C729 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1383f
C730 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.148207f
C731 SUNSAR_SAR8B_CV_0.XA2.XA11.Y a_7650_36828# 0.10248f
C732 a_8802_27500# VPWR 0.380119f
C733 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.129613f
C734 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.432466f
C735 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.153225f
C736 SUNSAR_SAR8B_CV_0.XA0.CEIN a_13950_4742# 0.156329f
C737 a_15210_36300# VPWR 0.395313f
C738 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.ENO 0.888066f
C739 a_13842_32956# VPWR 0.430937f
C740 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.175568f
C741 a_23922_28556# VPWR 0.496622f
C742 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<3> 0.1286f
C743 a_10170_37180# VPWR 0.470548f
C744 SUNSAR_SAR8B_CV_0.XA2.XA6.MP2.D VPWR 0.105892f
C745 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y 0.318734f
C746 a_16542_4918# VPWR 0.46774f
C747 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.257673f
C748 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y VPWR 0.748775f
C749 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_SAR8B_CV_0.D<4> 0.238616f
C750 a_10190_41000# VPWR 0.385576f
C751 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.356354f
C752 a_13842_35420# VPWR 0.396084f
C753 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR 6.57457f
C754 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.118226f
C755 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.EN 0.128277f
C756 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S 0.314697f
C757 SUNSAR_SAR8B_CV_0.XA0.CEIN a_12582_4742# 0.156329f
C758 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR 0.100103f
C759 a_13842_36300# VPWR 0.395565f
C760 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.33518f
C761 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.ENO 0.837821f
C762 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C763 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.205884f
C764 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.646191f
C765 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3334# 0.162056f
C766 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_3334# 0.111418f
C767 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.440597f
C768 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.521227f
C769 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VPWR 1.58781f
C770 a_8802_37180# VPWR 0.470672f
C771 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR 4.1452f
C772 a_15210_29612# VPWR 0.394799f
C773 SUNSAR_CAPT8B_CV_0.XG12.QN a_16382_43816# 0.129239f
C774 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_3728# 0.172147f
C775 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.153899f
C776 a_8822_41000# VPWR 0.385652f
C777 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.DONE 0.150309f
C778 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.220689f
C779 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.84356f
C780 a_23922_30844# VPWR 0.422642f
C781 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35420# 0.160931f
C782 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.527529f
C783 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.13041f
C784 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.2954f
C785 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.CMP_OP 7.91015f
C786 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR 0.100103f
C787 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_28556# 0.140127f
C788 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.ENO 0.905126f
C789 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.221348f
C790 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_3334# 0.118433f
C791 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.63636f
C792 a_13842_29612# VPWR 0.394799f
C793 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR 0.515447f
C794 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.424961f
C795 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C796 a_20270_43816# VPWR 0.38934f
C797 SUNSAR_SAR8B_CV_0.XA1.XA11.Y a_6282_36828# 0.104051f
C798 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_10170_35420# 0.133834f
C799 a_5130_27500# VPWR 0.380285f
C800 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.118161f
C801 a_10170_32956# VPWR 0.430937f
C802 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C803 a_20250_28556# VPWR 0.403733f
C804 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.440597f
C805 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<4> 0.129233f
C806 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C807 SUNSAR_SAR8B_CV_0.XA2.XA10.Y a_7650_36300# 0.13253f
C808 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VPWR 0.428795f
C809 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_6768# 0.105547f
C810 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.196077f
C811 a_18902_43816# VPWR 0.38934f
C812 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.07747f
C813 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.301485f
C814 ua[1] ua[0] 3.85014f
C815 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6267f
C816 a_10170_35420# VPWR 0.396084f
C817 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.377598f
C818 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR 2.3695f
C819 a_3762_27500# VPWR 0.380119f
C820 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.440597f
C821 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 5.16845f
C822 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.432466f
C823 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S 0.345133f
C824 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.157855f
C825 a_10170_36300# VPWR 0.395313f
C826 a_8802_32956# VPWR 0.430937f
C827 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_4038# 0.135341f
C828 a_18882_28556# VPWR 0.403733f
C829 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VPWR 1.58781f
C830 a_5130_37180# VPWR 0.470533f
C831 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR 4.15202f
C832 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.40651f
C833 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.127043f
C834 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.424961f
C835 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.28008f
C836 a_5150_41000# VPWR 0.385562f
C837 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.DONE 0.150615f
C838 a_8802_35420# VPWR 0.396084f
C839 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR 2.3676f
C840 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y a_2630_42408# 0.100131f
C841 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.12241f
C842 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR 0.100103f
C843 a_8802_36300# VPWR 0.395565f
C844 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3686# 0.163645f
C845 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3334# 0.162056f
C846 a_3762_37180# VPWR 0.470657f
C847 SUNSAR_SAR8B_CV_0.XA1.XA10.Y a_6282_36300# 0.13402f
C848 a_10170_29612# VPWR 0.394799f
C849 SUNSAR_CAPT8B_CV_0.XF11.QN a_12710_43816# 0.127669f
C850 a_9990_4918# VPWR 0.466169f
C851 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_4688# 0.172147f
C852 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.55788f
C853 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[0] 0.199387f
C854 a_3782_41000# VPWR 0.385652f
C855 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.270239f
C856 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1383f
C857 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR 2.3707f
C858 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_8802_35420# 0.133834f
C859 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.440597f
C860 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C861 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.SARP 5.15147f
C862 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR 0.100103f
C863 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.220575f
C864 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.233892f
C865 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<5> 0.1286f
C866 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y SUNSAR_CAPT8B_CV_0.XA3.A 0.297144f
C867 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y a_21422_41000# 0.115667f
C868 a_8802_29612# VPWR 0.394799f
C869 a_15230_43816# VPWR 0.38934f
C870 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.63098f
C871 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_SAR8B_CV_0.D<5> 0.238616f
C872 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.CEO 0.277778f
C873 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR 2.3707f
C874 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35420# 0.160931f
C875 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA8.A 0.527529f
C876 a_20250_27852# VPWR 0.357005f
C877 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.204048f
C878 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S 0.314697f
C879 a_5130_32956# VPWR 0.430937f
C880 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C881 a_15210_28556# VPWR 0.403733f
C882 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.175568f
C883 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VPWR 1.58781f
C884 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y a_20270_41000# 0.156079f
C885 SUNSAR_SAR8B_CV_0.XA1.XA6.MP2.D VPWR 0.105892f
C886 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43816# 0.129239f
C887 a_13862_43816# VPWR 0.38934f
C888 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.547785f
C889 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.301485f
C890 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22790_42760# 0.133036f
C891 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.D<5> 0.362034f
C892 clk ui_in[0] 0.169425f
C893 a_23942_41352# VPWR 0.373866f
C894 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.351225f
C895 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.DONE 0.150831f
C896 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.51035f
C897 a_5130_35420# VPWR 0.396084f
C898 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.148207f
C899 SUNSAR_SAR8B_CV_0.XA0.XA11.Y a_2610_36828# 0.10248f
C900 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR 2.3707f
C901 a_18882_27852# VPWR 0.357158f
C902 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.699044f
C903 a_5130_36300# VPWR 0.395313f
C904 a_3762_32956# VPWR 0.430937f
C905 a_13842_28556# VPWR 0.403733f
C906 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.379169p
C907 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.646191f
C908 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C909 a_20250_37532# VPWR 0.4511f
C910 SUNSAR_SAR8B_CV_0.XA0.XA6.MP2.D VPWR 0.105892f
C911 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.185068f
C912 a_16542_5270# VPWR 0.486169f
C913 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW clk 0.197555f
C914 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.63098f
C915 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA3.A 0.254583f
C916 a_3762_35420# VPWR 0.396084f
C917 SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR 2.3707f
C918 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C919 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.12241f
C920 SUNSAR_SAR8B_CV_0.XA0.CEIN a_13950_5094# 0.160184f
C921 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR 0.100103f
C922 a_3762_36300# VPWR 0.395565f
C923 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.CEO 0.300333f
C924 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C925 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3686# 0.163645f
C926 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.401945f
C927 SUNSAR_CAPT8B_CV_0.XA5.A clk 0.20527f
C928 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<6> 0.129233f
C929 a_18882_37532# VPWR 0.454256f
C930 a_5130_29612# VPWR 0.394799f
C931 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_5648# 0.172147f
C932 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.547785f
C933 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.220689f
C934 SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR 2.3707f
C935 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6267f
C936 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.31012f
C937 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.432466f
C938 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.Y 0.649845f
C939 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S 0.345133f
C940 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.228693f
C941 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.699044f
C942 SUNSAR_SAR8B_CV_0.XA0.CEIN a_12582_5094# 0.160184f
C943 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR 0.100103f
C944 SUNSAR_SAR8B_CV_0.XA6.ENO a_17730_28556# 0.132757f
C945 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR 4.78095f
C946 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.220593f
C947 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.133554f
C948 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y SUNSAR_CAPT8B_CV_0.XA3.Y 0.342913f
C949 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.63636f
C950 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VPWR 1.58781f
C951 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR 2.57982f
C952 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.51035f
C953 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.710435f
C954 a_3762_29612# VPWR 0.394799f
C955 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.428385f
C956 a_10190_43816# VPWR 0.38934f
C957 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.63098f
C958 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.24396f
C959 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.44051f
C960 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y a_15230_41880# 0.100592f
C961 a_20270_41352# VPWR 0.391367f
C962 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.356354f
C963 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.DONE 0.147658f
C964 SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR 2.3707f
C965 a_15210_27852# VPWR 0.357005f
C966 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.380687f
C967 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA5.Y 0.744161f
C968 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.232226f
C969 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.204048f
C970 a_23922_36652# VPWR 0.446957f
C971 a_23922_33132# VPWR 0.4125f
C972 a_10170_28556# VPWR 0.403733f
C973 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.154933f
C974 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.401945f
C975 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.440586f
C976 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C977 SUNSAR_SAR8B_CV_0.XA0.XA10.Y a_2610_36300# 0.13253f
C978 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C979 a_9990_5270# VPWR 0.48774f
C980 a_8822_43816# VPWR 0.38934f
C981 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.15919f
C982 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.547785f
C983 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.301485f
C984 uo_out[1] uo_out[0] 0.366518f
C985 a_18902_41352# VPWR 0.391367f
C986 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 3.51035f
C987 SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR 0.646249f
C988 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.377598f
C989 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35420# 0.160931f
C990 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.401945f
C991 a_13842_27852# VPWR 0.357158f
C992 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.699044f
C993 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.109021f
C994 SUNSAR_SAR8B_CV_0.XA5.ENO a_16362_28556# 0.135264f
C995 a_8802_28556# VPWR 0.403733f
C996 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y a_22790_43640# 0.127669f
C997 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<7> 0.162541f
C998 a_15210_37532# VPWR 0.455459f
C999 a_20250_34716# VPWR 0.393873f
C1000 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR 0.324956f
C1001 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR 0.796216f
C1002 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.428385f
C1003 SUNSAR_CAPT8B_CV_0.XI14.QN uo_out[0] 0.256493f
C1004 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.83572f
C1005 a_20250_31196# VPWR 0.431145f
C1006 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_5130_35420# 0.133834f
C1007 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.126085f
C1008 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C1009 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR 0.100103f
C1010 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR 0.705366f
C1011 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR 2.57273f
C1012 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C1013 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VPWR 1.58781f
C1014 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y a_18902_41000# 0.15757f
C1015 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<7> 0.274892f
C1016 a_13842_37532# VPWR 0.454304f
C1017 a_18882_34716# VPWR 0.396368f
C1018 a_23922_29964# VPWR 0.425757f
C1019 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C1020 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_6608# 0.172147f
C1021 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_2928# 0.105547f
C1022 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.241632f
C1023 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.D<6> 0.362018f
C1024 SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR 1.18991f
C1025 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.270239f
C1026 a_18882_31196# VPWR 0.433639f
C1027 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.51035f
C1028 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA8.A 0.527529f
C1029 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.401945f
C1030 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.11382f
C1031 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.432466f
C1032 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.699044f
C1033 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR 0.100103f
C1034 SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR 2.54505f
C1035 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.586572f
C1036 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CP0 0.318407f
C1037 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_4038# 0.135341f
C1038 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y a_17750_41000# 0.114097f
C1039 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 54.1913f
C1040 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.0194f
C1041 SUNSAR_CAPT8B_CV_0.XH13.QN uo_out[1] 0.252841f
C1042 a_5150_43816# VPWR 0.38934f
C1043 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_SAR8B_CV_0.D<6> 0.238616f
C1044 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y a_20270_42760# 0.111734f
C1045 VPWR ua[0] 0.425538f
C1046 a_15230_41352# VPWR 0.391367f
C1047 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR 0.903837f
C1048 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.CEO 0.277778f
C1049 a_10170_27852# VPWR 0.357005f
C1050 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.238103f
C1051 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.12241f
C1052 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR 0.112284f
C1053 SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR 2.54504f
C1054 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C1055 a_5130_28556# VPWR 0.403733f
C1056 a_16542_5622# VPWR 0.469729f
C1057 a_3782_43816# VPWR 0.38934f
C1058 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.301485f
C1059 VPWR ua[1] 0.188995f
C1060 uo_out[3] uo_out[2] 0.110015f
C1061 a_13862_41352# VPWR 0.391367f
C1062 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 54.1921f
C1063 SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR 1.19836f
C1064 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.148207f
C1065 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_3762_35420# 0.133834f
C1066 a_8802_27852# VPWR 0.357158f
C1067 a_23942_42408# VPWR 0.388942f
C1068 SUNSAR_SAR8B_CV_0.XA0.CEIN a_13950_5446# 0.102601f
C1069 SUNSAR_SAR8B_CV_0.XA4.ENO a_12690_28556# 0.132757f
C1070 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.108318f
C1071 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.699044f
C1072 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR 0.711145f
C1073 SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR 2.54505f
C1074 a_3762_28556# VPWR 0.403733f
C1075 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 0.635098f
C1076 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VPWR 1.58781f
C1077 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1078 a_10170_37532# VPWR 0.455561f
C1079 a_15210_34716# VPWR 0.396368f
C1080 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR 0.10219f
C1081 SUNSAR_CAPT8B_CV_0.XG12.QN uo_out[2] 0.253231f
C1082 VPWR ui_in[0] 1.07924f
C1083 SUNSAR_CAPT8B_CV_0.XA4.MP1.G clk 0.432892f
C1084 a_15210_31196# VPWR 0.433639f
C1085 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35420# 0.160931f
C1086 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.283764f
C1087 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.Y 0.744161f
C1088 SUNSAR_SAR8B_CV_0.XA0.CEIN a_12582_5446# 0.101031f
C1089 SUNSAR_SAR8B_CV_0.XA0.CEIN ua[0] 0.932378f
C1090 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR 0.708932f
C1091 SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR 2.54504f
C1092 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.244746f
C1093 SUNSAR_CAPT8B_CV_0.XA5.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.197749f
C1094 a_8802_37532# VPWR 0.454405f
C1095 a_13842_34716# VPWR 0.396368f
C1096 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VPWR 0.269339f
C1097 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C1098 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARP 0.177799f
C1099 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C1100 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_3888# 0.105547f
C1101 a_16542_5974# VPWR 0.44699f
C1102 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR 11.4501f
C1103 uo_out[4] uo_out[3] 0.857214f
C1104 VPWR clk 0.669028f
C1105 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.351225f
C1106 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR 0.908851f
C1107 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.220689f
C1108 a_13842_31196# VPWR 0.433639f
C1109 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.51035f
C1110 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA5.Y 0.649845f
C1111 SUNSAR_SAR8B_CV_0.XA3.ENO a_11322_28556# 0.135264f
C1112 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.733192f
C1113 SUNSAR_SAR8B_CV_0.XA0.CEIN ua[1] 0.658951f
C1114 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR 2.61784f
C1115 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.373421f
C1116 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.314981f
C1117 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.CKN 0.413022f
C1118 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.63636f
C1119 SUNSAR_CAPT8B_CV_0.XA5.A VPWR 1.17045f
C1120 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y a_16382_41000# 0.115667f
C1121 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.139824f
C1122 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 6.84356f
C1123 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.412248f
C1124 a_23942_43992# VPWR 0.339461f
C1125 SUNSAR_CAPT8B_CV_0.XF11.QN uo_out[3] 0.264123f
C1126 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y a_18902_42760# 0.113305f
C1127 VPWR uo_out[0] 1.14289f
C1128 a_10190_41352# VPWR 0.391367f
C1129 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.282403f
C1130 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA8.A 0.527529f
C1131 a_5130_27852# VPWR 0.357005f
C1132 a_20270_42408# VPWR 0.388814f
C1133 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.204048f
C1134 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR 0.112284f
C1135 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.154344f
C1136 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR 2.6168f
C1137 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C1138 a_20250_28908# VPWR 0.392546f
C1139 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C1140 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y a_15230_41000# 0.156079f
C1141 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1142 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR 0.796216f
C1143 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.22402f
C1144 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.301485f
C1145 VPWR uo_out[1] 0.986945f
C1146 uo_out[5] uo_out[4] 1.16561f
C1147 a_8822_41352# VPWR 0.391367f
C1148 SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR 1.19834f
C1149 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 6.84356f
C1150 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.377598f
C1151 a_3762_27852# VPWR 0.357158f
C1152 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.5424f
C1153 a_18902_42408# VPWR 0.388814f
C1154 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.734928f
C1155 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.106747f
C1156 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XA0.CEIN 4.16332f
C1157 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR 0.711145f
C1158 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR 2.61938f
C1159 a_18882_28908# VPWR 0.392546f
C1160 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.310451f
C1161 a_20270_43288# VPWR 0.39173f
C1162 a_5130_37532# VPWR 0.455509f
C1163 a_10170_34716# VPWR 0.396368f
C1164 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.771246f
C1165 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S 0.145483f
C1166 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO 0.144331f
C1167 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.412248f
C1168 SUNSAR_CAPT8B_CV_0.XI14.QN VPWR 0.882006f
C1169 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[4] 0.248279f
C1170 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.224581f
C1171 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_SAR8B_CV_0.D<7> 0.238616f
C1172 VPWR uo_out[2] 0.987117f
C1173 uo_out[6] uo_out[4] 0.815262f
C1174 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.356354f
C1175 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR 0.908827f
C1176 a_10170_31196# VPWR 0.433639f
C1177 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR 0.708932f
C1178 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.422121f
C1179 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.152326f
C1180 a_18902_43288# VPWR 0.39173f
C1181 a_3762_37532# VPWR 0.454354f
C1182 a_8802_34716# VPWR 0.396368f
C1183 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_4848# 0.105547f
C1184 a_9990_5622# VPWR 0.468158f
C1185 SUNSAR_CAPT8B_CV_0.XH13.QN VPWR 0.881997f
C1186 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.D<7> 0.362082f
C1187 VPWR uo_out[3] 1.19648f
C1188 uo_out[7] uo_out[4] 0.119113f
C1189 uo_out[6] uo_out[5] 0.317731f
C1190 SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR 1.19836f
C1191 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.270239f
C1192 a_8802_31196# VPWR 0.433639f
C1193 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.1913f
C1194 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.136678f
C1195 SUNSAR_SAR8B_CV_0.XA2.ENO a_7650_28556# 0.132757f
C1196 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.108318f
C1197 a_20250_33836# VPWR 0.40361f
C1198 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.315699f
C1199 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN 0.133554f
C1200 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.233892f
C1201 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.340483f
C1202 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 27.1383f
C1203 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S 0.145483f
C1204 SUNSAR_CAPT8B_CV_0.XG12.QN VPWR 0.881997f
C1205 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[5] 0.2482f
C1206 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y a_10190_41880# 0.100592f
C1207 VPWR uo_out[4] 0.993845f
C1208 uo_out[7] uo_out[5] 1.58097f
C1209 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP 0.435464f
C1210 a_5150_41352# VPWR 0.391367f
C1211 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.252557f
C1212 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.CEO 0.277778f
C1213 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.214181f
C1214 a_15230_42408# VPWR 0.388814f
C1215 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.DONE 0.367606f
C1216 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR 0.112284f
C1217 a_18882_33836# VPWR 0.405586f
C1218 a_15210_28908# VPWR 0.392546f
C1219 a_16542_2630# VPWR 0.446313f
C1220 a_23942_40296# VPWR 0.449779f
C1221 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VPWR 0.263064f
C1222 a_9990_5974# VPWR 0.448145f
C1223 SUNSAR_CAPT8B_CV_0.XF11.QN VPWR 0.881997f
C1224 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.301485f
C1225 VPWR uo_out[5] 0.992028f
C1226 uo_out[7] uo_out[6] 2.3808f
C1227 a_3782_41352# VPWR 0.391367f
C1228 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR 0.908851f
C1229 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 27.139301f
C1230 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.148207f
C1231 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.Y 0.649845f
C1232 a_13862_42408# VPWR 0.388814f
C1233 SUNSAR_SAR8B_CV_0.XA1.ENO a_6282_28556# 0.135264f
C1234 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR 0.711145f
C1235 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.CKN 0.190344f
C1236 a_13842_28908# VPWR 0.392546f
C1237 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.424961f
C1238 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARP 0.476511f
C1239 a_15230_43288# VPWR 0.39173f
C1240 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y a_22790_42408# 0.10248f
C1241 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1242 a_5130_34716# VPWR 0.396368f
C1243 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S 0.145483f
C1244 a_23922_26796# VPWR 0.440719f
C1245 SUNSAR_CAPT8B_CV_0.XE10.QN VPWR 0.881997f
C1246 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[6] 0.255878f
C1247 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y a_15230_42760# 0.111734f
C1248 VPWR uo_out[6] 1.27969f
C1249 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.27006f
C1250 a_5130_31196# VPWR 0.433639f
C1251 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA5.Y 0.744161f
C1252 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR 0.708932f
C1253 SUNSAR_SAR8B_CV_0.SARN ua[0] 0.953801f
C1254 a_13862_43288# VPWR 0.39173f
C1255 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y a_13862_41000# 0.15757f
C1256 a_3762_34716# VPWR 0.396368f
C1257 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35068# 0.129098f
C1258 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO 0.144331f
C1259 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_5808# 0.105547f
C1260 SUNSAR_CAPT8B_CV_0.XD09.QN VPWR 0.881997f
C1261 SUNSAR_CAPT8B_CV_0.XA5.A SUNSAR_CAPT8B_CV_0.XA5.XA1.Y 0.101177f
C1262 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.530413f
C1263 VPWR uo_out[7] 1.21778f
C1264 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR 0.624166f
C1265 SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR 1.19834f
C1266 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.84356f
C1267 a_3762_31196# VPWR 0.433639f
C1268 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA8.A 0.527529f
C1269 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.106747f
C1270 SUNSAR_SAR8B_CV_0.SARN ua[1] 0.757758f
C1271 a_15210_33836# VPWR 0.405586f
C1272 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.314981f
C1273 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.CKN 0.413022f
C1274 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.63636f
C1275 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_21422_42408# 0.113479f
C1276 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y a_12710_41000# 0.114097f
C1277 a_20270_40296# VPWR 0.452389f
C1278 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6267f
C1279 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105216f
C1280 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.31211f
C1281 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VPWR 0.263064f
C1282 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S 0.145483f
C1283 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.440597f
C1284 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.356301f
C1285 SUNSAR_CAPT8B_CV_0.XC08.QN VPWR 0.881997f
C1286 SUNSAR_CAPT8B_CV_0.XB07.QN uo_out[7] 0.260947f
C1287 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D 0.147973f
C1288 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR 0.908827f
C1289 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.104736f
C1290 a_10190_42408# VPWR 0.388814f
C1291 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR 0.112284f
C1292 a_13842_33836# VPWR 0.405586f
C1293 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 0.244746f
C1294 a_10170_28908# VPWR 0.392546f
C1295 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.424961f
C1296 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1297 a_18902_40296# VPWR 0.454411f
C1298 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR 3.86355f
C1299 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.195146f
C1300 a_20250_26796# VPWR 0.440138f
C1301 SUNSAR_CAPT8B_CV_0.XB07.QN VPWR 0.881997f
C1302 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.667435f
C1303 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.301485f
C1304 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.351092f
C1305 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.275206f
C1306 SUNSAR_SAR8B_CV_0.D<0> VPWR 4.8886f
C1307 SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR 1.19836f
C1308 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 13.6271f
C1309 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR 6.62954f
C1310 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA5.A 0.496756f
C1311 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.118266f
C1312 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.108318f
C1313 a_8822_42408# VPWR 0.388814f
C1314 SUNSAR_SAR8B_CV_0.XA0.ENO a_2610_28556# 0.132757f
C1315 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR 0.713544f
C1316 a_8802_28908# VPWR 0.392546f
C1317 a_9990_2630# VPWR 0.445157f
C1318 a_10190_43288# VPWR 0.39173f
C1319 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.152047f
C1320 a_23922_34892# VPWR 0.392835f
C1321 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S 0.145483f
C1322 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO 0.144331f
C1323 a_18882_26796# VPWR 0.441293f
C1324 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.440597f
C1325 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y a_13862_42760# 0.113305f
C1326 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D 0.146505f
C1327 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR 0.100103f
C1328 a_23922_31724# VPWR 0.409011f
C1329 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.161999f
C1330 SUNSAR_SAR8B_CV_0.XA0.CEIN VPWR 7.19758f
C1331 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 1.43616f
C1332 a_16542_2982# VPWR 0.487343f
C1333 a_8822_43288# VPWR 0.39173f
C1334 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.339883f
C1335 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.130369f
C1336 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.100252f
C1337 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.56776f
C1338 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_6768# 0.105547f
C1339 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.165155f
C1340 a_20270_44168# VPWR 0.338694f
C1341 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR 0.100103f
C1342 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR 0.908851f
C1343 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1383f
C1344 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.41354f
C1345 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S 0.142682f
C1346 a_10170_33836# VPWR 0.405586f
C1347 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.315699f
C1348 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_17750_42408# 0.111909f
C1349 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y a_11342_41000# 0.115667f
C1350 a_15230_40296# VPWR 0.452695f
C1351 SUNSAR_SAR8B_CV_0.XA7.ENO VPWR 4.36341f
C1352 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.51035f
C1353 SUNSAR_SAR8B_CV_0.XA0.CEIN SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.293873f
C1354 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S 0.145483f
C1355 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35068# 0.127528f
C1356 a_18902_44168# VPWR 0.339109f
C1357 SUNSAR_SAR8B_CV_0.D<1> VPWR 4.55777f
C1358 SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR 2.5308f
C1359 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA8.A 0.527529f
C1360 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.104736f
C1361 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.Y 0.744161f
C1362 a_5150_42408# VPWR 0.388814f
C1363 a_20250_36828# VPWR 0.389943f
C1364 a_8802_33836# VPWR 0.405586f
C1365 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.04737f
C1366 a_5130_28908# VPWR 0.392546f
C1367 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.132601f
C1368 SUNSAR_SAR8B_CV_0.XB2.XA3.B ua[0] 0.238743f
C1369 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y a_10190_41000# 0.156079f
C1370 a_13862_40296# VPWR 0.454411f
C1371 SUNSAR_SAR8B_CV_0.XA6.ENO VPWR 5.01862f
C1372 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.ENO 0.408515f
C1373 a_15210_26796# VPWR 0.440138f
C1374 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.779346f
C1375 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.20369f
C1376 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.301485f
C1377 SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR 1.19834f
C1378 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 3.52991f
C1379 SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR 2.52749f
C1380 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 0.588443f
C1381 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA5.Y 0.649845f
C1382 a_3782_42408# VPWR 0.388814f
C1383 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.10953f
C1384 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S 0.142644f
C1385 a_18882_36828# VPWR 0.392558f
C1386 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.128051f
C1387 a_3762_28908# VPWR 0.392546f
C1388 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S ua[0] 0.100365f
C1389 a_5150_43288# VPWR 0.39173f
C1390 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.154155f
C1391 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_16382_42408# 0.113479f
C1392 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1393 SUNSAR_SAR8B_CV_0.XA5.ENO VPWR 4.43046f
C1394 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.36023f
C1395 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S 0.145483f
C1396 a_13842_26796# VPWR 0.441293f
C1397 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.934205f
C1398 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D 0.150367f
C1399 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR 0.908827f
C1400 SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR 2.52762f
C1401 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.733529f
C1402 SUNSAR_SAR8B_CV_0.EN a_20250_29612# 0.142347f
C1403 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.133602f
C1404 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.242261f
C1405 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.201115f
C1406 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.428385f
C1407 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y uo_out[0] 0.245907f
C1408 a_3782_43288# VPWR 0.39173f
C1409 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.3401f
C1410 SUNSAR_SAR8B_CV_0.XA4.ENO VPWR 5.00372f
C1411 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.51035f
C1412 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VPWR 0.263064f
C1413 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO 0.144331f
C1414 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.965002f
C1415 a_15230_44168# VPWR 0.338694f
C1416 SUNSAR_SAR8B_CV_0.D<2> VPWR 4.58391f
C1417 SUNSAR_SAR8B_CV_0.XA7.XA2.A a_20250_30316# 0.127528f
C1418 SUNSAR_CAPT8B_CV_0.XA3.A a_22790_41000# 0.11811f
C1419 SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR 1.20157f
C1420 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6267f
C1421 SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR 2.52762f
C1422 SUNSAR_SAR8B_CV_0.EN a_18882_29612# 0.143511f
C1423 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y VPWR 0.675532f
C1424 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.111165f
C1425 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S 0.142624f
C1426 a_5130_33836# VPWR 0.405586f
C1427 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.12197f
C1428 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.63636f
C1429 SUNSAR_SAR8B_CV_0.XB1.XA3.B ua[1] 0.238743f
C1430 a_9990_2982# VPWR 0.488913f
C1431 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y uo_out[0] 0.307261f
C1432 a_10190_40296# VPWR 0.452786f
C1433 SUNSAR_SAR8B_CV_0.XA3.ENO VPWR 4.43046f
C1434 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S 0.17663f
C1435 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.401945f
C1436 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.356301f
C1437 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.885278f
C1438 a_13862_44168# VPWR 0.339109f
C1439 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y a_10190_42760# 0.111734f
C1440 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y a_5150_41880# 0.100592f
C1441 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.27006f
C1442 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D 0.146505f
C1443 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR 0.100103f
C1444 SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR 2.52762f
C1445 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.133602f
C1446 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR 0.877293f
C1447 a_15210_36828# VPWR 0.392437f
C1448 a_3762_33836# VPWR 0.405586f
C1449 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.61097f
C1450 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.ENO 0.791856f
C1451 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.318734f
C1452 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.428385f
C1453 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S ua[1] 0.100365f
C1454 a_16542_3334# VPWR 0.377065f
C1455 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.300065f
C1456 a_8822_40296# VPWR 0.454411f
C1457 SUNSAR_SAR8B_CV_0.XA2.ENO VPWR 5.00372f
C1458 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA10.Y 0.355906f
C1459 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.ENO 0.431783f
C1460 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35068# 0.129098f
C1461 a_10170_26796# VPWR 0.440138f
C1462 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.965002f
C1463 SUNSAR_SAR8B_CV_0.XA6.XA2.A a_18882_30316# 0.129098f
C1464 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR 0.100103f
C1465 ua[2] VGND 0.10961f
C1466 ua[3] VGND 0.10961f
C1467 ua[4] VGND 0.110707f
C1468 ua[5] VGND 0.111915f
C1469 ua[6] VGND 0.111915f
C1470 ua[7] VGND 0.103056f
C1471 ua[0] VGND 7.03068f
C1472 ua[1] VGND 6.38225f
C1473 ui_in[0] VGND 5.19924f
C1474 clk VGND 5.44899f
C1475 uo_out[0] VGND 2.73433f
C1476 uo_out[1] VGND 1.87119f
C1477 uo_out[2] VGND 1.57055f
C1478 uo_out[3] VGND 1.81511f
C1479 uo_out[4] VGND 1.73363f
C1480 uo_out[5] VGND 2.75265f
C1481 uo_out[6] VGND 2.5967f
C1482 uo_out[7] VGND 3.46094f
C1483 VPWR VGND 0.657889p
C1484 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 7.424201f
C1485 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 7.424201f
C1486 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 20.8457f
C1487 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 20.8457f
C1488 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 8.18329f
C1489 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 8.18329f
C1490 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 13.6417f
C1491 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 13.6417f
C1492 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 10.065901f
C1493 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 10.065901f
C1494 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 7.16564f
C1495 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 7.16564f
C1496 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 7.15659f
C1497 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 7.15659f
C1498 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 20.872f
C1499 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 20.872f
C1500 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 8.18273f
C1501 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 8.18273f
C1502 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 13.6417f
C1503 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 13.6417f
C1504 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 10.065901f
C1505 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 10.065901f
C1506 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 7.16564f
C1507 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 7.16564f
C1508 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 7.15659f
C1509 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 7.15659f
C1510 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 20.872599f
C1511 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 20.872599f
C1512 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 8.18273f
C1513 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 8.18273f
C1514 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 13.6417f
C1515 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 13.6417f
C1516 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 10.065901f
C1517 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 10.065901f
C1518 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 7.16564f
C1519 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 7.16564f
C1520 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 7.15659f
C1521 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 7.15659f
C1522 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 20.869598f
C1523 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 20.869598f
C1524 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 8.18273f
C1525 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 8.18273f
C1526 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 13.6439f
C1527 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 13.6439f
C1528 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 10.0691f
C1529 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 10.0719f
C1530 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.87363f
C1531 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.870339f
C1532 a_15390_2630# VGND 0.539466f $ **FLOATING
C1533 a_13950_2630# VGND 0.427094f $ **FLOATING
C1534 a_12582_2630# VGND 0.426679f $ **FLOATING
C1535 a_11142_2630# VGND 0.540621f $ **FLOATING
C1536 a_15390_2982# VGND 0.488855f $ **FLOATING
C1537 a_13950_2982# VGND 0.352472f $ **FLOATING
C1538 a_12582_2982# VGND 0.352472f $ **FLOATING
C1539 a_11142_2982# VGND 0.487284f $ **FLOATING
C1540 a_15390_3334# VGND 0.372888f $ **FLOATING
C1541 a_13950_3334# VGND 0.352438f $ **FLOATING
C1542 a_12582_3334# VGND 0.352438f $ **FLOATING
C1543 a_11142_3334# VGND 0.372888f $ **FLOATING
C1544 a_13950_3686# VGND 0.352418f $ **FLOATING
C1545 a_12582_3686# VGND 0.352418f $ **FLOATING
C1546 SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND 39.1318f
C1547 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.690451f
C1548 SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND 39.1318f
C1549 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.690451f
C1550 a_15390_4038# VGND 0.394414f $ **FLOATING
C1551 a_13950_4038# VGND 0.354407f $ **FLOATING
C1552 a_12582_4038# VGND 0.354407f $ **FLOATING
C1553 a_11142_4038# VGND 0.394414f $ **FLOATING
C1554 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VGND 36.5225f
C1555 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.33311f
C1556 a_13950_4390# VGND 0.352432f $ **FLOATING
C1557 a_12582_4390# VGND 0.352432f $ **FLOATING
C1558 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.33311f
C1559 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VGND 36.5225f
C1560 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VGND 2.95952f
C1561 a_15390_4566# VGND 0.38683f $ **FLOATING
C1562 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VGND 2.922f
C1563 a_11142_4566# VGND 0.38683f $ **FLOATING
C1564 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VGND 0.935058f
C1565 a_13950_4742# VGND 0.352456f $ **FLOATING
C1566 a_12582_4742# VGND 0.352456f $ **FLOATING
C1567 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND 0.78794f
C1568 a_15390_4918# VGND 0.467558f $ **FLOATING
C1569 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND 0.78794f
C1570 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VGND 0.935058f
C1571 a_11142_4918# VGND 0.469129f $ **FLOATING
C1572 a_13950_5094# VGND 0.353103f $ **FLOATING
C1573 a_12582_5094# VGND 0.353103f $ **FLOATING
C1574 a_15390_5270# VGND 0.490054f $ **FLOATING
C1575 a_11142_5270# VGND 0.488483f $ **FLOATING
C1576 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND 0.593399f
C1577 a_13950_5446# VGND 0.433341f $ **FLOATING
C1578 a_12582_5446# VGND 0.433756f $ **FLOATING
C1579 a_15390_5622# VGND 0.469507f $ **FLOATING
C1580 a_15390_5974# VGND 0.538415f $ **FLOATING
C1581 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND 0.593399f
C1582 a_11142_5622# VGND 0.471077f $ **FLOATING
C1583 a_11142_5974# VGND 0.53726f $ **FLOATING
C1584 a_22770_26796# VGND 0.52795f $ **FLOATING
C1585 a_21402_26796# VGND 0.530047f $ **FLOATING
C1586 a_17730_26796# VGND 0.529204f $ **FLOATING
C1587 a_16362_26796# VGND 0.53036f $ **FLOATING
C1588 a_12690_26796# VGND 0.529204f $ **FLOATING
C1589 a_11322_26796# VGND 0.53036f $ **FLOATING
C1590 a_7650_26796# VGND 0.528649f $ **FLOATING
C1591 a_6282_26796# VGND 0.529488f $ **FLOATING
C1592 a_2610_26796# VGND 0.529614f $ **FLOATING
C1593 a_22770_27148# VGND 0.497229f $ **FLOATING
C1594 a_21402_27148# VGND 0.465038f $ **FLOATING
C1595 a_17730_27148# VGND 0.468999f $ **FLOATING
C1596 a_16362_27148# VGND 0.465634f $ **FLOATING
C1597 a_12690_27148# VGND 0.468999f $ **FLOATING
C1598 a_11322_27148# VGND 0.465634f $ **FLOATING
C1599 a_7650_27148# VGND 0.467888f $ **FLOATING
C1600 a_6282_27148# VGND 0.463921f $ **FLOATING
C1601 a_2610_27148# VGND 0.468853f $ **FLOATING
C1602 a_21402_27500# VGND 0.383751f $ **FLOATING
C1603 a_17730_27500# VGND 0.385256f $ **FLOATING
C1604 a_16362_27500# VGND 0.384074f $ **FLOATING
C1605 a_12690_27500# VGND 0.385256f $ **FLOATING
C1606 a_11322_27500# VGND 0.384074f $ **FLOATING
C1607 a_7650_27500# VGND 0.384352f $ **FLOATING
C1608 a_6282_27500# VGND 0.382331f $ **FLOATING
C1609 a_2610_27500# VGND 0.385317f $ **FLOATING
C1610 a_21402_27852# VGND 0.367686f $ **FLOATING
C1611 a_17730_27852# VGND 0.368312f $ **FLOATING
C1612 a_16362_27852# VGND 0.366781f $ **FLOATING
C1613 a_12690_27852# VGND 0.368312f $ **FLOATING
C1614 a_11322_27852# VGND 0.366781f $ **FLOATING
C1615 a_7650_27852# VGND 0.367201f $ **FLOATING
C1616 a_6282_27852# VGND 0.365038f $ **FLOATING
C1617 a_2610_27852# VGND 0.368166f $ **FLOATING
C1618 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.D VGND 0.483793f
C1619 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.D VGND 0.480412f
C1620 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.D VGND 0.461451f
C1621 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.D VGND 0.480412f
C1622 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.D VGND 0.461451f
C1623 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.D VGND 0.480412f
C1624 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.D VGND 0.461451f
C1625 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.D VGND 0.480412f
C1626 a_21402_28204# VGND 0.402918f $ **FLOATING
C1627 a_17730_28204# VGND 0.403457f $ **FLOATING
C1628 a_16362_28204# VGND 0.403457f $ **FLOATING
C1629 a_12690_28204# VGND 0.403457f $ **FLOATING
C1630 a_11322_28204# VGND 0.403457f $ **FLOATING
C1631 a_7650_28204# VGND 0.402433f $ **FLOATING
C1632 a_6282_28204# VGND 0.401801f $ **FLOATING
C1633 a_2610_28204# VGND 0.403398f $ **FLOATING
C1634 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND 0.577116f
C1635 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN0.S VGND 0.734123f
C1636 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN0.S VGND 0.739788f
C1637 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN0.S VGND 0.729634f
C1638 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN0.S VGND 0.739788f
C1639 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN0.S VGND 0.729634f
C1640 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN0.S VGND 0.737472f
C1641 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN0.S VGND 0.725525f
C1642 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.S VGND 0.73983f
C1643 a_22770_28556# VGND 0.399356f $ **FLOATING
C1644 a_21402_28556# VGND 0.384985f $ **FLOATING
C1645 a_17730_28556# VGND 0.385524f $ **FLOATING
C1646 a_16362_28556# VGND 0.385524f $ **FLOATING
C1647 a_12690_28556# VGND 0.385524f $ **FLOATING
C1648 a_11322_28556# VGND 0.385524f $ **FLOATING
C1649 a_7650_28556# VGND 0.3845f $ **FLOATING
C1650 a_6282_28556# VGND 0.383868f $ **FLOATING
C1651 a_2610_28556# VGND 0.385465f $ **FLOATING
C1652 a_21402_28908# VGND 0.39155f $ **FLOATING
C1653 a_17730_28908# VGND 0.392089f $ **FLOATING
C1654 a_16362_28908# VGND 0.392089f $ **FLOATING
C1655 a_12690_28908# VGND 0.392089f $ **FLOATING
C1656 a_11322_28908# VGND 0.392089f $ **FLOATING
C1657 a_7650_28908# VGND 0.391065f $ **FLOATING
C1658 a_6282_28908# VGND 0.390433f $ **FLOATING
C1659 a_2610_28908# VGND 0.39203f $ **FLOATING
C1660 SUNSAR_SAR8B_CV_0.SARP VGND 0.143204p
C1661 a_21402_29612# VGND 0.393057f $ **FLOATING
C1662 a_17730_29612# VGND 0.393646f $ **FLOATING
C1663 a_16362_29612# VGND 0.393212f $ **FLOATING
C1664 a_12690_29612# VGND 0.393646f $ **FLOATING
C1665 a_11322_29612# VGND 0.393212f $ **FLOATING
C1666 a_7650_29612# VGND 0.392622f $ **FLOATING
C1667 a_6282_29612# VGND 0.391638f $ **FLOATING
C1668 a_2610_29612# VGND 0.393582f $ **FLOATING
C1669 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.299162f
C1670 a_22770_29964# VGND 0.398247f $ **FLOATING
C1671 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VGND 1.25305f
C1672 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VGND 1.24782f
C1673 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VGND 1.247f
C1674 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VGND 1.24782f
C1675 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VGND 1.247f
C1676 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VGND 1.24281f
C1677 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VGND 1.23805f
C1678 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VGND 1.2475f
C1679 a_21402_30316# VGND 0.399101f $ **FLOATING
C1680 a_17730_30316# VGND 0.398588f $ **FLOATING
C1681 a_16362_30316# VGND 0.398588f $ **FLOATING
C1682 a_12690_30316# VGND 0.398588f $ **FLOATING
C1683 a_11322_30316# VGND 0.398588f $ **FLOATING
C1684 a_7650_30316# VGND 0.397564f $ **FLOATING
C1685 a_6282_30316# VGND 0.396932f $ **FLOATING
C1686 a_2610_30316# VGND 0.398524f $ **FLOATING
C1687 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND 14.5848f
C1688 a_22770_30844# VGND 0.419082f $ **FLOATING
C1689 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND 2.22179f
C1690 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND 2.20473f
C1691 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND 2.20475f
C1692 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND 2.20473f
C1693 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND 2.20475f
C1694 SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND 2.19357f
C1695 SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND 2.18443f
C1696 SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND 2.20278f
C1697 a_21402_31196# VGND 0.422267f $ **FLOATING
C1698 a_17730_31196# VGND 0.422807f $ **FLOATING
C1699 a_16362_31196# VGND 0.422807f $ **FLOATING
C1700 a_12690_31196# VGND 0.422807f $ **FLOATING
C1701 a_11322_31196# VGND 0.422807f $ **FLOATING
C1702 a_7650_31196# VGND 0.421783f $ **FLOATING
C1703 a_6282_31196# VGND 0.421151f $ **FLOATING
C1704 a_2610_31196# VGND 0.422742f $ **FLOATING
C1705 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND 18.988f
C1706 a_22770_31724# VGND 0.420723f $ **FLOATING
C1707 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.95338f
C1708 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.93766f
C1709 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.93678f
C1710 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.93766f
C1711 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.93678f
C1712 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.34062f
C1713 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.010139f
C1714 a_21402_32076# VGND 0.422859f $ **FLOATING
C1715 a_17730_32076# VGND 0.423399f $ **FLOATING
C1716 a_16362_32076# VGND 0.423399f $ **FLOATING
C1717 a_12690_32076# VGND 0.423399f $ **FLOATING
C1718 a_11322_32076# VGND 0.423399f $ **FLOATING
C1719 a_7650_32076# VGND 0.423399f $ **FLOATING
C1720 a_6282_32076# VGND 0.423399f $ **FLOATING
C1721 a_2610_32076# VGND 0.423334f $ **FLOATING
C1722 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND 1.49316f
C1723 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.308787f
C1724 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND 3.10023f
C1725 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND 3.13373f
C1726 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND 3.13281f
C1727 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND 3.13373f
C1728 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND 3.13281f
C1729 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND 3.13084f
C1730 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND 3.12998f
C1731 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND 3.2189f
C1732 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND 2.66737f
C1733 a_21402_32956# VGND 0.422807f $ **FLOATING
C1734 a_17730_32956# VGND 0.422807f $ **FLOATING
C1735 a_16362_32956# VGND 0.422807f $ **FLOATING
C1736 a_12690_32956# VGND 0.422807f $ **FLOATING
C1737 a_11322_32956# VGND 0.422807f $ **FLOATING
C1738 a_7650_32956# VGND 0.422807f $ **FLOATING
C1739 a_6282_32956# VGND 0.422807f $ **FLOATING
C1740 a_2610_32956# VGND 0.422742f $ **FLOATING
C1741 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND 2.83208f
C1742 a_22770_33132# VGND 0.400772f $ **FLOATING
C1743 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 2.96363f
C1744 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 2.96825f
C1745 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 2.96834f
C1746 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 2.96825f
C1747 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 2.96834f
C1748 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.343029f
C1749 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.54721f
C1750 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 11.657901f
C1751 a_21402_33836# VGND 0.423443f $ **FLOATING
C1752 a_17730_33836# VGND 0.423443f $ **FLOATING
C1753 a_16362_33836# VGND 0.423443f $ **FLOATING
C1754 a_12690_33836# VGND 0.423443f $ **FLOATING
C1755 a_11322_33836# VGND 0.423443f $ **FLOATING
C1756 a_7650_33836# VGND 0.423443f $ **FLOATING
C1757 a_6282_33836# VGND 0.423443f $ **FLOATING
C1758 a_2610_33836# VGND 0.423291f $ **FLOATING
C1759 SUNSAR_SAR8B_CV_0.SARN VGND 0.144327p
C1760 SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.D VGND 0.146138f
C1761 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND 0.487114f
C1762 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.630399f
C1763 SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.D VGND 0.146138f
C1764 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.37303f
C1765 a_22770_34540# VGND 0.391469f $ **FLOATING
C1766 SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.D VGND 0.146138f
C1767 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 3.95932f
C1768 SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.D VGND 0.146138f
C1769 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.12911f
C1770 SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.D VGND 0.146138f
C1771 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.0789f
C1772 SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.D VGND 0.146138f
C1773 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.44242f
C1774 SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.D VGND 0.146138f
C1775 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 3.96126f
C1776 SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.D VGND 0.146138f
C1777 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 9.71945f
C1778 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 7.69803f
C1779 a_21402_34716# VGND 0.392167f $ **FLOATING
C1780 a_17730_34716# VGND 0.392167f $ **FLOATING
C1781 a_16362_34716# VGND 0.392167f $ **FLOATING
C1782 a_12690_34716# VGND 0.392167f $ **FLOATING
C1783 a_11322_34716# VGND 0.392167f $ **FLOATING
C1784 a_7650_34716# VGND 0.392167f $ **FLOATING
C1785 a_6282_34716# VGND 0.392167f $ **FLOATING
C1786 a_2610_34716# VGND 0.392102f $ **FLOATING
C1787 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND 4.73089f
C1788 a_22770_34892# VGND 0.391931f $ **FLOATING
C1789 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.65561f
C1790 SUNSAR_SAR8B_CV_0.XA6.ENO VGND 4.43303f
C1791 SUNSAR_SAR8B_CV_0.XA5.ENO VGND 4.33111f
C1792 SUNSAR_SAR8B_CV_0.XA4.ENO VGND 4.19979f
C1793 SUNSAR_SAR8B_CV_0.XA3.ENO VGND 4.37267f
C1794 SUNSAR_SAR8B_CV_0.XA2.ENO VGND 4.34942f
C1795 SUNSAR_SAR8B_CV_0.XA1.ENO VGND 4.31953f
C1796 SUNSAR_SAR8B_CV_0.XA0.ENO VGND 4.32115f
C1797 a_21402_35068# VGND 0.38696f $ **FLOATING
C1798 a_17730_35068# VGND 0.38696f $ **FLOATING
C1799 a_16362_35068# VGND 0.38696f $ **FLOATING
C1800 a_12690_35068# VGND 0.38696f $ **FLOATING
C1801 a_11322_35068# VGND 0.38696f $ **FLOATING
C1802 a_7650_35068# VGND 0.38696f $ **FLOATING
C1803 a_6282_35068# VGND 0.38696f $ **FLOATING
C1804 a_2610_35068# VGND 0.386896f $ **FLOATING
C1805 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND 4.48688f
C1806 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.531311f
C1807 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.520453f
C1808 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.531311f
C1809 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.520453f
C1810 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.531311f
C1811 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.520453f
C1812 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.542477f
C1813 a_22770_35420# VGND 0.392922f $ **FLOATING
C1814 a_21402_35420# VGND 0.386859f $ **FLOATING
C1815 a_17730_35420# VGND 0.386694f $ **FLOATING
C1816 a_16362_35420# VGND 0.387067f $ **FLOATING
C1817 a_12690_35420# VGND 0.386694f $ **FLOATING
C1818 a_11322_35420# VGND 0.387067f $ **FLOATING
C1819 a_7650_35420# VGND 0.386694f $ **FLOATING
C1820 a_6282_35420# VGND 0.387067f $ **FLOATING
C1821 a_2610_35420# VGND 0.386877f $ **FLOATING
C1822 SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND 1.05449f
C1823 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND 0.106067f
C1824 SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND 1.49344f
C1825 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VGND 1.48248f
C1826 SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND 1.4938f
C1827 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND 0.106067f
C1828 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VGND 1.48661f
C1829 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND 0.106067f
C1830 SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND 1.4942f
C1831 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VGND 1.47678f
C1832 SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND 1.4938f
C1833 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND 0.106067f
C1834 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VGND 1.48661f
C1835 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND 0.106067f
C1836 SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND 1.4942f
C1837 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VGND 1.47678f
C1838 SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND 1.4938f
C1839 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND 0.106067f
C1840 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VGND 1.48661f
C1841 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND 0.106067f
C1842 SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND 1.4942f
C1843 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VGND 1.47678f
C1844 SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND 1.50208f
C1845 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND 0.106067f
C1846 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VGND 1.55576f
C1847 a_22770_35948# VGND 0.411021f $ **FLOATING
C1848 a_21402_35948# VGND 0.388247f $ **FLOATING
C1849 a_17730_35948# VGND 0.388786f $ **FLOATING
C1850 a_16362_35948# VGND 0.388786f $ **FLOATING
C1851 a_12690_35948# VGND 0.388786f $ **FLOATING
C1852 a_11322_35948# VGND 0.388786f $ **FLOATING
C1853 a_7650_35948# VGND 0.388786f $ **FLOATING
C1854 a_6282_35948# VGND 0.388786f $ **FLOATING
C1855 a_2610_35948# VGND 0.388722f $ **FLOATING
C1856 SUNSAR_SAR8B_CV_0.XA20.XA10.B VGND 0.777474f
C1857 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.868472f
C1858 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.870095f
C1859 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.870155f
C1860 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.870095f
C1861 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.870155f
C1862 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.870095f
C1863 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.870155f
C1864 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.878758f
C1865 a_22770_36300# VGND 0.470018f $ **FLOATING
C1866 a_21402_36300# VGND 0.391211f $ **FLOATING
C1867 a_17730_36300# VGND 0.392024f $ **FLOATING
C1868 a_16362_36300# VGND 0.39175f $ **FLOATING
C1869 a_12690_36300# VGND 0.392004f $ **FLOATING
C1870 a_11322_36300# VGND 0.39175f $ **FLOATING
C1871 a_7650_36300# VGND 0.392002f $ **FLOATING
C1872 a_6282_36300# VGND 0.39175f $ **FLOATING
C1873 a_2610_36300# VGND 0.391937f $ **FLOATING
C1874 a_22770_36652# VGND 0.539269f $ **FLOATING
C1875 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND 0.867157f
C1876 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND 0.869383f
C1877 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND 0.862778f
C1878 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND 0.869362f
C1879 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND 0.862766f
C1880 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND 0.869361f
C1881 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND 0.862778f
C1882 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND 0.875877f
C1883 SUNSAR_SAR8B_CV_0.XA0.CEIN VGND 32.539497f
C1884 a_21402_36828# VGND 0.411129f $ **FLOATING
C1885 a_17730_36828# VGND 0.410959f $ **FLOATING
C1886 a_16362_36828# VGND 0.410719f $ **FLOATING
C1887 a_12690_36828# VGND 0.41095f $ **FLOATING
C1888 a_11322_36828# VGND 0.410718f $ **FLOATING
C1889 a_7650_36828# VGND 0.410952f $ **FLOATING
C1890 a_6282_36828# VGND 0.410719f $ **FLOATING
C1891 a_2610_36828# VGND 0.41074f $ **FLOATING
C1892 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND 1.07046f
C1893 SUNSAR_SAR8B_CV_0.XA7.CEO VGND 1.88576f
C1894 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND 1.08743f
C1895 SUNSAR_SAR8B_CV_0.XA6.CEO VGND 1.41392f
C1896 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND 1.05234f
C1897 SUNSAR_SAR8B_CV_0.XA5.CEO VGND 1.69845f
C1898 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND 1.08738f
C1899 SUNSAR_SAR8B_CV_0.XA4.CEO VGND 1.49292f
C1900 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND 1.05233f
C1901 SUNSAR_SAR8B_CV_0.XA3.CEO VGND 1.69844f
C1902 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND 1.08739f
C1903 SUNSAR_SAR8B_CV_0.XA2.CEO VGND 1.49293f
C1904 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND 1.05234f
C1905 SUNSAR_SAR8B_CV_0.XA1.CEO VGND 1.69844f
C1906 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND 1.09608f
C1907 SUNSAR_SAR8B_CV_0.XA0.CEO VGND 1.4987f
C1908 a_21402_37180# VGND 0.472605f $ **FLOATING
C1909 a_17730_37180# VGND 0.471966f $ **FLOATING
C1910 a_16362_37180# VGND 0.473517f $ **FLOATING
C1911 a_12690_37180# VGND 0.471951f $ **FLOATING
C1912 a_11322_37180# VGND 0.473516f $ **FLOATING
C1913 a_7650_37180# VGND 0.471954f $ **FLOATING
C1914 a_6282_37180# VGND 0.473517f $ **FLOATING
C1915 a_2610_37180# VGND 0.47159f $ **FLOATING
C1916 a_21402_37532# VGND 0.543507f $ **FLOATING
C1917 a_17730_37532# VGND 0.545679f $ **FLOATING
C1918 a_16362_37532# VGND 0.544363f $ **FLOATING
C1919 a_12690_37532# VGND 0.545542f $ **FLOATING
C1920 a_11322_37532# VGND 0.544363f $ **FLOATING
C1921 a_7650_37532# VGND 0.545576f $ **FLOATING
C1922 a_6282_37532# VGND 0.544365f $ **FLOATING
C1923 a_2610_37532# VGND 0.543853f $ **FLOATING
C1924 a_22790_40296# VGND 0.543886f $ **FLOATING
C1925 a_21422_40296# VGND 0.543054f $ **FLOATING
C1926 a_17750_40296# VGND 0.544048f $ **FLOATING
C1927 a_16382_40296# VGND 0.545201f $ **FLOATING
C1928 a_12710_40296# VGND 0.544048f $ **FLOATING
C1929 a_11342_40296# VGND 0.545204f $ **FLOATING
C1930 a_7670_40296# VGND 0.544046f $ **FLOATING
C1931 a_6302_40296# VGND 0.545201f $ **FLOATING
C1932 a_2630_40296# VGND 0.542813f $ **FLOATING
C1933 a_22790_40648# VGND 0.489516f $ **FLOATING
C1934 a_21422_40648# VGND 0.48751f $ **FLOATING
C1935 a_17750_40648# VGND 0.489596f $ **FLOATING
C1936 a_16382_40648# VGND 0.488025f $ **FLOATING
C1937 a_12710_40648# VGND 0.489596f $ **FLOATING
C1938 a_11342_40648# VGND 0.488025f $ **FLOATING
C1939 a_7670_40648# VGND 0.489596f $ **FLOATING
C1940 a_6302_40648# VGND 0.488025f $ **FLOATING
C1941 a_2630_40648# VGND 0.489995f $ **FLOATING
C1942 SUNSAR_SAR8B_CV_0.DONE VGND 20.345901f
C1943 a_22790_41000# VGND 0.386169f $ **FLOATING
C1944 a_21422_41000# VGND 0.385655f $ **FLOATING
C1945 a_17750_41000# VGND 0.385655f $ **FLOATING
C1946 a_16382_41000# VGND 0.385655f $ **FLOATING
C1947 a_12710_41000# VGND 0.385655f $ **FLOATING
C1948 a_11342_41000# VGND 0.385655f $ **FLOATING
C1949 a_7670_41000# VGND 0.385655f $ **FLOATING
C1950 a_6302_41000# VGND 0.385655f $ **FLOATING
C1951 a_2630_41000# VGND 0.386141f $ **FLOATING
C1952 a_22790_41352# VGND 0.372123f $ **FLOATING
C1953 a_21422_41352# VGND 0.390928f $ **FLOATING
C1954 a_17750_41352# VGND 0.390928f $ **FLOATING
C1955 a_16382_41352# VGND 0.390928f $ **FLOATING
C1956 a_12710_41352# VGND 0.390928f $ **FLOATING
C1957 a_11342_41352# VGND 0.390928f $ **FLOATING
C1958 a_7670_41352# VGND 0.390928f $ **FLOATING
C1959 a_6302_41352# VGND 0.390928f $ **FLOATING
C1960 a_2630_41352# VGND 0.391414f $ **FLOATING
C1961 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND 0.792386f
C1962 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND 0.100913f
C1963 SUNSAR_SAR8B_CV_0.D<0> VGND 5.62991f
C1964 SUNSAR_SAR8B_CV_0.D<1> VGND 13.1194f
C1965 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND 0.100821f
C1966 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND 0.100821f
C1967 SUNSAR_SAR8B_CV_0.D<2> VGND 12.0092f
C1968 SUNSAR_SAR8B_CV_0.D<3> VGND 10.9751f
C1969 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND 0.100821f
C1970 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND 0.100821f
C1971 SUNSAR_SAR8B_CV_0.D<4> VGND 11.348901f
C1972 SUNSAR_SAR8B_CV_0.D<5> VGND 12.1097f
C1973 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND 0.100821f
C1974 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND 0.100821f
C1975 SUNSAR_SAR8B_CV_0.D<6> VGND 11.5195f
C1976 SUNSAR_SAR8B_CV_0.D<7> VGND 16.6604f
C1977 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND 0.100821f
C1978 a_22790_41880# VGND 0.39234f $ **FLOATING
C1979 a_21422_41880# VGND 0.392571f $ **FLOATING
C1980 a_17750_41880# VGND 0.393111f $ **FLOATING
C1981 a_16382_41880# VGND 0.393111f $ **FLOATING
C1982 a_12710_41880# VGND 0.393111f $ **FLOATING
C1983 a_11342_41880# VGND 0.393111f $ **FLOATING
C1984 a_7670_41880# VGND 0.393111f $ **FLOATING
C1985 a_6302_41880# VGND 0.393111f $ **FLOATING
C1986 a_2630_41880# VGND 0.393486f $ **FLOATING
C1987 SUNSAR_CAPT8B_CV_0.XA3.A VGND 1.91068f
C1988 a_22790_42408# VGND 0.408132f $ **FLOATING
C1989 a_21422_42408# VGND 0.387221f $ **FLOATING
C1990 a_17750_42408# VGND 0.387761f $ **FLOATING
C1991 a_16382_42408# VGND 0.387761f $ **FLOATING
C1992 a_12710_42408# VGND 0.387761f $ **FLOATING
C1993 a_11342_42408# VGND 0.387761f $ **FLOATING
C1994 a_7670_42408# VGND 0.387761f $ **FLOATING
C1995 a_6302_42408# VGND 0.387761f $ **FLOATING
C1996 a_2630_42408# VGND 0.388136f $ **FLOATING
C1997 SUNSAR_CAPT8B_CV_0.XA5.XA1.Y VGND 1.01852f
C1998 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND 1.24489f
C1999 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND 1.23659f
C2000 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND 1.23659f
C2001 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND 1.23659f
C2002 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND 1.23659f
C2003 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND 1.23659f
C2004 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND 1.23659f
C2005 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND 1.2531f
C2006 a_22790_42760# VGND 0.376791f $ **FLOATING
C2007 a_21422_42760# VGND 0.390424f $ **FLOATING
C2008 a_17750_42760# VGND 0.390963f $ **FLOATING
C2009 a_16382_42760# VGND 0.390963f $ **FLOATING
C2010 a_12710_42760# VGND 0.390963f $ **FLOATING
C2011 a_11342_42760# VGND 0.390963f $ **FLOATING
C2012 a_7670_42760# VGND 0.390963f $ **FLOATING
C2013 a_6302_42760# VGND 0.390963f $ **FLOATING
C2014 a_2630_42760# VGND 0.391339f $ **FLOATING
C2015 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 23.963099f
C2016 SUNSAR_SAR8B_CV_0.EN VGND 10.3178f
C2017 a_22790_43112# VGND 0.38655f $ **FLOATING
C2018 SUNSAR_CAPT8B_CV_0.XI14.XA5.Y VGND 1.27898f
C2019 SUNSAR_CAPT8B_CV_0.XH13.XA5.Y VGND 1.28097f
C2020 SUNSAR_CAPT8B_CV_0.XG12.XA5.Y VGND 1.28097f
C2021 SUNSAR_CAPT8B_CV_0.XF11.XA5.Y VGND 1.28097f
C2022 SUNSAR_CAPT8B_CV_0.XE10.XA5.Y VGND 1.28097f
C2023 SUNSAR_CAPT8B_CV_0.XD09.XA5.Y VGND 1.28097f
C2024 SUNSAR_CAPT8B_CV_0.XC08.XA5.Y VGND 1.28097f
C2025 SUNSAR_CAPT8B_CV_0.XB07.XA5.Y VGND 1.28345f
C2026 SUNSAR_CAPT8B_CV_0.XA5.A VGND 2.23979f
C2027 a_21422_43288# VGND 0.391671f $ **FLOATING
C2028 a_17750_43288# VGND 0.392211f $ **FLOATING
C2029 a_16382_43288# VGND 0.392211f $ **FLOATING
C2030 a_12710_43288# VGND 0.392211f $ **FLOATING
C2031 a_11342_43288# VGND 0.392211f $ **FLOATING
C2032 a_7670_43288# VGND 0.392211f $ **FLOATING
C2033 a_6302_43288# VGND 0.392211f $ **FLOATING
C2034 a_2630_43288# VGND 0.392586f $ **FLOATING
C2035 SUNSAR_CAPT8B_CV_0.XA3.Y VGND 1.59466f
C2036 a_22790_43640# VGND 0.385751f $ **FLOATING
C2037 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND 0.106067f
C2038 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND 2.57238f
C2039 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VGND 1.67006f
C2040 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND 0.106067f
C2041 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VGND 1.67243f
C2042 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND 2.555f
C2043 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND 0.106067f
C2044 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND 2.55514f
C2045 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VGND 1.67243f
C2046 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND 0.106067f
C2047 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VGND 1.67243f
C2048 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND 2.555f
C2049 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND 0.106067f
C2050 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND 2.55514f
C2051 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VGND 1.67243f
C2052 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND 0.106067f
C2053 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VGND 1.67243f
C2054 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND 2.555f
C2055 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND 0.106067f
C2056 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND 2.55514f
C2057 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VGND 1.67243f
C2058 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND 0.106067f
C2059 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VGND 1.67194f
C2060 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND 2.62109f
C2061 SUNSAR_CAPT8B_CV_0.XA6.XA1.Y VGND 0.948554f
C2062 a_21422_43816# VGND 0.38804f $ **FLOATING
C2063 a_17750_43816# VGND 0.388579f $ **FLOATING
C2064 a_16382_43816# VGND 0.388579f $ **FLOATING
C2065 a_12710_43816# VGND 0.388579f $ **FLOATING
C2066 a_11342_43816# VGND 0.388579f $ **FLOATING
C2067 a_7670_43816# VGND 0.388579f $ **FLOATING
C2068 a_6302_43816# VGND 0.388579f $ **FLOATING
C2069 a_2630_43816# VGND 0.388955f $ **FLOATING
C2070 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 24.5001f
C2071 a_22790_43992# VGND 0.424176f $ **FLOATING
C2072 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.2375f
C2073 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.23686f
C2074 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.23686f
C2075 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.23686f
C2076 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.23686f
C2077 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.23686f
C2078 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.23686f
C2079 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.23702f
C2080 a_21422_44168# VGND 0.424488f $ **FLOATING
C2081 a_17750_44168# VGND 0.423472f $ **FLOATING
C2082 a_16382_44168# VGND 0.423887f $ **FLOATING
C2083 a_12710_44168# VGND 0.423472f $ **FLOATING
C2084 a_11342_44168# VGND 0.423887f $ **FLOATING
C2085 a_7670_44168# VGND 0.423472f $ **FLOATING
C2086 a_6302_44168# VGND 0.423887f $ **FLOATING
C2087 a_2630_44168# VGND 0.424073f $ **FLOATING
.ends

