* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

.subckt SUNTR_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 B G 0.33939f
C1 a_216_n18# B 0.330729f
C2 a_216_334# B 0.331144f
C3 B VSUBS 2.80592f
.ends

.subckt SUNTR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 G B 0.411913f
C1 a_324_n18# B 0.422415f
C2 a_324_334# B 0.422f
.ends

.subckt SUNTR_BFX1_CV Y AVDD AVSS MP1/B MN1/a_324_334# A MP1/a_216_334# VSUBS
XMP0 AVDD A MP1/G MP1/B MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNTR_PCHDL
XMP1 Y MP1/G AVDD MP1/B MP1/a_216_n18# MP1/a_216_334# VSUBS SUNTR_PCHDL
XMN0 AVSS A MP1/G VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNTR_NCHDL
XMN1 Y MP1/G AVSS VSUBS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 MP1/B MP1/a_216_n18# -0.310513f
C1 AVSS AVDD 0.10499f
C2 MP1/G AVSS 0.120067f
C3 A MP1/G 0.156853f
C4 MP1/B AVDD 0.181063f
C5 MP1/B MP1/G 0.178777f
C6 MP1/B A 0.109691f
C7 AVDD VSUBS 0.276075f
C8 AVSS VSUBS 0.45436f
C9 Y VSUBS 0.218882f
C10 MN1/a_324_n18# VSUBS 0.351938f
C11 MN1/a_324_334# VSUBS 0.422f
C12 MP1/G VSUBS 0.969276f
C13 A VSUBS 0.55997f
C14 MN0/a_324_n18# VSUBS 0.422415f
C15 MP1/B VSUBS 4.386796f
.ends

.subckt SUNTR_TIEH_CV Y AVDD AVSS MP0/B MP0/G MP0/a_216_334# MP0/a_216_n18# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y MP0/G AVDD MP0/B MP0/a_216_n18# MP0/a_216_334# VSUBS SUNTR_PCHDL
XMN0 MP0/G MP0/G AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNTR_NCHDL
C0 MP0/B MP0/G 0.112479f
C1 MP0/B AVDD 0.112171f
C2 AVDD VSUBS 0.260853f
C3 AVSS VSUBS 0.382267f
C4 MP0/G VSUBS 0.78444f
C5 MN0/a_324_n18# VSUBS 0.422415f
C6 MN0/a_324_334# VSUBS 0.422f
C7 MP0/B VSUBS 2.80738f
.ends

.subckt SUNTR_TAPCELLB_CV AVDD MN1/a_324_n18# MP1/a_216_n18# AVSS
XMP1 AVDD AVDD AVDD AVDD MP1/a_216_n18# MP1/a_216_334# AVSS SUNTR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 AVDD AVSS 0.107602f
C1 AVSS 0 1.064147f
C2 MN1/a_324_n18# 0 0.422415f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.146627f
.ends

.subckt tt_um_TT06_SAR_done DONE uio_out<0> uio_oe<0> VPWR VGND
Xx3 uio_out<0> VPWR VGND VPWR x4/MN0/a_324_n18# DONE x4/MP0/a_216_n18# VGND SUNTR_BFX1_CV
Xx4 uio_oe<0> VPWR VGND VPWR x4/MP0/G x5/MP1/a_216_n18# x4/MP0/a_216_n18# x4/MN0/a_324_n18#
+ VGND x5/MN1/a_324_n18# SUNTR_TIEH_CV
Xx5 VPWR x5/MN1/a_324_n18# x5/MP1/a_216_n18# VGND SUNTR_TAPCELLB_CV
C0 uio_oe<0> VPWR 0.524617f
C1 uio_out<0> VGND 0.294473f
C2 x4/MP0/G VGND 0.114893f
C3 VPWR x5/MP1/a_216_n18# -0.314359f
C4 x4/MP0/a_216_n18# VPWR -0.31151f
C5 VGND 0 0.898244f
C6 x5/MN1/a_324_334# 0 0.422f
C7 VPWR 0 7.717914f
C8 x4/MP0/G 0 0.782647f
C9 x5/MN1/a_324_n18# 0 0.360407f
C10 uio_oe<0> 0 0.133144f
C11 uio_out<0> 0 0.357519f
C12 x3/MN1/a_324_n18# 0 0.355196f
C13 x4/MN0/a_324_n18# 0 0.360407f
C14 x3/MP1/G 0 0.95314f
C15 DONE 0 0.720744f
C16 x3/MN0/a_324_n18# 0 0.422415f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_XS736D c1_n1946_n17480# m3_n1986_n17520# VSUBS
X0 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X1 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X2 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X3 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X4 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X5 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X6 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X7 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X8 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
C0 m3_n1986_n17520# c1_n1946_n17480# 0.265161p
C1 c1_n1946_n17480# VSUBS 9.109429f
C2 m3_n1986_n17520# VSUBS 65.3375f
.ends

.subckt SUNSAR_RM1 A B VSUBS
R0 A B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
.ends

.subckt SUNSAR_CAP32C_CV C1B C2 C4 C16 CTOP AVSS C1A XRES1A/B C8 XRES1B/B VSUBS
XXRES16 C16 XRES16/B VSUBS SUNSAR_RM1
XXRES2 C2 XRES2/B VSUBS SUNSAR_RM1
XXRES1A C1A XRES1A/B VSUBS SUNSAR_RM1
XXRES4 C4 XRES4/B VSUBS SUNSAR_RM1
XXRES1B C1B XRES1B/B VSUBS SUNSAR_RM1
XXRES8 C8 XRES8/B VSUBS SUNSAR_RM1
C0 XRES1A/B XRES16/B 0.437694f
C1 XRES1A/B AVSS 3.7558f
C2 XRES1B/B CTOP 3.552515f
C3 XRES8/B XRES2/B 0.419738f
C4 XRES8/B XRES4/B 0.449585f
C5 XRES16/B XRES2/B 0.441867f
C6 AVSS XRES2/B 4.083764f
C7 AVSS XRES4/B 4.927044f
C8 XRES1A/B CTOP 3.552515f
C9 AVSS XRES8/B 6.54197f
C10 AVSS XRES16/B 9.801106f
C11 XRES1B/B XRES4/B 0.40569f
C12 XRES2/B CTOP 6.866754f
C13 XRES1B/B AVSS 3.75982f
C14 XRES4/B CTOP 13.651895f
C15 XRES8/B CTOP 27.161474f
C16 XRES16/B CTOP 54.216488f
C17 AVSS CTOP 9.918658f
C18 CTOP VSUBS 7.76011f
C19 XRES2/B VSUBS 3.1129f
C20 XRES4/B VSUBS 3.516117f
C21 XRES8/B VSUBS 3.933522f
C22 XRES16/B VSUBS 4.664508f
C23 AVSS VSUBS 15.179144f
C24 C8 VSUBS 0.101745f
C25 XRES1B/B VSUBS 2.892833f
C26 C1B VSUBS 0.116997f
C27 C4 VSUBS 0.101745f
C28 XRES1A/B VSUBS 1.735354f
C29 C1A VSUBS 0.116997f
C30 C2 VSUBS 0.101745f
C31 C16 VSUBS 0.101745f
.ends

.subckt SUNSAR_CDAC7_CV CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0>
+ CTOP AVSS VSUBS
XX16ab CP<5> CP<5> CP<5> CP<6> CTOP AVSS CP<5> X16ab/XRES1A/B CP<4> X16ab/XRES1B/B
+ VSUBS SUNSAR_CAP32C_CV
XXC0 CP<9> CP<9> CP<9> CP<9> CTOP AVSS CP<9> XC0/XRES1A/B CP<9> XC0/XRES1B/B VSUBS
+ SUNSAR_CAP32C_CV
XXC1 CP<8> CP<8> CP<8> CP<8> CTOP AVSS CP<8> XC1/XRES1A/B CP<8> XC1/XRES1B/B VSUBS
+ SUNSAR_CAP32C_CV
XXC32a<0> CP<0> CP<1> CP<2> CP<7> CTOP AVSS AVSS XC32a<0>/XRES1A/B CP<3> XC32a<0>/XRES1B/B
+ VSUBS SUNSAR_CAP32C_CV
C0 CP<1> CP<3> 0.220707f
C1 CP<9> CP<5> 0.103206f
C2 XC1/XRES1B/B XC32a<0>/XRES1A/B 0.635098f
C3 X16ab/XRES1B/B XC0/XRES1A/B 0.635098f
C4 AVSS CTOP -1.633715f
C5 CP<5> CP<0> 0.20259f
C6 CP<7> CP<8> 2.575701f
C7 CP<8> CTOP 0.122672f
C8 CP<5> CP<8> 0.359484f
C9 CP<2> CP<3> 2.212231f
C10 CP<0> CP<1> 1.909476f
C11 X16ab/XRES1A/B XC32a<0>/XRES1B/B 0.635098f
C12 CP<2> CP<1> 1.995553f
C13 CP<5> CP<4> 1.57931f
C14 CP<5> CP<7> 0.394951f
C15 CP<9> AVSS 0.343312f
C16 CP<4> CP<3> 1.263888f
C17 CP<3> CP<7> 0.178438f
C18 CP<6> CP<7> 1.652261f
C19 CP<5> CP<3> 0.229397f
C20 CP<9> CP<8> 0.889573f
C21 CP<6> CP<5> 2.020583f
C22 CP<2> CP<0> 0.24075f
C23 CP<1> CP<7> 0.188755f
C24 CP<8> AVSS 0.71211f
C25 XC32a<0>/XRES2/B VSUBS 3.1129f
C26 XC32a<0>/XRES4/B VSUBS 3.516117f
C27 XC32a<0>/XRES8/B VSUBS 3.933522f
C28 XC32a<0>/XRES16/B VSUBS 4.664508f
C29 CP<3> VSUBS 1.126461f
C30 XC32a<0>/XRES1B/B VSUBS 2.892833f
C31 CP<0> VSUBS 1.167979f
C32 CP<2> VSUBS 0.834649f
C33 XC32a<0>/XRES1A/B VSUBS 1.735354f
C34 CP<1> VSUBS 1.392542f
C35 CP<7> VSUBS 1.060384f
C36 CTOP VSUBS 20.24516f
C37 XC1/XRES2/B VSUBS 3.1129f
C38 XC1/XRES4/B VSUBS 3.516117f
C39 XC1/XRES8/B VSUBS 3.933522f
C40 XC1/XRES16/B VSUBS 4.664508f
C41 AVSS VSUBS 51.996902f
C42 XC1/XRES1B/B VSUBS 2.892833f
C43 XC1/XRES1A/B VSUBS 1.735354f
C44 CP<8> VSUBS 3.823549f
C45 XC0/XRES2/B VSUBS 3.1129f
C46 XC0/XRES4/B VSUBS 3.516117f
C47 XC0/XRES8/B VSUBS 3.933522f
C48 XC0/XRES16/B VSUBS 4.664508f
C49 XC0/XRES1B/B VSUBS 2.892833f
C50 XC0/XRES1A/B VSUBS 1.735354f
C51 CP<5> VSUBS 2.378288f
C52 X16ab/XRES2/B VSUBS 3.1129f
C53 X16ab/XRES4/B VSUBS 3.516117f
C54 X16ab/XRES8/B VSUBS 3.933522f
C55 X16ab/XRES16/B VSUBS 4.664508f
C56 CP<4> VSUBS 0.757332f
C57 X16ab/XRES1B/B VSUBS 2.892833f
C58 X16ab/XRES1A/B VSUBS 1.735354f
C59 CP<6> VSUBS 0.645761f
C60 CP<9> VSUBS 2.290488f
.ends

.subckt SUNSAR_PCHDL D G S B a_216_n18# a_216_334# VSUBS
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 B G 0.341895f
C1 a_216_n18# B 0.330729f
C2 a_216_334# B 0.331144f
C3 B VSUBS 2.80584f
.ends

.subckt SUNSAR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 G B 0.415197f
C1 a_324_n18# B 0.422415f
C2 a_324_334# B 0.422f
.ends

.subckt SUNSAR_NDX1_CV Y AVDD AVSS MN1/a_324_334# B A BULKP MP0/a_216_n18# MP1/a_216_334#
+ MN0/a_324_n18# VSUBS
XMP0 Y A AVDD BULKP MP0/a_216_n18# B VSUBS SUNSAR_PCHDL
XMP1 AVDD B Y BULKP A MP1/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 Y B MN1/S VSUBS A MN1/a_324_334# SUNSAR_NCHDL
C0 A BULKP -0.246413f
C1 BULKP AVDD 0.154562f
C2 BULKP B -0.247362f
C3 AVSS VSUBS 0.392705f
C4 MN1/a_324_334# VSUBS 0.422f
C5 AVDD VSUBS 0.326781f
C6 MN0/a_324_n18# VSUBS 0.422415f
C7 Y VSUBS 0.252959f
C8 B VSUBS 0.538314f
C9 BULKP VSUBS 3.595964f
C10 A VSUBS 0.539194f
.ends

.subckt SUNSAR_NRX1_CV AVDD AVSS MN1/a_324_334# B BULKP MP0/a_216_n18# Y MP1/a_216_334#
+ A MN0/a_324_n18# VSUBS
XMP0 MP1/S A AVDD BULKP MP0/a_216_n18# B VSUBS SUNSAR_PCHDL
XMP1 Y B MP1/S BULKP A MP1/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 AVSS B Y VSUBS A MN1/a_324_334# SUNSAR_NCHDL
C0 A BULKP -0.246413f
C1 Y AVSS 0.112939f
C2 BULKP AVDD 0.122023f
C3 BULKP B -0.247362f
C4 AVSS VSUBS 0.506278f
C5 Y VSUBS 0.247181f
C6 MN1/a_324_334# VSUBS 0.422f
C7 MN0/a_324_n18# VSUBS 0.422415f
C8 AVDD VSUBS 0.25764f
C9 B VSUBS 0.538314f
C10 BULKP VSUBS 3.595964f
C11 A VSUBS 0.539194f
.ends

.subckt SUNSAR_IVX1_CV BULKP AVSS Y MP0/a_216_n18# MP0/a_216_334# AVDD A MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y A AVDD BULKP MP0/a_216_n18# MP0/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP A 0.109299f
C1 BULKP AVDD 0.103136f
C2 AVSS VSUBS 0.367376f
C3 A VSUBS 0.631634f
C4 Y VSUBS 0.268384f
C5 MN0/a_324_n18# VSUBS 0.422415f
C6 MN0/a_324_334# VSUBS 0.422f
C7 AVDD VSUBS 0.246592f
C8 BULKP VSUBS 2.80697f
.ends

.subckt SUNSAR_TAPCELLB_CV AVDD MN1/a_324_n18# MN1/a_324_334# MP1/a_216_334# MP1/a_216_n18#
+ AVSS
XMP1 AVDD AVDD AVDD AVDD MP1/a_216_n18# MP1/a_216_334# AVSS SUNSAR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.104949f
C1 AVSS 0 1.048908f
C2 MN1/a_324_n18# 0 0.422415f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.134387f
.ends

.subckt SUNSAR_SARKICKHX1_CV CI BULKP AVDD AVSS MP6_DMY/a_216_334# MN6/a_324_334#
+ CKN MP0/a_216_n18# CK MN0/a_324_n18# VSUBS
XMP1_DMY AVDD AVDD AVDD BULKP CKN AVDD VSUBS SUNSAR_PCHDL
XMP4_DMY AVDD AVDD AVDD BULKP AVDD AVDD VSUBS SUNSAR_PCHDL
XMP0 AVDD CKN MP0/S BULKP MP0/a_216_n18# AVDD VSUBS SUNSAR_PCHDL
XMN0 MP0/S CKN AVSS VSUBS MN0/a_324_n18# CI SUNSAR_NCHDL
XMN1 MP0/S CI MP0/S VSUBS CKN CI SUNSAR_NCHDL
XMN2 MP0/S CI MP0/S VSUBS CI CI SUNSAR_NCHDL
XMN3 MP0/S CI MP0/S VSUBS CI CI SUNSAR_NCHDL
XMN4 MP0/S CI MP0/S VSUBS CI CI SUNSAR_NCHDL
XMN6 AVDD CK MP0/S VSUBS CI MN6/a_324_334# SUNSAR_NCHDL
XMN5 MP0/S CI MP0/S VSUBS CI CK SUNSAR_NCHDL
XMP3_DMY AVDD AVDD AVDD BULKP AVDD AVDD VSUBS SUNSAR_PCHDL
XMP6_DMY AVDD AVDD AVDD BULKP AVDD MP6_DMY/a_216_334# VSUBS SUNSAR_PCHDL
XMP2_DMY AVDD AVDD AVDD BULKP AVDD AVDD VSUBS SUNSAR_PCHDL
XMP5_DMY AVDD AVDD AVDD BULKP AVDD AVDD VSUBS SUNSAR_PCHDL
C0 CKN BULKP -0.227092f
C1 BULKP AVDD -3.515122f
C2 MP0/S AVSS 0.208328f
C3 AVSS AVDD 0.180248f
C4 MP0/S AVDD 0.104608f
C5 MP0/S BULKP 0.11694f
C6 AVDD VSUBS 0.74157f
C7 BULKP VSUBS 7.544365f
C8 CK VSUBS 0.372036f
C9 MN6/a_324_334# VSUBS 0.422f
C10 CI VSUBS 1.791641f
C11 AVSS VSUBS 0.555322f
C12 MN0/a_324_n18# VSUBS 0.422415f
C13 MP0/S VSUBS 0.370985f
C14 CKN VSUBS 0.56349f
.ends

.subckt SUNSAR_SARCMPHX1_CV CI CK VMR N2 AVDD AVSS MP6/a_216_334# MN6/a_324_334# BULKP
+ MP0/a_216_n18# CO MN0/a_324_n18# VSUBS N1
XMP0 AVDD CK N1 BULKP MP0/a_216_n18# CK VSUBS SUNSAR_PCHDL
XMP1 N2 CK AVDD BULKP CK AVDD VSUBS SUNSAR_PCHDL
XMN0 N1 CK AVSS VSUBS MN0/a_324_n18# CI SUNSAR_NCHDL
XMP2 AVDD AVDD N2 BULKP CK CK VSUBS SUNSAR_PCHDL
XMN1 N2 CI N1 VSUBS CK CI SUNSAR_NCHDL
XMP3 CO CK AVDD BULKP AVDD VMR VSUBS SUNSAR_PCHDL
XMP4 AVDD VMR CO BULKP CK VMR VSUBS SUNSAR_PCHDL
XMN2 N1 CI N2 VSUBS CI CI SUNSAR_NCHDL
XMP5 CO VMR AVDD BULKP VMR VMR VSUBS SUNSAR_PCHDL
XMN3 N2 CI N1 VSUBS CI CI SUNSAR_NCHDL
XMN4 N1 CI N2 VSUBS CI CI SUNSAR_NCHDL
XMP6 AVDD VMR CO BULKP VMR MP6/a_216_334# VSUBS SUNSAR_PCHDL
XMN5 N2 CI N1 VSUBS CI VMR SUNSAR_NCHDL
XMN6 CO VMR N2 VSUBS CI MN6/a_324_334# SUNSAR_NCHDL
C0 BULKP CK -1.349649f
C1 N1 CI 0.175052f
C2 BULKP VMR -1.552184f
C3 AVDD CO 0.222193f
C4 AVDD BULKP -0.442314f
C5 AVDD AVSS 0.157463f
C6 N1 AVSS 0.158948f
C7 N1 N2 0.189549f
C8 AVSS VSUBS 0.533831f
C9 MN6/a_324_334# VSUBS 0.422f
C10 VMR VSUBS 0.606867f
C11 CI VSUBS 1.771056f
C12 CK VSUBS 0.626869f
C13 CO VSUBS 0.213838f
C14 BULKP VSUBS 7.544966f
C15 N2 VSUBS 0.221339f
C16 MN0/a_324_n18# VSUBS 0.422415f
C17 AVDD VSUBS 0.609607f
C18 N1 VSUBS 0.369132f
.ends

.subckt SUNSAR_IVX4_CV AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18#
+ Y A MN0/a_324_n18# VSUBS
XMP0 Y A AVDD BULKP MP0/a_216_n18# A VSUBS SUNSAR_PCHDL
XMP1 AVDD A Y BULKP A A VSUBS SUNSAR_PCHDL
XMP2 Y A AVDD BULKP A A VSUBS SUNSAR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 AVDD A Y BULKP A MP3/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 AVSS A Y VSUBS A A SUNSAR_NCHDL
XMN2 Y A AVSS VSUBS A A SUNSAR_NCHDL
XMN3 AVSS A Y VSUBS A MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.166303f
C1 Y AVSS 0.174863f
C2 BULKP A -1.606473f
C3 AVDD AVSS 0.131604f
C4 AVDD Y 0.146264f
C5 Y A 0.147008f
C6 A VSUBS 2.062361f
C7 AVSS VSUBS 0.622587f
C8 MN3/a_324_334# VSUBS 0.422f
C9 Y VSUBS 0.278637f
C10 MN0/a_324_n18# VSUBS 0.422415f
C11 AVDD VSUBS 0.372455f
C12 BULKP VSUBS 5.176431f
.ends

.subckt SUNSAR_SARCMPX1_CV CPI CNI CK_CMP CK_SAMPLE DONE XA9/A CPO AVDD CNO AVSS
XXA10 XA9/A AVDD AVSS XA11/MN0/a_324_n18# XA12/Y XA11/Y AVDD XA9/MP0/a_216_334# XA11/MP0/a_216_n18#
+ XA9/MN0/a_324_334# AVSS SUNSAR_NDX1_CV
XXA11 AVDD AVSS XA12/MN0/a_324_n18# DONE AVDD XA11/MP0/a_216_n18# XA11/Y XA12/MP0/a_216_n18#
+ CK_SAMPLE XA11/MN0/a_324_n18# AVSS SUNSAR_NRX1_CV
XXA12 AVDD AVSS XA12/Y XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD CK_CMP XA12/MN0/a_324_n18#
+ AVSS XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVDD XA13/MN1/a_324_n18# XA13/MN1/a_324_334# XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA1 CPI AVDD AVDD AVSS XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# XA9/A XA1/MP0/a_216_n18#
+ XA9/Y XA1/MN0/a_324_n18# AVSS SUNSAR_SARKICKHX1_CV
XXA2 CPI XA9/Y XA3/CO XA2/N2 AVDD AVSS XA2/MP6/a_216_334# XA2/MN6/a_324_334# AVDD
+ XA2/MP0/a_216_n18# XA3a/A XA2/MN0/a_324_n18# AVSS XA3/N1 SUNSAR_SARCMPHX1_CV
XXA3 CNI XA9/Y XA3a/A XA3/N2 AVDD AVSS XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVDD
+ XA3/MP0/a_216_n18# XA3/CO XA3/MN0/a_324_n18# AVSS XA3/N1 SUNSAR_SARCMPHX1_CV
XXA4 CNI AVDD AVDD AVSS XA9/MP0/a_216_n18# XA9/MN0/a_324_n18# XA9/A XA4/MP0/a_216_n18#
+ XA9/Y XA4/MN0/a_324_n18# AVSS SUNSAR_SARKICKHX1_CV
XXA3a AVDD AVSS XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVDD XA3a/MP0/a_216_n18# CNO
+ XA3a/A XA3a/MN0/a_324_n18# AVSS SUNSAR_IVX4_CV
XXA2a AVDD AVSS XA3a/MP0/a_216_n18# XA3a/MN0/a_324_n18# AVDD XA2/MP6/a_216_334# CPO
+ XA3/CO XA2/MN6/a_324_334# AVSS SUNSAR_IVX4_CV
XXA9 AVDD AVSS XA9/Y XA9/MP0/a_216_n18# XA9/MP0/a_216_334# AVDD XA9/A XA9/MN0/a_324_n18#
+ AVSS XA9/MN0/a_324_334# SUNSAR_IVX1_CV
C0 XA4/MP0/a_216_n18# AVDD -0.311987f
C1 XA9/Y XA3a/A 0.391167f
C2 XA3/MP0/a_216_n18# AVDD -0.313369f
C3 XA9/A AVDD 0.189383f
C4 XA3a/A CPO 0.108133f
C5 XA3/CO AVDD 1.166637f
C6 XA3/N1 AVDD 0.195531f
C7 XA2/MP6/a_216_334# AVDD -0.313518f
C8 XA12/Y CK_SAMPLE 0.106092f
C9 XA2/MP0/a_216_n18# AVDD -0.311986f
C10 XA3/CO XA9/A 0.141462f
C11 XA11/Y XA12/Y 0.130476f
C12 XA3a/MP0/a_216_n18# AVDD -0.312264f
C13 XA3/N1 CNO 0.113873f
C14 XA3/N1 XA3/CO 0.289212f
C15 CNI XA9/A 0.362147f
C16 XA12/MP0/a_216_n18# AVDD -0.312799f
C17 XA9/A CPI 0.297822f
C18 XA3a/A AVDD 0.912932f
C19 XA13/MP1/a_216_n18# AVDD -0.311986f
C20 XA3/N1 CPI 0.115376f
C21 XA3a/A XA9/A 0.136678f
C22 XA9/MP0/a_216_n18# AVDD -0.311986f
C23 XA3a/A XA3/CO 1.092423f
C24 XA12/Y AVDD 0.490048f
C25 XA9/Y AVDD 0.164728f
C26 XA3/N1 XA3a/A 0.309118f
C27 XA9/Y XA9/A 1.524979f
C28 XA9/Y XA3/CO 0.24121f
C29 XA9/MP0/a_216_334# AVDD -0.311309f
C30 XA11/Y XA9/A 0.268591f
C31 XA11/MP0/a_216_n18# AVDD -0.312939f
C32 XA3/N1 XA9/Y 0.106124f
C33 XA1/MP0/a_216_n18# AVDD -0.311986f
C34 XA9/Y CNI 0.382485f
C35 XA9/Y CPI 0.27081f
C36 XA9/MN0/a_324_n18# AVSS 0.355152f
C37 XA3/CO AVSS 2.700073f
C38 CPO AVSS 0.178234f
C39 XA2/MN6/a_324_334# AVSS 0.353692f
C40 XA3a/A AVSS 2.521704f
C41 XA3/MN0/a_324_n18# AVSS 0.353692f
C42 CNO AVSS 0.179699f
C43 XA3a/MN0/a_324_n18# AVSS 0.353692f
C44 XA4/MN0/a_324_n18# AVSS 0.3537f
C45 XA4/MP0/S AVSS 0.414246f
C46 CNI AVSS 3.621781f
C47 XA3/N2 AVSS 0.246915f
C48 XA9/Y AVSS 4.611301f
C49 XA2/N2 AVSS 0.246915f
C50 XA2/MN0/a_324_n18# AVSS 0.353761f
C51 XA3/N1 AVSS 1.207811f
C52 AVDD AVSS 46.225964f
C53 CPI AVSS 3.746344f
C54 XA1/MN0/a_324_n18# AVSS 0.356268f
C55 XA1/MP0/S AVSS 0.422681f
C56 XA9/A AVSS 4.708538f
C57 XA0/MN1/a_324_n18# AVSS 0.422415f
C58 XA13/MN1/a_324_n18# AVSS 0.356268f
C59 XA13/MN1/a_324_334# AVSS 0.422f
C60 CK_CMP AVSS 0.538462f
C61 XA12/MN0/a_324_n18# AVSS 0.356976f
C62 XA11/MN0/a_324_n18# AVSS 0.354241f
C63 DONE AVSS 0.474555f
C64 CK_SAMPLE AVSS 0.470196f
C65 XA9/MN0/a_324_334# AVSS 0.355744f
C66 XA12/Y AVSS 0.688417f
C67 XA11/Y AVSS 0.835238f
.ends

.subckt SUNSAR_NCHDLR D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 G B 0.415197f
C1 a_324_n18# B 0.422415f
C2 a_324_334# B 0.422f
.ends

.subckt SUNSAR_CAP_BSSW_CV A B VSUBS
R0 A m3_6948_120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R1 m3_252_280# B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
C0 A B 65.019196f
C1 m3_6948_120# B 0.172147f
C2 m3_252_280# A 0.105547f
C3 B VSUBS 13.2906f
C4 A VSUBS 13.2887f
.ends

.subckt SUNSAR_CAP_BSSW5_CV B A VSUBS
XXCAPB0 A B VSUBS SUNSAR_CAP_BSSW_CV
XXCAPB1 A B VSUBS SUNSAR_CAP_BSSW_CV
XXCAPB2 A B VSUBS SUNSAR_CAP_BSSW_CV
XXCAPB3 A B VSUBS SUNSAR_CAP_BSSW_CV
XXCAPB4 A B VSUBS SUNSAR_CAP_BSSW_CV
C0 A B 54.00426f
C1 B VSUBS 54.06679f
C2 A VSUBS 55.079098f
.ends

.subckt SUNSAR_TIEH_CV Y BULKP AVDD AVSS MP0/G MP0/a_216_n18# MP0/a_216_334# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 Y MP0/G AVDD BULKP MP0/a_216_n18# MP0/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 MP0/G MP0/G AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.106173f
C1 BULKP MP0/G 0.112786f
C2 AVDD VSUBS 0.24902f
C3 AVSS VSUBS 0.367715f
C4 MP0/G VSUBS 0.790179f
C5 MN0/a_324_n18# VSUBS 0.422415f
C6 MN0/a_324_334# VSUBS 0.422f
C7 BULKP VSUBS 2.806854f
.ends

.subckt SUNSAR_TIEL_CV BULKP AVDD AVSS MP0/G Y MP0/a_216_n18# MP0/a_216_334# MN0/a_324_n18#
+ VSUBS MN0/a_324_334#
XMP0 MP0/G MP0/G AVDD BULKP MP0/a_216_n18# MP0/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 Y MP0/G AVSS VSUBS MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.103703f
C1 BULKP MP0/G 0.161174f
C2 AVDD VSUBS 0.249049f
C3 AVSS VSUBS 0.370369f
C4 MP0/G VSUBS 0.708387f
C5 MN0/a_324_n18# VSUBS 0.422415f
C6 MN0/a_324_334# VSUBS 0.422f
C7 BULKP VSUBS 2.806659f
.ends

.subckt SUNSAR_TGPD_CV AVSS MP2/B MN2/a_324_334# MP0/S B MP0/a_216_n18# A C MP2/a_216_334#
+ MN0/a_324_n18# VSUBS AVDD
XMP1_DMY B AVDD AVDD MP2/B C C VSUBS SUNSAR_PCHDL
XMP0 AVDD C MP0/S MP2/B MP0/a_216_n18# AVDD VSUBS SUNSAR_PCHDL
XMN0 AVSS C MP0/S VSUBS MN0/a_324_n18# C SUNSAR_NCHDL
XMP2 A C B MP2/B AVDD MP2/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 B C AVSS VSUBS C MP0/S SUNSAR_NCHDL
XMN2 A MP0/S B VSUBS C MN2/a_324_334# SUNSAR_NCHDL
C0 C MP2/B -0.388363f
C1 C MP0/S 0.148714f
C2 MP2/B AVDD -0.506518f
C3 B A 0.108f
C4 AVDD VSUBS 0.478784f
C5 AVSS VSUBS 0.352742f
C6 A VSUBS 0.204323f
C7 MN2/a_324_334# VSUBS 0.422f
C8 MP2/B VSUBS 4.387254f
C9 MP0/S VSUBS 0.747699f
C10 MN0/a_324_n18# VSUBS 0.422415f
C11 C VSUBS 0.995573f
.ends

.subckt SUNSAR_SARBSSWCTRL_CV GN GNG TIE_H BULKP AVDD AVSS MN1/a_324_334# C MP0/a_216_n18#
+ MP1/a_216_334# MN0/a_324_n18# VSUBS
XMP0 GNG C GN BULKP MP0/a_216_n18# GN VSUBS SUNSAR_PCHDL
XMP1 AVDD GN GNG BULKP C MP1/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 MN1/S C AVSS VSUBS MN0/a_324_n18# TIE_H SUNSAR_NCHDL
XMN1 GN TIE_H MN1/S VSUBS C MN1/a_324_334# SUNSAR_NCHDL
C0 BULKP GN -0.16538f
C1 BULKP C -0.234337f
C2 C GN 0.105655f
C3 BULKP AVDD 0.119037f
C4 AVDD VSUBS 0.263047f
C5 AVSS VSUBS 0.384798f
C6 TIE_H VSUBS 0.37082f
C7 GN VSUBS 0.410388f
C8 MN1/a_324_334# VSUBS 0.422f
C9 C VSUBS 0.568156f
C10 MN0/a_324_n18# VSUBS 0.422415f
C11 BULKP VSUBS 3.595271f
.ends

.subckt SUNSAR_SARBSSW_CV VI CK CKN TIE_L VO1 M4/G VO2 XA3/B XA4/GNG AVDD AVSS
XM1 VI M4/G VO1 AVSS M1/a_324_n18# M2/a_324_n18# SUNSAR_NCHDLR
XM2 VI M4/G VO1 AVSS M2/a_324_n18# M3/a_324_n18# SUNSAR_NCHDLR
XM3 VI M4/G VO1 AVSS M3/a_324_n18# M4/a_324_n18# SUNSAR_NCHDLR
XM4 VI M4/G VO1 AVSS M4/a_324_n18# M5/a_324_n18# SUNSAR_NCHDLR
XM5 VI TIE_L VO2 AVSS M5/a_324_n18# M6/a_324_n18# SUNSAR_NCHDLR
XXCAPB1 XA3/B XA4/GNG AVSS SUNSAR_CAP_BSSW5_CV
XM6 VI TIE_L VO2 AVSS M6/a_324_n18# M7/a_324_n18# SUNSAR_NCHDLR
XM7 VI TIE_L VO2 AVSS M7/a_324_n18# M8/a_324_n18# SUNSAR_NCHDLR
XM8 VI TIE_L VO2 AVSS M8/a_324_n18# M8/a_324_334# SUNSAR_NCHDLR
XXA0 AVDD AVSS CKN XA0/MP0/a_216_n18# XA3/MP0/a_216_n18# AVDD CK XA0/MN0/a_324_n18#
+ AVSS XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA1 XA1/Y AVDD AVDD AVSS XA1/MP0/G XA4/MP1/a_216_334# XA7/MP1/a_216_n18# XA4/MN1/a_324_334#
+ AVSS XA7/MN1/a_324_n18# SUNSAR_TIEH_CV
XXA2 AVDD AVDD AVSS XA2/MP0/G TIE_L XA7/MP1/a_216_334# XA5/MP1/a_216_n18# XA7/MN1/a_324_334#
+ AVSS XA5/MN1/a_324_n18# SUNSAR_TIEL_CV
XXA3 AVSS AVDD XA4/MN0/a_324_n18# XA3/MP0/S XA3/B XA3/MP0/a_216_n18# VI CKN XA4/MP0/a_216_n18#
+ XA3/MN0/a_324_n18# AVSS AVDD SUNSAR_TGPD_CV
XXA5 AVDD XA5/MN1/a_324_n18# XA5/MN1/a_324_334# XA5/MP1/a_216_334# XA5/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA4 M4/G XA4/GNG XA1/Y AVDD AVDD AVSS XA4/MN1/a_324_334# CKN XA4/MP0/a_216_n18# XA4/MP1/a_216_334#
+ XA4/MN0/a_324_n18# AVSS SUNSAR_SARBSSWCTRL_CV
XXA5b AVDD XA5b/MN1/a_324_n18# XA0/MN0/a_324_n18# XA0/MP0/a_216_n18# XA5b/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA7 AVDD XA7/MN1/a_324_n18# XA7/MN1/a_324_334# XA7/MP1/a_216_334# XA7/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
C0 AVSS XA1/Y 0.269286f
C1 XA3/B AVDD 1.133969f
C2 XA5/MP1/a_216_n18# AVDD -0.311986f
C3 VO2 AVSS 0.115254f
C4 XA4/GNG AVDD 2.405915f
C5 TIE_L AVSS 0.570893f
C6 AVSS CKN 0.456081f
C7 M4/G VO1 0.121857f
C8 VI VO1 0.509495f
C9 VI M4/G 0.733023f
C10 AVDD XA1/Y 0.335195f
C11 AVDD XA7/MP1/a_216_n18# -0.314016f
C12 XA1/MP0/G XA1/Y 0.210055f
C13 AVDD CKN 0.381615f
C14 XA4/MP1/a_216_334# AVDD -0.310882f
C15 XA7/MP1/a_216_334# AVDD -0.311812f
C16 XA3/B CKN 0.220083f
C17 XA4/GNG CKN 0.13356f
C18 XA0/MP0/a_216_n18# AVDD -0.310529f
C19 VO1 AVSS 0.112136f
C20 M4/G AVSS 0.641192f
C21 VI AVSS 0.44414f
C22 AVDD XA4/MP0/a_216_n18# -0.315004f
C23 M4/G XA4/GNG 0.159364f
C24 M4/G XA1/Y 0.191529f
C25 VI VO2 0.402032f
C26 VI TIE_L 0.431895f
C27 M4/G CKN 0.164954f
C28 VI CKN 0.158203f
C29 AVDD AVSS 0.15268f
C30 AVDD XA3/MP0/a_216_n18# -0.315912f
C31 AVDD XA2/MP0/G 0.154505f
C32 XA3/MP0/S CKN 0.35416f
C33 XA7/MN1/a_324_n18# 0 0.359583f
C34 AVSS 0 2.93973f
C35 XA5b/MN1/a_324_n18# 0 0.422415f
C36 AVDD 0 16.012844f
C37 XA1/Y 0 0.690197f
C38 CKN 0 1.768971f
C39 XA4/MN0/a_324_n18# 0 0.359583f
C40 XA5/MN1/a_324_334# 0 0.422f
C41 XA3/MP0/S 0 0.743486f
C42 XA3/MN0/a_324_n18# 0 0.359583f
C43 XA2/MP0/G 0 0.708335f
C44 XA7/MN1/a_324_334# 0 0.359583f
C45 XA5/MN1/a_324_n18# 0 0.360407f
C46 XA1/MP0/G 0 0.788614f
C47 XA4/MN1/a_324_334# 0 0.359583f
C48 CK 0 0.513823f
C49 XA0/MN0/a_324_n18# 0 0.359583f
C50 M8/a_324_n18# 0 0.356977f
C51 M8/a_324_334# 0 0.422f
C52 M6/a_324_n18# 0 0.356977f
C53 M7/a_324_n18# 0 0.356977f
C54 XA3/B 0 54.41209f
C55 XA4/GNG 0 53.065117f
C56 VO2 0 0.317444f
C57 TIE_L 0 2.408263f
C58 M5/a_324_n18# 0 0.356977f
C59 M3/a_324_n18# 0 0.356977f
C60 M4/a_324_n18# 0 0.356977f
C61 VO1 0 0.370636f
C62 M4/G 0 2.475647f
C63 VI 0 1.254522f
C64 M1/a_324_n18# 0 0.422415f
C65 M2/a_324_n18# 0 0.356977f
.ends

.subckt SUNSAR_SAREMX1_CV B EN ENO AVDD MP3/a_216_334# MN3/a_324_334# A BULKP MP0/a_216_n18#
+ AVSS RST_N MN0/a_324_n18# VSUBS
XMP0 AVDD RST_N MP3/G BULKP MP0/a_216_n18# MP1/a_216_n18# VSUBS SUNSAR_PCHDL
XMP1 MP2/S B ENO BULKP MP1/a_216_n18# MP2/a_216_n18# VSUBS SUNSAR_PCHDL
XMP2 MP3/S A MP2/S BULKP MP2/a_216_n18# MP3/a_216_n18# VSUBS SUNSAR_PCHDL
XMN0 MN2/S EN MP3/G VSUBS MN0/a_324_n18# MN1/a_324_n18# SUNSAR_NCHDL
XMP3 AVDD MP3/G MP3/S BULKP MP3/a_216_n18# MP3/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 MN2/S B AVSS VSUBS MN1/a_324_n18# MN2/a_324_n18# SUNSAR_NCHDL
XMN2 AVSS A MN2/S VSUBS MN2/a_324_n18# MN3/a_324_n18# SUNSAR_NCHDL
XMN3 ENO MP3/G AVSS VSUBS MN3/a_324_n18# MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP A 0.108551f
C1 BULKP B 0.113772f
C2 ENO MP3/G 0.133485f
C3 MP3/G AVDD 0.124994f
C4 BULKP MP3/a_216_n18# -0.311038f
C5 MN2/S AVSS 0.206972f
C6 BULKP MP3/G 0.480172f
C7 BULKP MP2/a_216_n18# -0.311038f
C8 ENO AVDD 0.155663f
C9 BULKP ENO 0.182005f
C10 BULKP MP1/a_216_n18# -0.311038f
C11 AVSS AVDD 0.157524f
C12 MP3/G A 0.105132f
C13 BULKP AVDD 0.233317f
C14 AVDD VSUBS 0.390025f
C15 AVSS VSUBS 0.695296f
C16 MN3/a_324_n18# VSUBS 0.35253f
C17 MN3/a_324_334# VSUBS 0.422f
C18 A VSUBS 0.498033f
C19 MN2/a_324_n18# VSUBS 0.352522f
C20 B VSUBS 0.513991f
C21 MN1/a_324_n18# VSUBS 0.352522f
C22 MP3/G VSUBS 0.827536f
C23 EN VSUBS 0.386445f
C24 MN2/S VSUBS 0.207484f
C25 MN0/a_324_n18# VSUBS 0.422415f
C26 ENO VSUBS 0.246284f
C27 BULKP VSUBS 7.539519f
.ends

.subckt SUNSAR_SARLTX1_CV RST_N EN LCK_N AVDD AVSS MN2/a_324_334# A BULKP MP0/a_216_n18#
+ CHL MP2/a_216_334# MN0/a_324_n18# VSUBS
XMP0 MP1/S RST_N AVDD BULKP MP0/a_216_n18# RST_N VSUBS SUNSAR_PCHDL
XMP1 MP2/S RST_N MP1/S BULKP RST_N RST_N VSUBS SUNSAR_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# LCK_N SUNSAR_NCHDL
XMP2 CHL RST_N MP2/S BULKP RST_N MP2/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 MN2/S LCK_N MN1/S VSUBS A EN SUNSAR_NCHDL
XMN2 CHL EN MN2/S VSUBS LCK_N MN2/a_324_334# SUNSAR_NCHDL
C0 BULKP RST_N -1.319845f
C1 AVDD BULKP 0.143379f
C2 EN VSUBS 0.372036f
C3 MN2/a_324_334# VSUBS 0.422f
C4 LCK_N VSUBS 0.335836f
C5 AVSS VSUBS 0.428199f
C6 RST_N VSUBS 0.123012f
C7 CHL VSUBS 0.260933f
C8 BULKP VSUBS 4.387078f
C9 A VSUBS 0.372036f
C10 MN0/a_324_n18# VSUBS 0.422415f
C11 AVDD VSUBS 0.276832f
.ends

.subckt SUNSAR_SARMRYX1_CV CMP_OP CHL_OP CHL_ON RST_N XA5/MP2/a_216_334# ENO XA5/MN2/a_324_334#
+ CMP_ON AVDD AVSS XA2/Y EN
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA1 CMP_ON EN ENO AVDD XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# CMP_OP AVDD XA1/MP0/a_216_n18#
+ AVSS RST_N XA1/MN0/a_324_n18# AVSS SUNSAR_SAREMX1_CV
XXA2 AVDD AVSS XA2/Y XA2/MP0/a_216_n18# XA4/MP0/a_216_n18# AVDD ENO XA2/MN0/a_324_n18#
+ AVSS XA4/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA4 RST_N EN XA2/Y AVDD AVSS XA5/MN0/a_324_n18# CMP_OP AVDD XA4/MP0/a_216_n18# CHL_OP
+ XA5/MP0/a_216_n18# XA4/MN0/a_324_n18# AVSS SUNSAR_SARLTX1_CV
XXA5 RST_N EN XA2/Y AVDD AVSS XA5/MN2/a_324_334# CMP_ON AVDD XA5/MP0/a_216_n18# CHL_ON
+ XA5/MP2/a_216_334# XA5/MN0/a_324_n18# AVSS SUNSAR_SARLTX1_CV
C0 AVDD XA4/MP0/a_216_n18# -0.31403f
C1 EN XA2/Y 0.114038f
C2 EN CMP_OP 0.196887f
C3 AVDD XA5/MP0/a_216_n18# -0.31403f
C4 ENO CMP_OP 0.15365f
C5 XA2/MP0/a_216_n18# AVDD -0.31403f
C6 XA1/MP0/a_216_n18# AVDD -0.311986f
C7 XA2/Y CMP_ON 0.130187f
C8 AVDD RST_N 1.195814f
C9 CMP_OP XA2/Y 0.183507f
C10 EN CMP_ON 0.54292f
C11 XA5/MN2/a_324_334# AVSS 0.422f
C12 CHL_ON AVSS 0.232377f
C13 CMP_ON AVSS 1.822119f
C14 XA5/MN0/a_324_n18# AVSS 0.3537f
C15 RST_N AVSS 0.223373f
C16 CHL_OP AVSS 0.170032f
C17 XA4/MN0/a_324_n18# AVSS 0.3537f
C18 XA2/Y AVSS 1.191276f
C19 XA2/MN0/a_324_n18# AVSS 0.353715f
C20 XA1/MN3/a_324_n18# AVSS 0.352733f
C21 CMP_OP AVSS 1.302224f
C22 XA1/MN2/a_324_n18# AVSS 0.353381f
C23 XA1/MN1/a_324_n18# AVSS 0.358f
C24 XA1/MP3/G AVSS 0.885586f
C25 EN AVSS 2.425524f
C26 XA1/MN2/S AVSS 0.199983f
C27 XA1/MN0/a_324_n18# AVSS 0.356268f
C28 ENO AVSS 0.8336f
C29 XA0/MN1/a_324_n18# AVSS 0.422415f
C30 AVDD AVSS 17.159056f
.ends

.subckt SUNSAR_SWX4_CV MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18# Y AVSS A
+ MN0/a_324_n18# VREF VSUBS
XMP0 Y A VREF BULKP MP0/a_216_n18# A VSUBS SUNSAR_PCHDL
XMP1 VREF A Y BULKP A A VSUBS SUNSAR_PCHDL
XMP2 Y A VREF BULKP A A VSUBS SUNSAR_PCHDL
XMN0 Y A AVSS VSUBS MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 VREF A Y BULKP A MP3/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 AVSS A Y VSUBS A A SUNSAR_NCHDL
XMN2 Y A AVSS VSUBS A A SUNSAR_NCHDL
XMN3 AVSS A Y VSUBS A MN3/a_324_334# SUNSAR_NCHDL
C0 A VREF 0.184236f
C1 Y VREF 0.133073f
C2 Y A 0.147007f
C3 BULKP VREF 0.281929f
C4 BULKP A -1.606473f
C5 Y AVSS 0.180645f
C6 AVSS VSUBS 0.66508f
C7 MN3/a_324_334# VSUBS 0.422f
C8 VREF VSUBS 0.501044f
C9 A VSUBS 2.06236f
C10 Y VSUBS 0.278638f
C11 MN0/a_324_n18# VSUBS 0.422415f
C12 BULKP VSUBS 5.176431f
.ends

.subckt SUNSAR_SARCEX1_CV B Y RST AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18#
+ A MN0/a_324_n18# VSUBS
XMP0 MP1/S A Y BULKP MP0/a_216_n18# A VSUBS SUNSAR_PCHDL
XMP1 AVDD A MP1/S BULKP A B VSUBS SUNSAR_PCHDL
XMP2 MP3/S B AVDD BULKP A B VSUBS SUNSAR_PCHDL
XMN0 MN1/S RST AVSS VSUBS MN0/a_324_n18# RST SUNSAR_NCHDL
XMP3 Y B MP3/S BULKP B MP3/a_216_334# VSUBS SUNSAR_PCHDL
XMN1 AVSS RST MN1/S VSUBS RST RST SUNSAR_NCHDL
XMN2 MN3/S RST AVSS VSUBS RST RST SUNSAR_NCHDL
XMN3 Y RST MN3/S VSUBS RST MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP A -1.005062f
C1 AVDD BULKP 0.114602f
C2 BULKP Y 0.191403f
C3 AVDD AVSS 0.106506f
C4 AVSS Y 0.129646f
C5 BULKP B -1.00547f
C6 AVDD VSUBS 0.247044f
C7 Y VSUBS 0.484249f
C8 MN3/a_324_334# VSUBS 0.422f
C9 AVSS VSUBS 0.495556f
C10 RST VSUBS 1.501372f
C11 MN0/a_324_n18# VSUBS 0.422415f
C12 BULKP VSUBS 5.174408f
.ends

.subckt SUNSAR_SARDIGEX4_CV CMP_OP CMP_ON CP0 CP1 CN1 XA9/B DONE CN0 RST_N XA11/A
+ CEO XA4/A CKS ENO EN VREF CEIN XA12/A AVSS AVDD
XXA10 AVDD AVSS XA11/A XA9/MP1/a_216_334# XA11/MP0/a_216_n18# AVDD XA9/Y XA9/MN1/a_324_334#
+ AVSS XA11/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA11 AVDD AVSS XA12/MN0/a_324_n18# CEIN AVDD XA11/MP0/a_216_n18# XA12/A XA12/MP0/a_216_n18#
+ XA11/A XA11/MN0/a_324_n18# AVSS SUNSAR_NRX1_CV
XXA12 AVDD AVSS CEO XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD XA12/A XA12/MN0/a_324_n18#
+ AVSS XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVDD XA13/MN1/a_324_n18# XA13/MN1/a_324_334# XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA1 CMP_OP XA4/A XA2/A RST_N XA2/MP0/a_216_n18# ENO XA2/MN0/a_324_n18# CMP_ON AVDD
+ AVSS XA1/XA2/Y EN SUNSAR_SARMRYX1_CV
XXA2 XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVDD XA2/MP0/a_216_n18# CN1 AVSS XA2/A
+ XA2/MN0/a_324_n18# VREF AVSS SUNSAR_SWX4_CV
XXA3 XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVDD XA3/MP0/a_216_n18# CP1 AVSS CN1 XA3/MN0/a_324_n18#
+ VREF AVSS SUNSAR_SWX4_CV
XXA5 XA6/MP0/a_216_n18# XA6/MN0/a_324_n18# AVDD XA5/MP0/a_216_n18# CN0 AVSS CP0 XA5/MN0/a_324_n18#
+ VREF AVSS SUNSAR_SWX4_CV
XXA4 XA5/MP0/a_216_n18# XA5/MN0/a_324_n18# AVDD XA4/MP0/a_216_n18# CP0 AVSS XA4/A
+ XA4/MN0/a_324_n18# VREF AVSS SUNSAR_SWX4_CV
XXA6 CP1 XA9/B CKS AVDD AVSS XA7/MP0/a_216_n18# XA7/MN0/a_324_n18# AVDD XA6/MP0/a_216_n18#
+ CN0 XA6/MN0/a_324_n18# AVSS SUNSAR_SARCEX1_CV
XXA7 AVDD AVSS XA9/A XA7/MP0/a_216_n18# XA8/MP0/a_216_n18# AVDD ENO XA7/MN0/a_324_n18#
+ AVSS XA8/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA8 AVDD AVSS DONE XA8/MP0/a_216_n18# XA9/MP0/a_216_n18# AVDD XA9/A XA8/MN0/a_324_n18#
+ AVSS XA9/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA9 XA9/Y AVDD AVSS XA9/MN1/a_324_334# XA9/B XA9/A AVDD XA9/MP0/a_216_n18# XA9/MP1/a_216_334#
+ XA9/MN0/a_324_n18# AVSS SUNSAR_NDX1_CV
C0 AVDD XA8/MP0/a_216_n18# -0.311987f
C1 CEIN XA12/A 0.110841f
C2 AVDD CN1 0.114213f
C3 AVDD CP1 0.743971f
C4 XA11/MP0/a_216_n18# AVDD -0.311842f
C5 CP0 XA4/A 0.350838f
C6 XA13/MP1/a_216_n18# AVDD -0.311986f
C7 EN XA4/A 0.118846f
C8 AVDD ENO 2.495094f
C9 CN1 XA4/A 0.466806f
C10 CP1 XA4/A 0.193274f
C11 XA2/A VREF 0.115624f
C12 AVDD XA5/MP0/a_216_n18# -0.298676f
C13 ENO XA4/A 0.119578f
C14 XA2/A CN1 0.327387f
C15 ENO RST_N 0.661116f
C16 AVDD XA9/MP1/a_216_334# -0.311908f
C17 AVDD XA3/MP0/a_216_n18# -0.298153f
C18 AVDD XA2/MP0/a_216_n18# -0.306139f
C19 XA9/Y XA11/A 0.134948f
C20 AVDD XA4/A 0.106262f
C21 CN0 CP0 0.298273f
C22 XA9/A XA9/B 0.245863f
C23 CP1 CP0 0.176643f
C24 AVDD XA2/A 0.202922f
C25 CP1 CN0 0.319562f
C26 AVDD XA9/MP0/a_216_n18# -0.311986f
C27 CP1 VREF 1.096312f
C28 CP1 CN1 0.208539f
C29 XA1/XA2/Y XA4/A 0.161989f
C30 ENO VREF 0.694105f
C31 XA2/A XA4/A 0.111482f
C32 XA9/Y XA9/B 0.108031f
C33 ENO CP1 0.402013f
C34 AVDD XA7/MP0/a_216_n18# -0.311987f
C35 XA12/MP0/a_216_n18# AVDD -0.311309f
C36 AVDD XA6/MP0/a_216_n18# -0.306081f
C37 AVDD XA4/MP0/a_216_n18# -0.298676f
C38 AVDD CP0 0.163708f
C39 AVDD CN0 0.409213f
C40 AVDD VREF 2.204398f
C41 XA9/MN1/a_324_334# AVSS 0.355152f
C42 XA9/MN0/a_324_n18# AVSS 0.3539f
C43 XA9/A AVSS 1.385171f
C44 DONE AVSS 0.144639f
C45 XA7/MN0/a_324_n18# AVSS 0.354718f
C46 XA8/MN0/a_324_n18# AVSS 0.355152f
C47 XA9/B AVSS 1.502326f
C48 CKS AVSS 1.45158f
C49 XA6/MN0/a_324_n18# AVSS 0.356268f
C50 XA4/A AVSS 3.131355f
C51 XA4/MN0/a_324_n18# AVSS 0.355744f
C52 CP0 AVSS 2.560386f
C53 CN0 AVSS 0.340136f
C54 XA5/MN0/a_324_n18# AVSS 0.355152f
C55 VREF AVSS 0.8336f
C56 CN1 AVSS 2.510553f
C57 CP1 AVSS 0.513004f
C58 XA3/MN0/a_324_n18# AVSS 0.355152f
C59 XA2/A AVSS 2.066712f
C60 XA2/MN0/a_324_n18# AVSS 0.355744f
C61 CMP_ON AVSS 1.344542f
C62 XA1/XA5/MN0/a_324_n18# AVSS 0.359841f
C63 RST_N AVSS 0.189551f
C64 XA1/XA4/MN0/a_324_n18# AVSS 0.360407f
C65 XA1/XA2/Y AVSS 1.04564f
C66 XA1/XA2/MN0/a_324_n18# AVSS 0.360407f
C67 XA1/XA1/MN3/a_324_n18# AVSS 0.355196f
C68 CMP_OP AVSS 1.158538f
C69 XA1/XA1/MN2/a_324_n18# AVSS 0.355196f
C70 XA1/XA1/MN1/a_324_n18# AVSS 0.355196f
C71 XA1/XA1/MP3/G AVSS 0.827195f
C72 EN AVSS 2.11207f
C73 XA1/XA1/MN2/S AVSS 0.200627f
C74 XA1/XA1/MN0/a_324_n18# AVSS 0.360407f
C75 ENO AVSS 1.875766f
C76 XA1/XA0/MN1/a_324_n18# AVSS 0.422415f
C77 AVDD AVSS 49.97179f
C78 XA13/MN1/a_324_334# AVSS 0.422f
C79 CEO AVSS 0.198916f
C80 XA12/MN0/a_324_n18# AVSS 0.355467f
C81 XA13/MN1/a_324_n18# AVSS 0.356268f
C82 XA12/A AVSS 0.87316f
C83 XA11/MN0/a_324_n18# AVSS 0.355152f
C84 CEIN AVSS 0.470391f
C85 XA11/A AVSS 0.773693f
C86 XA9/Y AVSS 0.833f
.ends

.subckt SUNSAR_SAR8B_CV SAR_IP SAR_IN DONE D<7> D<4> D<1> EN CK_SAMPLE_BSSW XA6/CN0
+ XA6/CP0 XA3/CN0 XA3/CP0 CK_SAMPLE D<0> XA7/CP0 XA0/CEIN XA4/CN0 D<3> XA4/CP0 XA1/CN0
+ D<6> XA1/CP0 SARP XA5/CN0 D<2> XA5/CP0 XA2/CN0 D<5> VREF XA2/CP0 SARN AVDD AVSS
XXDAC1 XA0/CP1 XA0/CP0 D<6> XA1/CP0 D<5> XA2/CP0 D<4> D<3> D<2> D<1> SARP AVSS AVSS
+ SUNSAR_CDAC7_CV
XXDAC2 D<7> XA0/CN0 XA1/CN1 XA1/CN0 XA2/CN1 XA2/CN0 XA3/CN0 XA4/CN0 XA5/CN0 XA6/CN0
+ SARN AVSS AVSS SUNSAR_CDAC7_CV
XXA20 SARP SARN XA7/CEO CK_SAMPLE DONE XA20/XA9/A XA20/CPO AVDD XA20/CNO AVSS SUNSAR_SARCMPX1_CV
XXB1 SAR_IP CK_SAMPLE_BSSW XB1/CKN XA0/CEIN SARP XB1/M4/G SARN XB1/XA3/B XB1/XA4/GNG
+ AVDD AVSS SUNSAR_SARBSSW_CV
XXA0 XA20/CPO XA20/CNO XA0/CP0 XA0/CP1 D<7> XA0/XA9/B XA0/DONE XA0/CN0 EN XA0/XA11/A
+ XA0/CEO XA0/XA4/A CK_SAMPLE XA1/EN EN VREF XA0/CEIN XA0/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXB2 SAR_IN CK_SAMPLE_BSSW XB2/CKN XA0/CEIN SARN XB2/M4/G SARP XB2/XA3/B XB2/XA4/GNG
+ AVDD AVSS SUNSAR_SARBSSW_CV
XXA1 XA20/CPO XA20/CNO XA1/CP0 D<6> XA1/CN1 XA1/XA9/B XA1/DONE XA1/CN0 EN XA1/XA11/A
+ XA1/CEO XA1/XA4/A CK_SAMPLE XA2/EN XA1/EN VREF XA0/CEO XA1/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA2 XA20/CPO XA20/CNO XA2/CP0 D<5> XA2/CN1 XA2/XA9/B XA2/DONE XA2/CN0 EN XA2/XA11/A
+ XA2/CEO XA2/XA4/A CK_SAMPLE XA3/EN XA2/EN VREF XA1/CEO XA2/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA3 XA20/CPO XA20/CNO XA3/CP0 D<4> XA3/CN1 XA3/XA9/B XA3/DONE XA3/CN0 EN XA3/XA11/A
+ XA3/CEO XA3/XA4/A CK_SAMPLE XA4/EN XA3/EN VREF XA2/CEO XA3/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA4 XA20/CPO XA20/CNO XA4/CP0 D<3> XA4/CN1 XA4/XA9/B XA4/DONE XA4/CN0 EN XA4/XA11/A
+ XA4/CEO XA4/XA4/A CK_SAMPLE XA5/EN XA4/EN VREF XA3/CEO XA4/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA5 XA20/CPO XA20/CNO XA5/CP0 D<2> XA5/CN1 XA5/XA9/B XA5/DONE XA5/CN0 EN XA5/XA11/A
+ XA5/CEO XA5/XA4/A CK_SAMPLE XA6/EN XA5/EN VREF XA4/CEO XA5/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA6 XA20/CPO XA20/CNO XA6/CP0 D<1> XA6/CN1 XA6/XA9/B XA6/DONE XA6/CN0 EN XA6/XA11/A
+ XA6/CEO XA6/XA4/A CK_SAMPLE XA7/EN XA6/EN VREF XA5/CEO XA6/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA7 XA20/CPO XA20/CNO XA7/CP0 D<0> XA7/CN1 XA7/XA9/B DONE XA7/CN0 EN XA7/XA11/A XA7/CEO
+ XA7/XA4/A CK_SAMPLE XA7/ENO XA7/EN VREF XA6/CEO XA7/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
C0 XA0/CP1 CK_SAMPLE 0.100695f
C1 XA5/CEO XA5/XA11/A 0.13078f
C2 XA7/ENO XA7/EN 0.779051f
C3 AVSS XA2/CEO 0.266939f
C4 XA20/CNO XA3/XA4/A 0.286128f
C5 XA5/CEO AVSS 0.43736f
C6 EN XA20/CNO 2.032689f
C7 XA1/EN XA20/CPO 0.251162f
C8 XA6/CN0 XA5/CN0 1.883929f
C9 AVSS D<3> 1.876198f
C10 XA2/CN0 XA2/CN1 0.583006f
C11 XA2/CP0 D<4> 0.835772f
C12 XA6/CN0 AVDD 2.589874f
C13 AVSS XA4/CN0 0.234489f
C14 XA20/CPO XA6/EN 0.378571f
C15 SARN XA0/CEIN 0.265285f
C16 D<1> D<3> 0.181155f
C17 XA2/CN1 D<2> 0.137975f
C18 VREF XA0/CEO 0.348781f
C19 XA2/CN0 XA1/CN0 2.065852f
C20 CK_SAMPLE D<2> 0.1008f
C21 XA1/CP0 XA2/CN1 0.143675f
C22 XA20/XA9/A XA20/CNO 0.101825f
C23 XA20/XA9/A XA7/XA4/A 0.11382f
C24 XA20/CPO XA2/EN 0.378571f
C25 EN VREF 0.66498f
C26 AVSS XA20/CPO 1.947881f
C27 XA1/CN0 XA2/CN1 0.547507f
C28 AVSS XA3/EN 0.214912f
C29 XA3/CEO AVSS 0.437359f
C30 VREF XA2/CEO 0.348781f
C31 XA1/CN0 XA1/CP0 3.345594f
C32 XDAC1/XC1/XRES16/B XB1/XA4/GNG 0.107427f
C33 CK_SAMPLE D<0> 0.102094f
C34 XA0/CEIN AVDD 9.065545f
C35 AVDD XA0/CEO 1.256112f
C36 XA20/CPO XA20/CNO 6.984268f
C37 XDAC1/XC1/XRES1A/B XB1/XA4/GNG 0.386137f
C38 XA1/CEO AVDD 0.342105f
C39 XA20/XA3/CO XA20/CPO 0.104539f
C40 XA20/CNO XA3/EN 0.302924f
C41 XA1/CEO XA1/XA12/A 0.264746f
C42 XA20/XA9/A SARN 0.113134f
C43 XA7/CEO AVDD 0.348014f
C44 AVDD EN 2.755226f
C45 AVSS XA2/CP0 0.193422f
C46 XA6/CN0 XA6/CP0 0.125928f
C47 XA5/EN XA6/EN 1.263077f
C48 XA0/CP1 XA1/CN1 0.268769f
C49 AVDD XA2/CEO 1.256112f
C50 XA5/CEO AVDD 0.342105f
C51 XA0/CP1 D<6> 1.561198f
C52 AVSS XA3/DONE 0.267946f
C53 D<5> XA0/CP0 0.306186f
C54 XA4/CN0 XA5/CN0 1.362054f
C55 XA4/CN0 XA4/CP0 0.125928f
C56 VREF XA3/EN 0.175304f
C57 AVDD XA4/CN0 2.483943f
C58 AVSS XA5/EN 0.218031f
C59 D<4> XA3/CN0 1.581234f
C60 XA6/CEO AVSS 0.276115f
C61 XA1/CN1 XA2/CN1 2.837019f
C62 XA20/CNO XA5/EN 0.302925f
C63 XA0/CN0 XA1/CP0 0.398101f
C64 AVDD XA20/CPO 2.513656f
C65 XA1/CN1 XA1/CP0 0.174582f
C66 D<6> XA2/CN1 0.199516f
C67 XB1/M4/G SARP 0.144008f
C68 AVDD XA3/EN 0.79199f
C69 XA6/CN0 XA4/CN0 0.14269f
C70 XA20/CNO XA2/XA4/A 0.212166f
C71 XA3/CEO AVDD 0.342105f
C72 CK_SAMPLE D<6> 0.1008f
C73 AVSS XA7/EN 0.231176f
C74 XA0/CN0 XA1/CN0 2.961017f
C75 XA1/CN1 XA1/CN0 0.608838f
C76 D<6> XA1/CP0 4.060233f
C77 SAR_IP SARP 0.279047f
C78 XA1/CEO XA0/CEO 0.431792f
C79 XA0/CP1 D<7> 0.831597f
C80 XA20/CNO XA7/EN 0.39054f
C81 XDAC2/XC1/XRES1A/B XB2/XA4/GNG 0.386137f
C82 VREF XA5/EN 0.175304f
C83 AVSS XA4/EN 0.355405f
C84 XA6/CEO VREF 0.348791f
C85 AVSS XA3/CN0 0.25506f
C86 DONE AVSS 0.493308f
C87 XB1/M4/G SARN 0.156031f
C88 XA20/CNO XA4/EN 0.457818f
C89 XA5/CEO XA5/XA12/A 0.264747f
C90 SAR_IP SARN 0.203945f
C91 AVDD XA5/EN 0.791989f
C92 VREF XA7/EN 0.175304f
C93 CK_SAMPLE D<4> 0.1008f
C94 XA6/CEO AVDD 1.255434f
C95 XA1/CP0 D<4> 0.174549f
C96 AVSS XA5/DONE 0.267946f
C97 D<5> XA2/CP0 3.965242f
C98 EN XA2/XA2/A 0.11426f
C99 XA0/CP1 AVSS 1.87901f
C100 XA0/CN0 XA1/CN1 0.495948f
C101 D<3> XA4/CN0 1.470811f
C102 XB1/XA3/B AVSS 1.491396f
C103 VREF XA4/EN 0.175304f
C104 XA20/CPO EN 0.728023f
C105 XA6/CN0 XA5/EN 0.115359f
C106 AVDD XA7/EN 0.809492f
C107 SARP XB1/XA4/GNG 1.624342f
C108 EN XA3/EN 0.311923f
C109 D<6> XA1/CN1 0.616721f
C110 XB1/XA4/GNG AVSS 1.208553f
C111 XDAC2/XC1/XRES16/B XB2/XA4/GNG 0.107427f
C112 XA3/CEO XA2/CEO 0.431793f
C113 AVSS XA2/CN0 0.127755f
C114 XA2/EN XA2/CN1 0.336738f
C115 XA20/CNO XA1/XA4/A 0.286129f
C116 AVDD XA4/EN 0.11184f
C117 AVSS D<2> 1.856228f
C118 XA6/CEO XA7/XA12/A 0.115411f
C119 AVSS XA2/CN1 1.031315f
C120 XA20/XA9/A XA20/CPO 0.365673f
C121 AVDD XA3/CN0 2.477465f
C122 AVSS CK_SAMPLE 2.799086f
C123 AVSS XA1/CP0 0.19218f
C124 D<1> D<2> 1.784246f
C125 XA2/EN XA1/CN0 0.127391f
C126 XA20/CNO XA2/CN1 0.188581f
C127 D<1> CK_SAMPLE 0.100705f
C128 AVSS XA1/CN0 0.126506f
C129 XA0/CN0 D<7> 0.494507f
C130 D<7> XA1/CN1 2.492607f
C131 XA4/CEO AVSS 0.266939f
C132 XA20/CPO XA3/EN 0.251162f
C133 EN XA5/EN 0.311923f
C134 XA6/CEO XA7/CEO 0.137785f
C135 XA0/CEIN XB2/CKN 0.100038f
C136 XB1/M4/G XA0/CEIN 0.110451f
C137 XB1/XA3/B AVDD 0.185337f
C138 XA3/CEO XA3/XA12/A 0.264747f
C139 XA1/EN XA1/CN1 0.231611f
C140 XA20/CNO XA0/XA4/A 0.212166f
C141 VREF CK_SAMPLE 1.866437f
C142 EN XA7/EN 0.173811f
C143 XA20/XA3a/A XA20/CNO 0.119511f
C144 AVDD XA2/CN0 2.508129f
C145 EN XA3/XA2/A 0.11418f
C146 XA6/XA4/A XA20/CNO 0.212166f
C147 D<2> XA5/CN0 1.58415f
C148 XA20/XA3/N1 SARN 0.135724f
C149 XA4/CEO VREF 0.348781f
C150 AVSS XA4/DONE 0.2733f
C151 XA20/CPO XA5/EN 0.251162f
C152 EN XA4/EN 0.235383f
C153 XA2/EN XA1/CN1 0.107883f
C154 AVDD CK_SAMPLE 4.279234f
C155 XA0/CN0 AVSS 0.144488f
C156 AVSS XA1/CN1 1.316495f
C157 XA20/XA9/A XA7/EN 0.291697f
C158 XA7/CEO DONE 0.119439f
C159 XA0/CEIN XB1/CKN 0.100039f
C160 EN XA5/XA2/A 0.11418f
C161 AVDD XA1/CN0 2.473342f
C162 AVSS D<6> 1.853472f
C163 D<1> XA0/CN0 0.232115f
C164 XA0/CP1 XA0/CP0 4.153562f
C165 XA20/CNO XA1/CN1 0.19102f
C166 XA4/CEO AVDD 1.256112f
C167 XA6/CN0 D<2> 0.155398f
C168 XA20/CPO XA7/EN 0.251284f
C169 XA3/CN0 XA4/CN0 1.410099f
C170 XA0/CN0 SARN 0.109275f
C171 XA7/ENO VREF 0.175304f
C172 D<5> XA2/CN1 0.490947f
C173 D<5> CK_SAMPLE 0.100705f
C174 XA20/CPO XA4/EN 0.378571f
C175 D<5> XA1/CP0 0.762697f
C176 XA0/CP0 XA2/CN1 0.144778f
C177 XA3/EN XA4/EN 1.263078f
C178 SARP D<7> 0.187721f
C179 AVSS D<7> 1.140293f
C180 XA0/CP0 XA1/CP0 1.795396f
C181 EN XA4/XA2/A 0.11426f
C182 AVSS D<4> 1.856228f
C183 AVSS XA1/DONE 0.267946f
C184 XA20/CNO XA5/XA4/A 0.286129f
C185 XA20/CNO D<7> 0.17726f
C186 XA0/CN0 AVDD 2.477148f
C187 XA1/EN XA2/EN 1.263077f
C188 AVSS XA1/EN 0.167653f
C189 D<3> D<2> 0.983626f
C190 AVSS XA6/EN 0.355405f
C191 XA2/CN1 D<3> 0.105016f
C192 XA1/EN XA20/CNO 0.302765f
C193 CK_SAMPLE D<3> 0.100705f
C194 XA20/CNO XA6/EN 0.457818f
C195 XA20/XA9/A CK_SAMPLE 0.169353f
C196 XA5/CEO XA4/CEO 0.431793f
C197 AVSS XA2/EN 0.296958f
C198 SARP AVSS 0.540564f
C199 AVSS XA0/DONE 0.27339f
C200 XA20/CPO XA2/CN1 0.255235f
C201 XA20/CNO XA2/EN 0.457819f
C202 DONE XA7/XA9/B 0.27523f
C203 D<1> AVSS 1.876198f
C204 CK_SAMPLE_BSSW AVSS 0.75049f
C205 XA0/CN0 XA0/CP0 3.564212f
C206 SARN SAR_IN 0.271831f
C207 D<5> D<6> 1.055163f
C208 XA1/EN VREF 0.175304f
C209 AVSS XA20/CNO 2.172184f
C210 XA0/CP0 XA1/CN1 0.139477f
C211 XA2/CN0 XA2/CP0 3.180098f
C212 SARN XB2/M4/G 0.24502f
C213 XA0/CP0 D<6> 0.81476f
C214 VREF XA6/EN 0.175304f
C215 XB2/XA3/B AVSS 1.491396f
C216 XA20/CNO XA7/XA4/A 0.304482f
C217 XA3/CN0 XA3/CP0 0.125928f
C218 XA2/CN1 XA2/CP0 0.110086f
C219 XB2/XA4/GNG AVSS 1.208553f
C220 XA5/CN0 XA5/CP0 0.125928f
C221 SARN SARP 5.1717f
C222 XA6/DONE AVSS 0.2733f
C223 SARN AVSS 3.513515f
C224 XA1/CP0 XA2/CP0 1.213936f
C225 XA4/EN XA3/CN0 0.13801f
C226 AVDD XA1/EN 0.791991f
C227 VREF XA2/EN 0.175304f
C228 XA6/EN XA5/CN0 0.13801f
C229 AVSS VREF 1.049192f
C230 AVDD XA6/EN 0.11184f
C231 XA20/CNO XA4/XA4/A 0.212166f
C232 D<5> D<4> 0.356702f
C233 AVDD XA2/EN 0.11184f
C234 XA0/CP0 D<7> 0.111006f
C235 AVSS XA5/CN0 0.234223f
C236 SARN XB2/XA4/GNG 1.624341f
C237 XA0/XA2/A EN 0.11426f
C238 AVDD AVSS 7.430067f
C239 XA0/CP0 D<4> 0.207798f
C240 CK_SAMPLE_BSSW AVDD 14.874317f
C241 AVDD XA20/CNO 2.72258f
C242 XA20/CPO XA1/CN1 0.267213f
C243 EN D<7> 0.334727f
C244 AVSS XA2/DONE 0.2733f
C245 AVDD XB2/XA3/B 0.185337f
C246 XA6/CN0 AVSS 0.279681f
C247 EN XA1/XA2/A 0.11418f
C248 XA2/CN0 XA3/CN0 2.194395f
C249 XA6/XA2/A EN 0.11426f
C250 XA6/CN0 D<1> 2.256405f
C251 XA0/CN0 XA2/CP0 1.220085f
C252 D<5> AVSS 1.873407f
C253 D<4> D<3> 0.665607f
C254 AVDD VREF 15.778251f
C255 XA1/EN EN 0.315013f
C256 XA0/CEIN XB2/M4/G 0.111673f
C257 SARP XA0/CP0 0.107476f
C258 AVSS XA0/CP0 0.207167f
C259 EN XA6/EN 0.235384f
C260 XA1/CEO XA1/XA11/A 0.13078f
C261 XA3/CEO XA3/XA11/A 0.13078f
C262 SARP XA0/CEIN 0.431405f
C263 XA0/CEIN AVSS 2.00975f
C264 AVSS XA0/CEO 0.267201f
C265 XA20/CPO D<7> 0.239708f
C266 AVDD XA5/CN0 2.476604f
C267 XA1/CEO AVSS 0.43736f
C268 EN XA2/EN 0.235383f
C269 XA7/CEO AVSS 0.539406f
C270 XA0/CEIN CK_SAMPLE_BSSW 6.834396f
C271 XA0/CP1 XA2/CN1 1.265362f
C272 AVSS EN 1.655709f
C273 XA7/XA9/MN1/a_324_334# 0 0.360407f
C274 XA7/XA9/MN0/a_324_n18# 0 0.360407f
C275 XA7/XA9/A 0 1.250075f
C276 XA7/XA7/MN0/a_324_n18# 0 0.360407f
C277 XA7/XA8/MN0/a_324_n18# 0 0.360407f
C278 XA7/XA9/B 0 1.158058f
C279 XA7/XA6/MN0/a_324_n18# 0 0.360407f
C280 XA7/XA4/A 0 2.621765f
C281 XA7/XA4/MN0/a_324_n18# 0 0.360407f
C282 XA7/CP0 0 2.4163f
C283 XA7/CN0 0 0.312365f
C284 XA7/XA5/MN0/a_324_n18# 0 0.360407f
C285 XA7/CN1 0 2.428168f
C286 D<0> 0 0.412798f
C287 XA7/XA3/MN0/a_324_n18# 0 0.360407f
C288 XA7/XA2/A 0 2.030764f
C289 XA7/XA2/MN0/a_324_n18# 0 0.360407f
C290 XA7/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C291 XA7/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C292 XA7/XA1/XA2/Y 0 1.060197f
C293 XA7/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C294 XA7/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C295 XA7/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C296 XA7/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C297 XA7/XA1/XA1/MP3/G 0 0.827484f
C298 XA7/XA1/XA1/MN2/S 0 0.200627f
C299 XA7/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C300 XA7/ENO 0 1.582724f
C301 XA7/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C302 XA7/XA13/MN1/a_324_334# 0 0.422f
C303 XA7/XA12/MN0/a_324_n18# 0 0.360407f
C304 XA7/XA13/MN1/a_324_n18# 0 0.360407f
C305 XA7/XA12/A 0 0.755669f
C306 XA7/XA11/MN0/a_324_n18# 0 0.360407f
C307 XA6/CEO 0 1.009021f
C308 XA7/XA11/A 0 0.662715f
C309 XA7/XA9/Y 0 0.718246f
C310 XA6/XA9/MN1/a_324_334# 0 0.360407f
C311 XA6/XA9/MN0/a_324_n18# 0 0.360407f
C312 XA6/XA9/A 0 1.250075f
C313 XA6/DONE 0 0.13094f
C314 XA6/XA7/MN0/a_324_n18# 0 0.360407f
C315 XA6/XA8/MN0/a_324_n18# 0 0.360407f
C316 XA6/XA9/B 0 1.158058f
C317 XA6/XA6/MN0/a_324_n18# 0 0.360407f
C318 XA6/XA4/A 0 2.621765f
C319 XA6/XA4/MN0/a_324_n18# 0 0.360407f
C320 XA6/CP0 0 2.4163f
C321 XA6/CN0 0 4.160099f
C322 XA6/XA5/MN0/a_324_n18# 0 0.360407f
C323 XA6/CN1 0 2.428168f
C324 D<1> 0 4.424545f
C325 XA6/XA3/MN0/a_324_n18# 0 0.360407f
C326 XA6/XA2/A 0 2.030764f
C327 XA6/XA2/MN0/a_324_n18# 0 0.360407f
C328 XA6/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C329 XA6/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C330 XA6/XA1/XA2/Y 0 1.060197f
C331 XA6/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C332 XA6/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C333 XA6/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C334 XA6/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C335 XA6/XA1/XA1/MP3/G 0 0.827484f
C336 XA6/XA1/XA1/MN2/S 0 0.200627f
C337 XA6/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C338 XA7/EN 0 3.856368f
C339 XA6/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C340 XA6/XA13/MN1/a_324_334# 0 0.422f
C341 XA6/XA12/MN0/a_324_n18# 0 0.360407f
C342 XA6/XA13/MN1/a_324_n18# 0 0.360407f
C343 XA6/XA12/A 0 0.755669f
C344 XA6/XA11/MN0/a_324_n18# 0 0.360407f
C345 XA5/CEO 0 1.104751f
C346 XA6/XA11/A 0 0.662715f
C347 XA6/XA9/Y 0 0.718246f
C348 XA5/XA9/MN1/a_324_334# 0 0.360407f
C349 XA5/XA9/MN0/a_324_n18# 0 0.360407f
C350 XA5/XA9/A 0 1.250075f
C351 XA5/DONE 0 0.123486f
C352 XA5/XA7/MN0/a_324_n18# 0 0.360407f
C353 XA5/XA8/MN0/a_324_n18# 0 0.360407f
C354 XA5/XA9/B 0 1.158058f
C355 XA5/XA6/MN0/a_324_n18# 0 0.360407f
C356 XA5/XA4/A 0 2.621765f
C357 XA5/XA4/MN0/a_324_n18# 0 0.360407f
C358 XA5/CP0 0 2.4163f
C359 XA5/CN0 0 3.052303f
C360 XA5/XA5/MN0/a_324_n18# 0 0.360407f
C361 XA5/CN1 0 2.428168f
C362 D<2> 0 3.706573f
C363 XA5/XA3/MN0/a_324_n18# 0 0.360407f
C364 XA5/XA2/A 0 2.030764f
C365 XA5/XA2/MN0/a_324_n18# 0 0.360407f
C366 XA5/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C367 XA5/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C368 XA5/XA1/XA2/Y 0 1.060197f
C369 XA5/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C370 XA5/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C371 XA5/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C372 XA5/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C373 XA5/XA1/XA1/MP3/G 0 0.827484f
C374 XA5/XA1/XA1/MN2/S 0 0.200627f
C375 XA5/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C376 XA6/EN 0 3.679756f
C377 XA5/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C378 XA5/XA13/MN1/a_324_334# 0 0.422f
C379 XA5/XA12/MN0/a_324_n18# 0 0.360407f
C380 XA5/XA13/MN1/a_324_n18# 0 0.360407f
C381 XA5/XA12/A 0 0.755669f
C382 XA5/XA11/MN0/a_324_n18# 0 0.360407f
C383 XA4/CEO 0 1.086041f
C384 XA5/XA11/A 0 0.662715f
C385 XA5/XA9/Y 0 0.718246f
C386 XA4/XA9/MN1/a_324_334# 0 0.360407f
C387 XA4/XA9/MN0/a_324_n18# 0 0.360407f
C388 XA4/XA9/A 0 1.250075f
C389 XA4/DONE 0 0.13094f
C390 XA4/XA7/MN0/a_324_n18# 0 0.360407f
C391 XA4/XA8/MN0/a_324_n18# 0 0.360407f
C392 XA4/XA9/B 0 1.158058f
C393 XA4/XA6/MN0/a_324_n18# 0 0.360407f
C394 XA4/XA4/A 0 2.621765f
C395 XA4/XA4/MN0/a_324_n18# 0 0.360407f
C396 XA4/CP0 0 2.4163f
C397 XA4/CN0 0 2.237548f
C398 XA4/XA5/MN0/a_324_n18# 0 0.360407f
C399 XA4/CN1 0 2.428168f
C400 D<3> 0 2.560026f
C401 XA4/XA3/MN0/a_324_n18# 0 0.360407f
C402 XA4/XA2/A 0 2.030764f
C403 XA4/XA2/MN0/a_324_n18# 0 0.360407f
C404 XA4/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C405 XA4/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C406 XA4/XA1/XA2/Y 0 1.060197f
C407 XA4/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C408 XA4/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C409 XA4/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C410 XA4/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C411 XA4/XA1/XA1/MP3/G 0 0.827484f
C412 XA4/XA1/XA1/MN2/S 0 0.200627f
C413 XA4/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C414 XA5/EN 0 3.635208f
C415 XA4/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C416 XA4/XA13/MN1/a_324_334# 0 0.422f
C417 XA4/XA12/MN0/a_324_n18# 0 0.360407f
C418 XA4/XA13/MN1/a_324_n18# 0 0.360407f
C419 XA4/XA12/A 0 0.755669f
C420 XA4/XA11/MN0/a_324_n18# 0 0.360407f
C421 XA3/CEO 0 1.107611f
C422 XA4/XA11/A 0 0.662715f
C423 XA4/XA9/Y 0 0.718246f
C424 XA3/XA9/MN1/a_324_334# 0 0.360407f
C425 XA3/XA9/MN0/a_324_n18# 0 0.360407f
C426 XA3/XA9/A 0 1.250075f
C427 XA3/DONE 0 0.123486f
C428 XA3/XA7/MN0/a_324_n18# 0 0.360407f
C429 XA3/XA8/MN0/a_324_n18# 0 0.360407f
C430 XA3/XA9/B 0 1.158058f
C431 XA3/XA6/MN0/a_324_n18# 0 0.360407f
C432 XA3/XA4/A 0 2.621765f
C433 XA3/XA4/MN0/a_324_n18# 0 0.360407f
C434 XA3/CP0 0 2.4163f
C435 XA3/CN0 0 3.224855f
C436 XA3/XA5/MN0/a_324_n18# 0 0.360407f
C437 XA3/CN1 0 2.428168f
C438 D<4> 0 3.08566f
C439 XA3/XA3/MN0/a_324_n18# 0 0.360407f
C440 XA3/XA2/A 0 2.030764f
C441 XA3/XA2/MN0/a_324_n18# 0 0.360407f
C442 XA3/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C443 XA3/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C444 XA3/XA1/XA2/Y 0 1.060197f
C445 XA3/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C446 XA3/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C447 XA3/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C448 XA3/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C449 XA3/XA1/XA1/MP3/G 0 0.827484f
C450 XA3/XA1/XA1/MN2/S 0 0.200627f
C451 XA3/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C452 XA4/EN 0 3.720665f
C453 XA3/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C454 XA3/XA13/MN1/a_324_334# 0 0.422f
C455 XA3/XA12/MN0/a_324_n18# 0 0.360407f
C456 XA3/XA13/MN1/a_324_n18# 0 0.360407f
C457 XA3/XA12/A 0 0.755669f
C458 XA3/XA11/MN0/a_324_n18# 0 0.360407f
C459 XA2/CEO 0 1.085281f
C460 XA3/XA11/A 0 0.662715f
C461 XA3/XA9/Y 0 0.718246f
C462 XA2/XA9/MN1/a_324_334# 0 0.360407f
C463 XA2/XA9/MN0/a_324_n18# 0 0.360407f
C464 XA2/XA9/A 0 1.250075f
C465 XA2/DONE 0 0.13094f
C466 XA2/XA7/MN0/a_324_n18# 0 0.360407f
C467 XA2/XA8/MN0/a_324_n18# 0 0.360407f
C468 XA2/XA9/B 0 1.158058f
C469 XA2/XA6/MN0/a_324_n18# 0 0.360407f
C470 XA2/XA4/A 0 2.621765f
C471 XA2/XA4/MN0/a_324_n18# 0 0.360407f
C472 XA2/CP0 0 4.49437f
C473 XA2/CN0 0 2.820252f
C474 XA2/XA5/MN0/a_324_n18# 0 0.360407f
C475 XA2/CN1 0 6.112935f
C476 XA2/XA3/MN0/a_324_n18# 0 0.360407f
C477 XA2/XA2/A 0 2.030764f
C478 XA2/XA2/MN0/a_324_n18# 0 0.360407f
C479 XA2/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C480 XA2/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C481 XA2/XA1/XA2/Y 0 1.060197f
C482 XA2/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C483 XA2/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C484 XA2/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C485 XA2/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C486 XA2/XA1/XA1/MP3/G 0 0.827484f
C487 XA2/XA1/XA1/MN2/S 0 0.200627f
C488 XA2/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C489 XA3/EN 0 3.784028f
C490 XA2/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C491 XA2/XA13/MN1/a_324_334# 0 0.422f
C492 XA2/XA12/MN0/a_324_n18# 0 0.360407f
C493 XA2/XA13/MN1/a_324_n18# 0 0.360407f
C494 XA2/XA12/A 0 0.755669f
C495 XA2/XA11/MN0/a_324_n18# 0 0.360407f
C496 XA1/CEO 0 1.104751f
C497 XA2/XA11/A 0 0.662715f
C498 XA2/XA9/Y 0 0.718246f
C499 XA1/XA9/MN1/a_324_334# 0 0.360407f
C500 XA1/XA9/MN0/a_324_n18# 0 0.360407f
C501 XA1/XA9/A 0 1.250075f
C502 XA1/DONE 0 0.123486f
C503 XA1/XA7/MN0/a_324_n18# 0 0.360407f
C504 XA1/XA8/MN0/a_324_n18# 0 0.360407f
C505 XA1/XA9/B 0 1.158058f
C506 XA1/XA6/MN0/a_324_n18# 0 0.360407f
C507 XA1/XA4/A 0 2.621765f
C508 XA1/XA4/MN0/a_324_n18# 0 0.360407f
C509 XA1/CP0 0 4.486094f
C510 XA1/CN0 0 2.798774f
C511 XA1/XA5/MN0/a_324_n18# 0 0.360407f
C512 XA1/CN1 0 4.70217f
C513 D<6> 0 2.989828f
C514 XA1/XA3/MN0/a_324_n18# 0 0.360407f
C515 XA1/XA2/A 0 2.030764f
C516 XA1/XA2/MN0/a_324_n18# 0 0.360407f
C517 XA1/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C518 XA1/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C519 XA1/XA1/XA2/Y 0 1.060197f
C520 XA1/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C521 XA1/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C522 XA1/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C523 XA1/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C524 XA1/XA1/XA1/MP3/G 0 0.827484f
C525 XA1/XA1/XA1/MN2/S 0 0.200627f
C526 XA1/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C527 XA2/EN 0 3.720665f
C528 XA1/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C529 XA1/XA13/MN1/a_324_334# 0 0.422f
C530 XA1/XA12/MN0/a_324_n18# 0 0.360407f
C531 XA1/XA13/MN1/a_324_n18# 0 0.360407f
C532 XA1/XA12/A 0 0.755669f
C533 XA1/XA11/MN0/a_324_n18# 0 0.360407f
C534 XA0/CEO 0 1.083361f
C535 XA1/XA11/A 0 0.662715f
C536 XA1/XA9/Y 0 0.718246f
C537 XB2/XA7/MN1/a_324_n18# 0 0.359583f
C538 XB2/XA5b/MN1/a_324_n18# 0 0.422415f
C539 XB2/XA1/Y 0 0.690197f
C540 XB2/CKN 0 1.768971f
C541 XB2/XA4/MN0/a_324_n18# 0 0.359583f
C542 XB2/XA5/MN1/a_324_334# 0 0.422f
C543 XB2/XA3/MP0/S 0 0.743486f
C544 XB2/XA3/MN0/a_324_n18# 0 0.359583f
C545 XB2/XA2/MP0/G 0 0.708335f
C546 XB2/XA7/MN1/a_324_334# 0 0.359583f
C547 XB2/XA5/MN1/a_324_n18# 0 0.360407f
C548 XB2/XA1/MP0/G 0 0.788614f
C549 XB2/XA4/MN1/a_324_334# 0 0.359583f
C550 XB2/XA0/MN0/a_324_n18# 0 0.359583f
C551 XB2/M8/a_324_n18# 0 0.356977f
C552 XB2/M8/a_324_334# 0 0.422f
C553 XB2/M6/a_324_n18# 0 0.356977f
C554 XB2/M7/a_324_n18# 0 0.356977f
C555 XB2/XA3/B 0 54.41209f
C556 XB2/XA4/GNG 0 53.065117f
C557 XB2/M5/a_324_n18# 0 0.356977f
C558 XB2/M3/a_324_n18# 0 0.356977f
C559 XB2/M4/a_324_n18# 0 0.356977f
C560 XB2/M4/G 0 2.475647f
C561 SAR_IN 0 1.184896f
C562 XB2/M1/a_324_n18# 0 0.422415f
C563 XB2/M2/a_324_n18# 0 0.356977f
C564 XA0/XA9/MN1/a_324_334# 0 0.360407f
C565 XA0/XA9/MN0/a_324_n18# 0 0.360407f
C566 XA0/XA9/A 0 1.250075f
C567 XA0/DONE 0 0.134046f
C568 XA0/XA7/MN0/a_324_n18# 0 0.360407f
C569 XA0/XA8/MN0/a_324_n18# 0 0.360407f
C570 XA0/XA9/B 0 1.158058f
C571 CK_SAMPLE 0 15.793598f
C572 XA0/XA6/MN0/a_324_n18# 0 0.360407f
C573 XA0/XA4/A 0 2.621765f
C574 XA0/XA4/MN0/a_324_n18# 0 0.360407f
C575 XA0/CP0 0 8.48089f
C576 XA0/XA5/MN0/a_324_n18# 0 0.360407f
C577 VREF 0 27.717136f
C578 D<7> 0 7.541619f
C579 XA0/XA3/MN0/a_324_n18# 0 0.360407f
C580 XA0/XA2/A 0 2.030764f
C581 XA0/XA2/MN0/a_324_n18# 0 0.360407f
C582 XA20/CNO 0 12.667546f
C583 XA0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C584 EN 0 4.718864f
C585 XA0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C586 XA0/XA1/XA2/Y 0 1.060197f
C587 XA0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C588 XA0/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C589 XA20/CPO 0 11.091676f
C590 XA0/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C591 XA0/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C592 XA0/XA1/XA1/MP3/G 0 0.827484f
C593 XA0/XA1/XA1/MN2/S 0 0.200627f
C594 XA0/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C595 XA1/EN 0 3.794638f
C596 XA0/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C597 AVDD 0 0.517971p
C598 XA0/XA13/MN1/a_324_334# 0 0.422f
C599 XA0/XA12/MN0/a_324_n18# 0 0.360407f
C600 XA0/XA13/MN1/a_324_n18# 0 0.360407f
C601 XA0/XA12/A 0 0.755669f
C602 XA0/XA11/MN0/a_324_n18# 0 0.360407f
C603 XA0/XA11/A 0 0.662715f
C604 XA0/XA9/Y 0 0.718246f
C605 XB1/XA7/MN1/a_324_n18# 0 0.359583f
C606 AVSS 0 0.14072p
C607 XB1/XA5b/MN1/a_324_n18# 0 0.422415f
C608 XB1/XA1/Y 0 0.690197f
C609 XB1/CKN 0 1.768971f
C610 XB1/XA4/MN0/a_324_n18# 0 0.359583f
C611 XB1/XA5/MN1/a_324_334# 0 0.422f
C612 XB1/XA3/MP0/S 0 0.743486f
C613 XB1/XA3/MN0/a_324_n18# 0 0.359583f
C614 XB1/XA2/MP0/G 0 0.708335f
C615 XB1/XA7/MN1/a_324_334# 0 0.359583f
C616 XB1/XA5/MN1/a_324_n18# 0 0.360407f
C617 XB1/XA1/MP0/G 0 0.788614f
C618 XB1/XA4/MN1/a_324_334# 0 0.359583f
C619 CK_SAMPLE_BSSW 0 3.70264f
C620 XB1/XA0/MN0/a_324_n18# 0 0.359583f
C621 XB1/M8/a_324_n18# 0 0.356977f
C622 XB1/M8/a_324_334# 0 0.422f
C623 XB1/M6/a_324_n18# 0 0.356977f
C624 XB1/M7/a_324_n18# 0 0.356977f
C625 XB1/XA3/B 0 54.41209f
C626 XB1/XA4/GNG 0 53.065117f
C627 XA0/CEIN 0 19.901903f
C628 XB1/M5/a_324_n18# 0 0.356977f
C629 XB1/M3/a_324_n18# 0 0.356977f
C630 XB1/M4/a_324_n18# 0 0.356977f
C631 XB1/M4/G 0 2.475647f
C632 SAR_IP 0 1.184896f
C633 XB1/M1/a_324_n18# 0 0.422415f
C634 XB1/M2/a_324_n18# 0 0.356977f
C635 XA20/XA9/MN0/a_324_n18# 0 0.360407f
C636 XA20/XA3/CO 0 2.703497f
C637 XA20/XA2/MN6/a_324_334# 0 0.360407f
C638 XA20/XA3a/A 0 2.536943f
C639 XA20/XA3/MN0/a_324_n18# 0 0.360407f
C640 XA20/XA3a/MN0/a_324_n18# 0 0.360407f
C641 XA20/XA4/MN0/a_324_n18# 0 0.360407f
C642 XA20/XA4/MP0/S 0 0.397005f
C643 SARN 0 29.964926f
C644 XA20/XA3/N2 0 0.234927f
C645 XA20/XA9/Y 0 3.176436f
C646 XA20/XA2/N2 0 0.234927f
C647 XA20/XA2/MN0/a_324_n18# 0 0.360407f
C648 XA20/XA3/N1 0 0.905385f
C649 SARP 0 30.549707f
C650 XA20/XA1/MN0/a_324_n18# 0 0.360407f
C651 XA20/XA1/MP0/S 0 0.397005f
C652 XA20/XA9/A 0 3.508213f
C653 XA20/XA0/MN1/a_324_n18# 0 0.422415f
C654 XA20/XA13/MN1/a_324_n18# 0 0.360407f
C655 XA20/XA13/MN1/a_324_334# 0 0.422f
C656 XA7/CEO 0 1.316615f
C657 XA20/XA12/MN0/a_324_n18# 0 0.360407f
C658 XA20/XA11/MN0/a_324_n18# 0 0.360407f
C659 DONE 0 0.902344f
C660 XA20/XA9/MN0/a_324_334# 0 0.360407f
C661 XA20/XA12/Y 0 0.623343f
C662 XA20/XA11/Y 0 0.759616f
C663 XDAC2/XC32a<0>/XRES2/B 0 3.1129f
C664 XDAC2/XC32a<0>/XRES4/B 0 3.516117f
C665 XDAC2/XC32a<0>/XRES8/B 0 3.933522f
C666 XDAC2/XC32a<0>/XRES16/B 0 4.664508f
C667 XDAC2/XC32a<0>/XRES1B/B 0 2.892833f
C668 XDAC2/XC32a<0>/XRES1A/B 0 1.735354f
C669 XDAC2/XC1/XRES2/B 0 3.1129f
C670 XDAC2/XC1/XRES4/B 0 3.516117f
C671 XDAC2/XC1/XRES8/B 0 3.933522f
C672 XDAC2/XC1/XRES16/B 0 4.664508f
C673 XDAC2/XC1/XRES1B/B 0 2.892833f
C674 XDAC2/XC1/XRES1A/B 0 1.735354f
C675 XA0/CN0 0 6.776559f
C676 XDAC2/XC0/XRES2/B 0 3.1129f
C677 XDAC2/XC0/XRES4/B 0 3.516117f
C678 XDAC2/XC0/XRES8/B 0 3.933522f
C679 XDAC2/XC0/XRES16/B 0 4.664508f
C680 XDAC2/XC0/XRES1B/B 0 2.892833f
C681 XDAC2/XC0/XRES1A/B 0 1.735354f
C682 XDAC2/X16ab/XRES2/B 0 3.1129f
C683 XDAC2/X16ab/XRES4/B 0 3.516117f
C684 XDAC2/X16ab/XRES8/B 0 3.933522f
C685 XDAC2/X16ab/XRES16/B 0 4.664508f
C686 XDAC2/X16ab/XRES1B/B 0 2.892833f
C687 XDAC2/X16ab/XRES1A/B 0 1.735354f
C688 XDAC1/XC32a<0>/XRES2/B 0 3.1129f
C689 XDAC1/XC32a<0>/XRES4/B 0 3.516117f
C690 XDAC1/XC32a<0>/XRES8/B 0 3.933522f
C691 XDAC1/XC32a<0>/XRES16/B 0 4.664508f
C692 XDAC1/XC32a<0>/XRES1B/B 0 2.892833f
C693 XDAC1/XC32a<0>/XRES1A/B 0 1.735354f
C694 XDAC1/XC1/XRES2/B 0 3.1129f
C695 XDAC1/XC1/XRES4/B 0 3.516117f
C696 XDAC1/XC1/XRES8/B 0 3.933522f
C697 XDAC1/XC1/XRES16/B 0 4.664508f
C698 XDAC1/XC1/XRES1B/B 0 2.892833f
C699 XDAC1/XC1/XRES1A/B 0 1.735354f
C700 XDAC1/XC0/XRES2/B 0 3.1129f
C701 XDAC1/XC0/XRES4/B 0 3.516117f
C702 XDAC1/XC0/XRES8/B 0 3.933522f
C703 XDAC1/XC0/XRES16/B 0 4.664508f
C704 XDAC1/XC0/XRES1B/B 0 2.892833f
C705 XDAC1/XC0/XRES1A/B 0 1.735354f
C706 D<5> 0 4.36517f
C707 XDAC1/X16ab/XRES2/B 0 3.1129f
C708 XDAC1/X16ab/XRES4/B 0 3.516117f
C709 XDAC1/X16ab/XRES8/B 0 3.933522f
C710 XDAC1/X16ab/XRES16/B 0 4.664508f
C711 XDAC1/X16ab/XRES1B/B 0 2.892833f
C712 XDAC1/X16ab/XRES1A/B 0 1.735354f
C713 XA0/CP1 0 4.930175f
.ends

.subckt SUNSAR_IVTRIX1_CV CN AVDD AVSS MN1/a_324_334# C Y BULKP MP0/a_216_n18# MP1/a_216_334#
+ A MN0/a_324_n18# VSUBS
XMP0 MP1/S A AVDD BULKP MP0/a_216_n18# CN VSUBS SUNSAR_PCHDL
XMP1 Y CN MP1/S BULKP A MP1/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 MN1/S A AVSS VSUBS MN0/a_324_n18# C SUNSAR_NCHDL
XMN1 Y C MN1/S VSUBS A MN1/a_324_334# SUNSAR_NCHDL
C0 BULKP A -0.231483f
C1 BULKP CN -0.345553f
C2 BULKP AVDD 0.123213f
C3 AVDD VSUBS 0.259844f
C4 AVSS VSUBS 0.395374f
C5 C VSUBS 0.372036f
C6 Y VSUBS 0.262859f
C7 MN1/a_324_334# VSUBS 0.422f
C8 A VSUBS 0.569283f
C9 MN0/a_324_n18# VSUBS 0.422415f
C10 BULKP VSUBS 3.597147f
.ends

.subckt SUNSAR_DFQNX1_CV Q QN XA7/C CK D AVDD AVSS
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA1 AVDD AVSS XA7/C XA1/MP0/a_216_n18# XA2/MP0/a_216_n18# AVDD CK XA1/MN0/a_324_n18#
+ AVSS XA2/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA2 AVDD AVSS XA6/C XA2/MP0/a_216_n18# XA3/MP0/a_216_n18# AVDD XA7/C XA2/MN0/a_324_n18#
+ AVSS XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA3 XA6/C AVDD AVSS XA4/MN0/a_324_n18# XA7/C XA5/A AVDD XA3/MP0/a_216_n18# XA4/MP0/a_216_n18#
+ D XA3/MN0/a_324_n18# AVSS SUNSAR_IVTRIX1_CV
XXA4 XA7/C AVDD AVSS XA5/MN0/a_324_n18# XA6/C XA5/A AVDD XA4/MP0/a_216_n18# XA5/MP0/a_216_n18#
+ XA6/A XA4/MN0/a_324_n18# AVSS SUNSAR_IVTRIX1_CV
XXA5 AVDD AVSS XA6/A XA5/MP0/a_216_n18# XA6/MP0/a_216_n18# AVDD XA5/A XA5/MN0/a_324_n18#
+ AVSS XA6/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA6 XA7/C AVDD AVSS XA7/MN0/a_324_n18# XA6/C QN AVDD XA6/MP0/a_216_n18# XA7/MP0/a_216_n18#
+ XA6/A XA6/MN0/a_324_n18# AVSS SUNSAR_IVTRIX1_CV
XXA7 XA6/C AVDD AVSS XA8/MN0/a_324_n18# XA7/C QN AVDD XA7/MP0/a_216_n18# XA8/MP0/a_216_n18#
+ Q XA7/MN0/a_324_n18# AVSS SUNSAR_IVTRIX1_CV
XXA8 AVDD AVSS Q XA8/MP0/a_216_n18# XA8/MP0/a_216_334# AVDD QN XA8/MN0/a_324_n18#
+ AVSS XA8/MN0/a_324_334# SUNSAR_IVX1_CV
C0 AVDD XA6/MP0/a_216_n18# -0.315634f
C1 AVDD XA5/MP0/a_216_n18# -0.313035f
C2 XA6/C XA5/A 0.400241f
C3 XA6/C XA6/A 0.511866f
C4 XA6/C Q 0.188983f
C5 XA6/C XA7/C 0.555229f
C6 AVDD XA6/C 0.894074f
C7 AVSS QN 0.208618f
C8 AVDD XA3/MP0/a_216_n18# -0.313035f
C9 AVDD XA7/MP0/a_216_n18# -0.314611f
C10 CK XA7/C 0.13667f
C11 AVSS XA5/A 0.31114f
C12 Q QN 0.164289f
C13 XA7/C QN 0.28651f
C14 AVDD QN 0.152707f
C15 XA6/A XA5/A 0.225387f
C16 AVSS XA7/C 0.523585f
C17 XA7/C XA6/A 0.41755f
C18 AVDD XA5/A 0.149071f
C19 AVDD XA6/A 0.50597f
C20 AVDD XA2/MP0/a_216_n18# -0.31496f
C21 XA7/C Q 0.128539f
C22 AVDD Q 0.337452f
C23 AVDD XA7/C 1.562268f
C24 XA6/C D 0.110712f
C25 AVDD XA8/MP0/a_216_n18# -0.312509f
C26 XA1/MP0/a_216_n18# AVDD -0.311986f
C27 D XA7/C 0.117769f
C28 AVDD XA4/MP0/a_216_n18# -0.313035f
C29 AVSS XA6/C 0.2601f
C30 XA7/C 0 2.352415f
C31 QN 0 0.966414f
C32 Q 0 0.838602f
C33 XA8/MN0/a_324_334# 0 0.422f
C34 XA8/MN0/a_324_n18# 0 0.360407f
C35 XA7/MN0/a_324_n18# 0 0.360407f
C36 XA6/MN0/a_324_n18# 0 0.360407f
C37 XA5/A 0 0.896691f
C38 XA6/A 0 1.098676f
C39 XA5/MN0/a_324_n18# 0 0.360407f
C40 XA4/MN0/a_324_n18# 0 0.360407f
C41 D 0 0.487386f
C42 XA3/MN0/a_324_n18# 0 0.360407f
C43 XA6/C 0 1.328497f
C44 XA2/MN0/a_324_n18# 0 0.360407f
C45 CK 0 0.515118f
C46 XA1/MN0/a_324_n18# 0 0.360407f
C47 AVSS 0 -0.115052f
C48 XA0/MN1/a_324_n18# 0 0.422415f
C49 AVDD 0 18.699612f
.ends

.subckt SUNSAR_ORX1_CV AVDD AVSS B XA1/MP0/a_216_n18# XA1/MN0/a_324_n18# XA2/MP0/a_216_334#
+ A BULKP XA2/MN0/a_324_334# VSUBS Y
XXA1 AVDD AVSS XA2/MN0/a_324_n18# B BULKP XA1/MP0/a_216_n18# XA2/A XA2/MP0/a_216_n18#
+ A XA1/MN0/a_324_n18# VSUBS SUNSAR_NRX1_CV
XXA2 BULKP AVSS Y XA2/MP0/a_216_n18# XA2/MP0/a_216_334# AVDD XA2/A XA2/MN0/a_324_n18#
+ VSUBS XA2/MN0/a_324_334# SUNSAR_IVX1_CV
C0 BULKP XA2/MP0/a_216_n18# -0.310513f
C1 B XA2/A 0.110841f
C2 Y VSUBS 0.217477f
C3 XA2/MN0/a_324_n18# VSUBS 0.357149f
C4 XA2/MN0/a_324_334# VSUBS 0.422f
C5 AVDD VSUBS 0.321354f
C6 AVSS VSUBS 0.551073f
C7 XA2/A VSUBS 0.902459f
C8 XA1/MN0/a_324_n18# VSUBS 0.422415f
C9 B VSUBS 0.472321f
C10 BULKP VSUBS 5.173117f
C11 A VSUBS 0.541859f
.ends

.subckt SUNSAR_BFX1_CV Y AVDD AVSS MN1/a_324_334# MP1/G A BULKP MP0/a_216_n18# MP1/a_216_334#
+ MN0/a_324_n18# VSUBS
XMP0 AVDD A MP1/G BULKP MP0/a_216_n18# MP1/G VSUBS SUNSAR_PCHDL
XMP1 Y MP1/G AVDD BULKP A MP1/a_216_334# VSUBS SUNSAR_PCHDL
XMN0 AVSS A MP1/G VSUBS MN0/a_324_n18# MP1/G SUNSAR_NCHDL
XMN1 Y MP1/G AVSS VSUBS A MN1/a_324_334# SUNSAR_NCHDL
C0 BULKP MP1/G -0.189656f
C1 A MP1/G 0.120372f
C2 A BULKP -0.246947f
C3 AVSS VSUBS 0.330762f
C4 Y VSUBS 0.213901f
C5 MN1/a_324_334# VSUBS 0.422f
C6 AVDD VSUBS 0.225252f
C7 MN0/a_324_n18# VSUBS 0.422415f
C8 MP1/G VSUBS 0.888781f
C9 BULKP VSUBS 3.596797f
C10 A VSUBS 0.536396f
.ends

.subckt SUNSAR_ANX1_CV B XA1/MP0/a_216_n18# XA2/A XA1/MN0/a_324_n18# XA2/MP0/a_216_334#
+ A BULKP XA2/MN0/a_324_334# AVDD AVSS VSUBS Y
XXA1 XA2/A AVDD AVSS XA2/MN0/a_324_n18# B A BULKP XA1/MP0/a_216_n18# XA2/MP0/a_216_n18#
+ XA1/MN0/a_324_n18# VSUBS SUNSAR_NDX1_CV
XXA2 BULKP AVSS Y XA2/MP0/a_216_n18# XA2/MP0/a_216_334# AVDD XA2/A XA2/MN0/a_324_n18#
+ VSUBS XA2/MN0/a_324_334# SUNSAR_IVX1_CV
C0 XA2/MP0/a_216_n18# BULKP -0.310513f
C1 Y VSUBS 0.219919f
C2 XA2/MN0/a_324_n18# VSUBS 0.357149f
C3 XA2/MN0/a_324_334# VSUBS 0.422f
C4 AVSS VSUBS 0.513075f
C5 AVDD VSUBS 0.340245f
C6 XA1/MN0/a_324_n18# VSUBS 0.422415f
C7 XA2/A VSUBS 0.881651f
C8 B VSUBS 0.474445f
C9 BULKP VSUBS 5.173117f
C10 A VSUBS 0.541859f
.ends

.subckt SUNSAR_CAPT8B_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN D<7> D<6> D<5> D<4>
+ D<3> D<2> D<1> D<0> DO<7> DO<6> DO<5> DO<4> DO<3> DO<2> DO<1> DO<0> TIE_L DONE AVDD
+ AVSS
XXD09 DO<5> XD09/QN XD09/XA7/C DONE D<5> AVDD AVSS SUNSAR_DFQNX1_CV
XXB07 DO<7> XB07/QN XB07/XA7/C DONE D<7> AVDD AVSS SUNSAR_DFQNX1_CV
XSUNSAR_IVX1_CV_0 AVDD AVSS XA5/B XA1/MP1/a_216_334# XA3/MP0/a_216_n18# AVDD ENABLE
+ XA1/MN1/a_324_334# AVSS XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXI14 DO<0> XI14/QN XI14/XA7/C DONE D<0> AVDD AVSS SUNSAR_DFQNX1_CV
XXG12 DO<2> XG12/QN XG12/XA7/C DONE D<2> AVDD AVSS SUNSAR_DFQNX1_CV
XXE10 DO<4> XE10/QN XE10/XA7/C DONE D<4> AVDD AVSS SUNSAR_DFQNX1_CV
XXC08 DO<6> XC08/QN XC08/XA7/C DONE D<6> AVDD AVSS SUNSAR_DFQNX1_CV
XXA1 AVDD XA1/MN1/a_324_n18# XA1/MN1/a_324_334# XA1/MP1/a_216_334# XA1/MP1/a_216_n18#
+ AVSS SUNSAR_TAPCELLB_CV
XXA2 AVDD AVDD AVSS XA2/MP0/G TIE_L XA2/MP0/a_216_n18# XA2/MP0/a_216_334# XA2/MN0/a_324_n18#
+ AVSS XA2/MN0/a_324_334# SUNSAR_TIEL_CV
XXA5a AVDD AVSS EN XA5a/MP0/a_216_n18# XA5a/MP0/a_216_334# AVDD CK_SAMPLE XA5a/MN0/a_324_n18#
+ AVSS XA5a/MN0/a_324_334# SUNSAR_IVX1_CV
XXA3 AVDD AVSS XA6/B XA3/MP0/a_216_n18# XA4/MP0/a_216_n18# AVDD XA5/B XA3/MN0/a_324_n18#
+ AVSS XA4/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA5 AVDD AVSS XA5/B XA4/MP1/a_216_334# XA4/MN1/a_324_334# XA5a/MP0/a_216_n18# XA6/A
+ AVDD XA5a/MN0/a_324_n18# AVSS CK_SAMPLE SUNSAR_ORX1_CV
XXA4 XA6/A AVDD AVSS XA4/MN1/a_324_334# XA4/MP1/G CKS AVDD XA4/MP0/a_216_n18# XA4/MP1/a_216_334#
+ XA4/MN0/a_324_n18# AVSS SUNSAR_BFX1_CV
XXH13 DO<1> XH13/QN XH13/XA7/C DONE D<1> AVDD AVSS SUNSAR_DFQNX1_CV
XXA6 XA6/B XA5a/MP0/a_216_334# XA6/XA2/A XA5a/MN0/a_324_334# XA2/MP0/a_216_n18# XA6/A
+ AVDD XA2/MN0/a_324_n18# AVDD AVSS AVSS CK_SAMPLE_BSSW SUNSAR_ANX1_CV
XXF11 DO<3> XF11/QN XF11/XA7/C DONE D<3> AVDD AVSS SUNSAR_DFQNX1_CV
C0 DO<0> AVSS 0.192871f
C1 XA5/B XA4/MP1/G 0.138434f
C2 D<4> AVSS 0.301985f
C3 XA5/B XA6/B 0.187691f
C4 DO<7> AVSS 0.186597f
C5 D<3> D<4> 0.12805f
C6 XH13/XA7/C XI14/XA7/C 0.233892f
C7 EN AVSS 0.334598f
C8 DO<3> AVSS 0.187665f
C9 D<5> AVDD 0.137402f
C10 XA5/B CKS 0.210661f
C11 D<5> D<6> 0.12805f
C12 D<5> DONE 0.295113f
C13 DO<2> AVSS 0.187666f
C14 XA4/MP1/a_216_334# AVDD -0.311908f
C15 XG12/XA7/C XF11/XA7/C 0.233892f
C16 TIE_L AVSS 0.167035f
C17 ENABLE AVSS 0.410372f
C18 XA6/B XA6/XA2/A 0.172524f
C19 D<4> AVDD 0.137402f
C20 DO<1> AVSS 0.187666f
C21 EN AVDD 0.458465f
C22 DONE D<4> 0.295113f
C23 D<0> AVSS 0.32707f
C24 EN XA6/B 0.176334f
C25 XA3/MP0/a_216_n18# AVDD -0.311309f
C26 EN CK_SAMPLE 0.28401f
C27 ENABLE AVDD 0.145509f
C28 AVSS DO<4> 0.187665f
C29 XA6/A AVSS 0.540389f
C30 D<2> AVSS 0.301985f
C31 D<3> AVSS 0.301985f
C32 D<0> AVDD 0.142353f
C33 D<0> XI14/XA7/C 0.159126f
C34 D<1> AVSS 0.301985f
C35 D<1> D<2> 0.12805f
C36 DONE D<0> 0.29654f
C37 DO<6> AVSS 0.187666f
C38 XA2/MP0/a_216_n18# AVDD -0.313603f
C39 XA5/B ENABLE 0.10479f
C40 DO<5> AVSS 0.187665f
C41 AVDD AVSS 6.228554f
C42 D<2> AVDD 0.137402f
C43 AVSS D<6> 0.301985f
C44 XC08/XA7/C D<6> 0.159126f
C45 XA4/MP0/a_216_n18# AVDD -0.311772f
C46 D<4> XE10/XA7/C 0.159127f
C47 D<3> AVDD 0.137402f
C48 XA6/A XA6/B 0.223197f
C49 D<7> AVSS 0.290141f
C50 DONE AVSS 7.136209f
C51 DONE D<2> 0.295113f
C52 XA6/B AVSS 0.54117f
C53 XA6/A CK_SAMPLE 0.103062f
C54 XC08/XA7/C XB07/XA7/C 0.233892f
C55 D<1> AVDD 0.137402f
C56 D<3> DONE 0.295113f
C57 CK_SAMPLE AVSS 0.395202f
C58 D<5> XD09/XA7/C 0.159126f
C59 XA6/A CKS 0.198582f
C60 CKS AVSS 1.512398f
C61 D<1> DONE 0.295113f
C62 CK_SAMPLE_BSSW AVSS 0.339545f
C63 XA5a/MP0/a_216_n18# AVDD -0.313603f
C64 XA6/A XA5/B 0.263519f
C65 D<2> XG12/XA7/C 0.159126f
C66 XA5/B AVSS 0.356101f
C67 XA6/B XA5/XA2/A 0.134182f
C68 AVDD D<6> 0.137402f
C69 XA1/MP1/a_216_334# AVDD -0.311986f
C70 CK_SAMPLE XA5/XA2/A 0.123914f
C71 D<3> XF11/XA7/C 0.159126f
C72 D<7> AVDD 0.129858f
C73 DONE AVDD 2.494628f
C74 XA6/B AVDD 0.218203f
C75 DONE D<6> 0.295113f
C76 XD09/XA7/C XE10/XA7/C 0.233892f
C77 CK_SAMPLE AVDD 0.496932f
C78 D<5> AVSS 0.301985f
C79 D<7> DONE 0.292286f
C80 XA6/B XA4/MP1/G 0.300066f
C81 D<7> XB07/XA7/C 0.159126f
C82 CK_SAMPLE_BSSW AVDD 0.508937f
C83 XA5a/MP0/a_216_334# AVDD -0.313603f
C84 CK_SAMPLE XA6/B 0.199415f
C85 D<1> XH13/XA7/C 0.159126f
C86 XF11/XA7/C 0 2.352415f
C87 XF11/QN 0 0.966414f
C88 DO<3> 0 0.963071f
C89 XF11/XA8/MN0/a_324_334# 0 0.422f
C90 XF11/XA8/MN0/a_324_n18# 0 0.360407f
C91 XF11/XA7/MN0/a_324_n18# 0 0.360407f
C92 XF11/XA6/MN0/a_324_n18# 0 0.360407f
C93 XF11/XA5/A 0 0.896691f
C94 XF11/XA6/A 0 1.098676f
C95 XF11/XA5/MN0/a_324_n18# 0 0.360407f
C96 XF11/XA4/MN0/a_324_n18# 0 0.360407f
C97 D<3> 0 0.918631f
C98 XF11/XA3/MN0/a_324_n18# 0 0.360407f
C99 XF11/XA6/C 0 1.328497f
C100 XF11/XA2/MN0/a_324_n18# 0 0.360407f
C101 XF11/XA1/MN0/a_324_n18# 0 0.360407f
C102 XF11/XA0/MN1/a_324_n18# 0 0.422415f
C103 CK_SAMPLE_BSSW 0 0.351307f
C104 XA6/XA2/MN0/a_324_n18# 0 0.360407f
C105 XA2/MN0/a_324_n18# 0 0.359492f
C106 XA5a/MN0/a_324_334# 0 0.359492f
C107 XA6/XA2/A 0 0.871363f
C108 XA6/B 0 1.026139f
C109 XH13/XA7/C 0 2.352415f
C110 XH13/QN 0 0.966414f
C111 DO<1> 0 0.963071f
C112 XH13/XA8/MN0/a_324_334# 0 0.422f
C113 XH13/XA8/MN0/a_324_n18# 0 0.360407f
C114 XH13/XA7/MN0/a_324_n18# 0 0.360407f
C115 XH13/XA6/MN0/a_324_n18# 0 0.360407f
C116 XH13/XA5/A 0 0.896691f
C117 XH13/XA6/A 0 1.098676f
C118 XH13/XA5/MN0/a_324_n18# 0 0.360407f
C119 XH13/XA4/MN0/a_324_n18# 0 0.360407f
C120 D<1> 0 0.918631f
C121 XH13/XA3/MN0/a_324_n18# 0 0.360407f
C122 XH13/XA6/C 0 1.328497f
C123 XH13/XA2/MN0/a_324_n18# 0 0.360407f
C124 XH13/XA1/MN0/a_324_n18# 0 0.360407f
C125 XH13/XA0/MN1/a_324_n18# 0 0.422415f
C126 XA4/MP1/G 0 0.884568f
C127 CKS 0 0.801993f
C128 CK_SAMPLE 0 0.805485f
C129 XA5/XA2/MN0/a_324_n18# 0 0.360407f
C130 XA5a/MN0/a_324_n18# 0 0.359492f
C131 XA5/XA2/A 0 0.888056f
C132 XA4/MN1/a_324_334# 0 0.359492f
C133 XA5/B 0 1.456308f
C134 XA6/A 0 1.690751f
C135 XA3/MN0/a_324_n18# 0 0.359492f
C136 XA4/MN0/a_324_n18# 0 0.359492f
C137 EN 0 0.153136f
C138 XA2/MP0/G 0 0.708335f
C139 TIE_L 0 0.1839f
C140 XA2/MN0/a_324_334# 0 0.422f
C141 XA1/MN1/a_324_n18# 0 0.422415f
C142 XC08/XA7/C 0 2.352415f
C143 XC08/QN 0 0.966414f
C144 DO<6> 0 0.963071f
C145 XC08/XA8/MN0/a_324_334# 0 0.422f
C146 XC08/XA8/MN0/a_324_n18# 0 0.360407f
C147 XC08/XA7/MN0/a_324_n18# 0 0.360407f
C148 XC08/XA6/MN0/a_324_n18# 0 0.360407f
C149 XC08/XA5/A 0 0.896691f
C150 XC08/XA6/A 0 1.098676f
C151 XC08/XA5/MN0/a_324_n18# 0 0.360407f
C152 XC08/XA4/MN0/a_324_n18# 0 0.360407f
C153 D<6> 0 0.918631f
C154 XC08/XA3/MN0/a_324_n18# 0 0.360407f
C155 XC08/XA6/C 0 1.328497f
C156 XC08/XA2/MN0/a_324_n18# 0 0.360407f
C157 XC08/XA1/MN0/a_324_n18# 0 0.360407f
C158 AVSS 0 -8.464535f
C159 XC08/XA0/MN1/a_324_n18# 0 0.422415f
C160 AVDD 0 0.152305p
C161 XE10/XA7/C 0 2.352415f
C162 XE10/QN 0 0.966414f
C163 DO<4> 0 0.963071f
C164 XE10/XA8/MN0/a_324_334# 0 0.422f
C165 XE10/XA8/MN0/a_324_n18# 0 0.360407f
C166 XE10/XA7/MN0/a_324_n18# 0 0.360407f
C167 XE10/XA6/MN0/a_324_n18# 0 0.360407f
C168 XE10/XA5/A 0 0.896691f
C169 XE10/XA6/A 0 1.098676f
C170 XE10/XA5/MN0/a_324_n18# 0 0.360407f
C171 XE10/XA4/MN0/a_324_n18# 0 0.360407f
C172 D<4> 0 0.918631f
C173 XE10/XA3/MN0/a_324_n18# 0 0.360407f
C174 XE10/XA6/C 0 1.328497f
C175 XE10/XA2/MN0/a_324_n18# 0 0.360407f
C176 XE10/XA1/MN0/a_324_n18# 0 0.360407f
C177 XE10/XA0/MN1/a_324_n18# 0 0.422415f
C178 XG12/XA7/C 0 2.352415f
C179 XG12/QN 0 0.966414f
C180 DO<2> 0 0.963071f
C181 XG12/XA8/MN0/a_324_334# 0 0.422f
C182 XG12/XA8/MN0/a_324_n18# 0 0.360407f
C183 XG12/XA7/MN0/a_324_n18# 0 0.360407f
C184 XG12/XA6/MN0/a_324_n18# 0 0.360407f
C185 XG12/XA5/A 0 0.896691f
C186 XG12/XA6/A 0 1.098676f
C187 XG12/XA5/MN0/a_324_n18# 0 0.360407f
C188 XG12/XA4/MN0/a_324_n18# 0 0.360407f
C189 D<2> 0 0.918631f
C190 XG12/XA3/MN0/a_324_n18# 0 0.360407f
C191 XG12/XA6/C 0 1.328497f
C192 XG12/XA2/MN0/a_324_n18# 0 0.360407f
C193 XG12/XA1/MN0/a_324_n18# 0 0.360407f
C194 XG12/XA0/MN1/a_324_n18# 0 0.422415f
C195 XI14/XA7/C 0 2.352415f
C196 XI14/QN 0 0.966414f
C197 DO<0> 0 0.960285f
C198 XI14/XA8/MN0/a_324_334# 0 0.422f
C199 XI14/XA8/MN0/a_324_n18# 0 0.360407f
C200 XI14/XA7/MN0/a_324_n18# 0 0.360407f
C201 XI14/XA6/MN0/a_324_n18# 0 0.360407f
C202 XI14/XA5/A 0 0.896691f
C203 XI14/XA6/A 0 1.098676f
C204 XI14/XA5/MN0/a_324_n18# 0 0.360407f
C205 XI14/XA4/MN0/a_324_n18# 0 0.360407f
C206 D<0> 0 1.011141f
C207 XI14/XA3/MN0/a_324_n18# 0 0.360407f
C208 XI14/XA6/C 0 1.328497f
C209 XI14/XA2/MN0/a_324_n18# 0 0.360407f
C210 XI14/XA1/MN0/a_324_n18# 0 0.360407f
C211 XI14/XA0/MN1/a_324_n18# 0 0.422415f
C212 ENABLE 0 0.918187f
C213 XA1/MN1/a_324_334# 0 0.359492f
C214 XB07/XA7/C 0 2.352415f
C215 XB07/QN 0 0.966414f
C216 DO<7> 0 0.973878f
C217 XB07/XA8/MN0/a_324_334# 0 0.422f
C218 XB07/XA8/MN0/a_324_n18# 0 0.360407f
C219 XB07/XA7/MN0/a_324_n18# 0 0.360407f
C220 XB07/XA6/MN0/a_324_n18# 0 0.360407f
C221 XB07/XA5/A 0 0.896691f
C222 XB07/XA6/A 0 1.098676f
C223 XB07/XA5/MN0/a_324_n18# 0 0.360407f
C224 XB07/XA4/MN0/a_324_n18# 0 0.360407f
C225 D<7> 0 1.10231f
C226 XB07/XA3/MN0/a_324_n18# 0 0.360407f
C227 XB07/XA6/C 0 1.328497f
C228 XB07/XA2/MN0/a_324_n18# 0 0.360407f
C229 DONE 0 9.575078f
C230 XB07/XA1/MN0/a_324_n18# 0 0.360407f
C231 XB07/XA0/MN1/a_324_n18# 0 0.422415f
C232 XD09/XA7/C 0 2.352415f
C233 XD09/QN 0 0.966414f
C234 DO<5> 0 0.965307f
C235 XD09/XA8/MN0/a_324_334# 0 0.422f
C236 XD09/XA8/MN0/a_324_n18# 0 0.360407f
C237 XD09/XA7/MN0/a_324_n18# 0 0.360407f
C238 XD09/XA6/MN0/a_324_n18# 0 0.360407f
C239 XD09/XA5/A 0 0.896691f
C240 XD09/XA6/A 0 1.098676f
C241 XD09/XA5/MN0/a_324_n18# 0 0.360407f
C242 XD09/XA4/MN0/a_324_n18# 0 0.360407f
C243 D<5> 0 0.918631f
C244 XD09/XA3/MN0/a_324_n18# 0 0.360407f
C245 XD09/XA6/C 0 1.328497f
C246 XD09/XA2/MN0/a_324_n18# 0 0.360407f
C247 XD09/XA1/MN0/a_324_n18# 0 0.360407f
C248 XD09/XA0/MN1/a_324_n18# 0 0.422415f
.ends

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
*+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
*+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
*+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
*+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
*+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
*+ VPWR VGND
Xtt_um_TT06_SAR_done_0 SUNSAR_SAR8B_CV_0/DONE uio_out[0] uio_oe[0] VPWR VGND tt_um_TT06_SAR_done
Xsky130_fd_pr__cap_mim_m3_1_XS736D_0 VPWR VGND VGND sky130_fd_pr__cap_mim_m3_1_XS736D
XSUNSAR_SAR8B_CV_0 ua[1] ua[0] SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/D<4>
+ SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0/XA6/CN0
+ SUNSAR_SAR8B_CV_0/XA6/CP0 SUNSAR_SAR8B_CV_0/XA3/CN0 SUNSAR_SAR8B_CV_0/XA3/CP0 SUNSAR_SAR8B_CV_0/CK_SAMPLE
+ SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/XA7/CP0 SUNSAR_SAR8B_CV_0/XA0/CEIN SUNSAR_SAR8B_CV_0/XA4/CN0
+ SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/CP0 SUNSAR_SAR8B_CV_0/XA1/CN0 SUNSAR_SAR8B_CV_0/D<6>
+ SUNSAR_SAR8B_CV_0/XA1/CP0 SUNSAR_SAR8B_CV_0/SARP SUNSAR_SAR8B_CV_0/XA5/CN0 SUNSAR_SAR8B_CV_0/D<2>
+ SUNSAR_SAR8B_CV_0/XA5/CP0 SUNSAR_SAR8B_CV_0/XA2/CN0 SUNSAR_SAR8B_CV_0/D<5> VPWR
+ SUNSAR_SAR8B_CV_0/XA2/CP0 SUNSAR_SAR8B_CV_0/SARN VPWR VGND SUNSAR_SAR8B_CV
XSUNSAR_CAPT8B_CV_0 clk ui_in[0] SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW
+ SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/D<5>
+ SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/D<1>
+ SUNSAR_SAR8B_CV_0/D<0> uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2]
+ uo_out[1] uo_out[0] TIE_L SUNSAR_SAR8B_CV_0/DONE VPWR VGND SUNSAR_CAPT8B_CV
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R1 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R2 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R3 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R4 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R5 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R6 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R7 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R8 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R9 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R10 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R11 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R12 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R13 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R14 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R15 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
C0 SUNSAR_SAR8B_CV_0/DONE ui_in[0] 0.159434f
C1 uio_oe[0] TIE_L1 0.902557f
C2 SUNSAR_SAR8B_CV_0/D<5> VGND 3.751857f
C3 SUNSAR_SAR8B_CV_0/D<5> VPWR 1.686887f
C4 TIE_L uo_out[4] 0.31941f
C5 TIE_L uo_out[7] 0.471918f
C6 VGND SUNSAR_SAR8B_CV_0/D<3> 3.719566f
C7 VGND SUNSAR_SAR8B_CV_0/D<2> 3.643656f
C8 VPWR SUNSAR_SAR8B_CV_0/D<3> 1.692954f
C9 VPWR SUNSAR_SAR8B_CV_0/D<2> 1.705346f
C10 SUNSAR_SAR8B_CV_0/XA0/CEIN VPWR 1.427229f
C11 SUNSAR_SAR8B_CV_0/XA0/CEIN ua[0] 0.982813f
C12 VGND SUNSAR_SAR8B_CV_0/XA6/CN0 -0.260744f
C13 TIE_L uo_out[3] 0.185334f
C14 SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/EN 0.131506f
C15 SUNSAR_SAR8B_CV_0/D<5> SUNSAR_SAR8B_CV_0/XA2/CP0 0.477434f
C16 SUNSAR_SAR8B_CV_0/EN ui_in[0] 0.968121f
C17 uo_out[7] uo_out[4] 0.121648f
C18 uo_out[1] uo_out[0] 0.328349f
C19 TIE_L VGND 0.100247f
C20 TIE_L VPWR 0.370965f
C21 clk TIE_L 0.13612f
C22 TIE_L uo_out[0] 0.278654f
C23 uio_oe[0] uo_out[5] 1.553295f
C24 uio_out[0] VGND 0.376081f
C25 SUNSAR_SAR8B_CV_0/XA7/CP0 SUNSAR_SAR8B_CV_0/D<0> 0.155245f
C26 uio_out[0] VPWR 0.145655f
C27 clk uio_out[0] 0.120689f
C28 uio_out[0] uo_out[0] 0.201579f
C29 SUNSAR_SAR8B_CV_0/D<6> VGND 3.637564f
C30 VGND SUNSAR_SAR8B_CV_0/XA4/CN0 -0.260744f
C31 SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/DONE 0.193713f
C32 SUNSAR_SAR8B_CV_0/D<6> VPWR 1.725454f
C33 uo_out[4] uo_out[3] 0.846609f
C34 VGND SUNSAR_SAR8B_CV_0/XA5/CN0 -0.26062f
C35 VPWR uo_out[7] 0.253367f
C36 uio_oe[0] uo_out[1] 0.432143f
C37 SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA1/CP0 0.476574f
C38 uio_oe[0] TIE_L 1.219126f
C39 SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA1/CN0 0.252238f
C40 VPWR uo_out[3] 0.234367f
C41 SUNSAR_SAR8B_CV_0/XA0/CEIN ua[1] 0.312742f
C42 SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/EN 0.315767f
C43 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW VGND 3.201681f
C44 VPWR SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0.187124f
C45 ua[0] SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0.437286f
C46 uio_oe[0] uio_out[0] 1.555271f
C47 TIE_L1 uo_out[5] 0.275794f
C48 uo_out[6] uo_out[5] 0.318994f
C49 TIE_L uo_out[2] 0.156661f
C50 ua[0] VGND 0.825069f
C51 VPWR VGND 24.256954f
C52 clk VGND 0.13736f
C53 ua[0] VPWR 0.537238f
C54 clk VPWR 0.185197f
C55 VGND SUNSAR_SAR8B_CV_0/XA3/CN0 -0.26062f
C56 SUNSAR_SAR8B_CV_0/CK_SAMPLE VGND 0.679252f
C57 uio_oe[0] uo_out[4] 0.550054f
C58 SUNSAR_SAR8B_CV_0/D<5> SUNSAR_SAR8B_CV_0/XA2/CN0 0.251493f
C59 SUNSAR_SAR8B_CV_0/CK_SAMPLE VPWR 2.139971f
C60 uio_oe[0] uo_out[7] 0.43252f
C61 SUNSAR_SAR8B_CV_0/XA0/XA4/A SUNSAR_SAR8B_CV_0/D<7> 0.103251f
C62 SUNSAR_SAR8B_CV_0/XA3/CP0 SUNSAR_SAR8B_CV_0/D<4> 0.151875f
C63 SUNSAR_SAR8B_CV_0/XA2/CP0 VGND -0.222661f
C64 SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/XA6/CP0 0.151117f
C65 SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/XA6/CN0 0.410141f
C66 SUNSAR_SAR8B_CV_0/XA1/CP0 VGND -0.221564f
C67 uio_oe[0] uo_out[3] 0.21235f
C68 SUNSAR_SAR8B_CV_0/XA1/CN0 VGND -0.15266f
C69 TIE_L TIE_L1 0.257793f
C70 TIE_L uo_out[6] 0.204625f
C71 uio_oe[0] VGND 0.340526f
C72 uio_oe[0] VPWR 1.039709f
C73 uio_oe[0] clk 0.260056f
C74 uio_oe[0] uo_out[0] 0.670799f
C75 SUNSAR_SAR8B_CV_0/DONE VGND 1.34648f
C76 ua[1] SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0.221633f
C77 TIE_L1 uo_out[7] 0.206895f
C78 VGND SUNSAR_SAR8B_CV_0/D<4> 3.598254f
C79 SUNSAR_SAR8B_CV_0/DONE VPWR 0.952355f
C80 uo_out[6] uo_out[4] 0.843602f
C81 VPWR SUNSAR_SAR8B_CV_0/D<4> 1.689756f
C82 uo_out[6] uo_out[7] 2.362091f
C83 ua[1] VGND 0.26469f
C84 ua[0] ua[1] 3.839995f
C85 ua[1] VPWR 0.257135f
C86 VGND ui_in[0] 0.483125f
C87 VPWR ui_in[0] 1.386636f
C88 clk ui_in[0] 0.134532f
C89 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA5/CP0 0.151875f
C90 SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/XA3/CN0 0.411522f
C91 TIE_L2 uo_out[7] 0.100011f
C92 TIE_L uo_out[5] 1.309194f
C93 uio_out[0] uo_out[5] 0.109219f
C94 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0/EN 0.127626f
C95 TIE_L1 VPWR 0.114647f
C96 uo_out[6] VGND 0.199834f
C97 uo_out[6] VPWR 0.323007f
C98 VGND SUNSAR_SAR8B_CV_0/D<1> 3.727024f
C99 VGND SUNSAR_SAR8B_CV_0/EN 0.490858f
C100 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/CP0 0.151117f
C101 VPWR SUNSAR_SAR8B_CV_0/D<1> 1.714778f
C102 VPWR SUNSAR_SAR8B_CV_0/EN 7.947423f
C103 uio_oe[0] uo_out[2] 0.267753f
C104 SUNSAR_SAR8B_CV_0/XA2/CN0 VGND -0.152784f
C105 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/CN0 0.410141f
C106 uo_out[5] uo_out[4] 1.133807f
C107 uo_out[5] uo_out[7] 1.578182f
C108 VGND SUNSAR_SAR8B_CV_0/D<7> 1.927649f
C109 VPWR SUNSAR_SAR8B_CV_0/D<7> 0.570534f
C110 TIE_L uo_out[1] 0.50141f
C111 SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/XA7/CEO 0.123345f
C112 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/EN 0.494615f
C113 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA5/CN0 0.411523f
C114 SUNSAR_SAR8B_CV_0/D<0> VGND 3.041315f
C115 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<7> 0.174845f
C116 SUNSAR_SAR8B_CV_0/D<0> VPWR 1.952988f
C117 uio_out[0] TIE_L 0.44106f
C118 ua[2] 0 0.119794f
C119 ua[3] 0 0.119794f
C120 ua[4] 0 0.121038f
C121 ua[5] 0 0.122428f
C122 ua[6] 0 0.122428f
C123 ua[7] 0 0.111009f
C124 TIE_L1 0 1.51307f
C125 TIE_L2 0 1.83212f
C126 m1_14848_7490# 0 0.145721f $ **FLOATING
C127 SUNSAR_CAPT8B_CV_0/XF11/XA7/C 0 2.352415f
C128 SUNSAR_CAPT8B_CV_0/XF11/QN 0 0.966414f
C129 uo_out[3] 0 1.33751f
C130 SUNSAR_CAPT8B_CV_0/XF11/XA8/MN0/a_324_334# 0 0.422f
C131 SUNSAR_CAPT8B_CV_0/XF11/XA8/MN0/a_324_n18# 0 0.360407f
C132 SUNSAR_CAPT8B_CV_0/XF11/XA7/MN0/a_324_n18# 0 0.360407f
C133 SUNSAR_CAPT8B_CV_0/XF11/XA6/MN0/a_324_n18# 0 0.360407f
C134 SUNSAR_CAPT8B_CV_0/XF11/XA5/A 0 0.896691f
C135 SUNSAR_CAPT8B_CV_0/XF11/XA6/A 0 1.098676f
C136 SUNSAR_CAPT8B_CV_0/XF11/XA5/MN0/a_324_n18# 0 0.360407f
C137 SUNSAR_CAPT8B_CV_0/XF11/XA4/MN0/a_324_n18# 0 0.360407f
C138 SUNSAR_CAPT8B_CV_0/XF11/XA3/MN0/a_324_n18# 0 0.360407f
C139 SUNSAR_CAPT8B_CV_0/XF11/XA6/C 0 1.328497f
C140 SUNSAR_CAPT8B_CV_0/XF11/XA2/MN0/a_324_n18# 0 0.360407f
C141 SUNSAR_CAPT8B_CV_0/XF11/XA1/MN0/a_324_n18# 0 0.360407f
C142 SUNSAR_CAPT8B_CV_0/XF11/XA0/MN1/a_324_n18# 0 0.422415f
C143 SUNSAR_CAPT8B_CV_0/XA6/XA2/MN0/a_324_n18# 0 0.360407f
C144 SUNSAR_CAPT8B_CV_0/XA2/MN0/a_324_n18# 0 0.359492f
C145 SUNSAR_CAPT8B_CV_0/XA5a/MN0/a_324_334# 0 0.359492f
C146 SUNSAR_CAPT8B_CV_0/XA6/XA2/A 0 0.871363f
C147 SUNSAR_CAPT8B_CV_0/XA6/B 0 1.026139f
C148 SUNSAR_CAPT8B_CV_0/XH13/XA7/C 0 2.352415f
C149 SUNSAR_CAPT8B_CV_0/XH13/QN 0 0.966414f
C150 uo_out[1] 0 1.194172f
C151 SUNSAR_CAPT8B_CV_0/XH13/XA8/MN0/a_324_334# 0 0.422f
C152 SUNSAR_CAPT8B_CV_0/XH13/XA8/MN0/a_324_n18# 0 0.360407f
C153 SUNSAR_CAPT8B_CV_0/XH13/XA7/MN0/a_324_n18# 0 0.360407f
C154 SUNSAR_CAPT8B_CV_0/XH13/XA6/MN0/a_324_n18# 0 0.360407f
C155 SUNSAR_CAPT8B_CV_0/XH13/XA5/A 0 0.896691f
C156 SUNSAR_CAPT8B_CV_0/XH13/XA6/A 0 1.098676f
C157 SUNSAR_CAPT8B_CV_0/XH13/XA5/MN0/a_324_n18# 0 0.360407f
C158 SUNSAR_CAPT8B_CV_0/XH13/XA4/MN0/a_324_n18# 0 0.360407f
C159 SUNSAR_CAPT8B_CV_0/XH13/XA3/MN0/a_324_n18# 0 0.360407f
C160 SUNSAR_CAPT8B_CV_0/XH13/XA6/C 0 1.328497f
C161 SUNSAR_CAPT8B_CV_0/XH13/XA2/MN0/a_324_n18# 0 0.360407f
C162 SUNSAR_CAPT8B_CV_0/XH13/XA1/MN0/a_324_n18# 0 0.360407f
C163 SUNSAR_CAPT8B_CV_0/XH13/XA0/MN1/a_324_n18# 0 0.422415f
C164 SUNSAR_CAPT8B_CV_0/XA4/MP1/G 0 0.884568f
C165 clk 0 2.385743f
C166 SUNSAR_CAPT8B_CV_0/XA5/XA2/MN0/a_324_n18# 0 0.360407f
C167 SUNSAR_CAPT8B_CV_0/XA5a/MN0/a_324_n18# 0 0.359492f
C168 SUNSAR_CAPT8B_CV_0/XA5/XA2/A 0 0.888056f
C169 SUNSAR_CAPT8B_CV_0/XA4/MN1/a_324_334# 0 0.359492f
C170 SUNSAR_CAPT8B_CV_0/XA5/B 0 1.456308f
C171 SUNSAR_CAPT8B_CV_0/XA6/A 0 1.690751f
C172 SUNSAR_CAPT8B_CV_0/XA3/MN0/a_324_n18# 0 0.359492f
C173 SUNSAR_CAPT8B_CV_0/XA4/MN0/a_324_n18# 0 0.359492f
C174 SUNSAR_CAPT8B_CV_0/XA2/MP0/G 0 0.708335f
C175 TIE_L 0 0.99989f
C176 SUNSAR_CAPT8B_CV_0/XA2/MN0/a_324_334# 0 0.422f
C177 SUNSAR_CAPT8B_CV_0/XA1/MN1/a_324_n18# 0 0.422415f
C178 SUNSAR_CAPT8B_CV_0/XC08/XA7/C 0 2.352415f
C179 SUNSAR_CAPT8B_CV_0/XC08/QN 0 0.966414f
C180 uo_out[6] 0 1.372751f
C181 SUNSAR_CAPT8B_CV_0/XC08/XA8/MN0/a_324_334# 0 0.422f
C182 SUNSAR_CAPT8B_CV_0/XC08/XA8/MN0/a_324_n18# 0 0.360407f
C183 SUNSAR_CAPT8B_CV_0/XC08/XA7/MN0/a_324_n18# 0 0.360407f
C184 SUNSAR_CAPT8B_CV_0/XC08/XA6/MN0/a_324_n18# 0 0.360407f
C185 SUNSAR_CAPT8B_CV_0/XC08/XA5/A 0 0.896691f
C186 SUNSAR_CAPT8B_CV_0/XC08/XA6/A 0 1.098676f
C187 SUNSAR_CAPT8B_CV_0/XC08/XA5/MN0/a_324_n18# 0 0.360407f
C188 SUNSAR_CAPT8B_CV_0/XC08/XA4/MN0/a_324_n18# 0 0.360407f
C189 SUNSAR_CAPT8B_CV_0/XC08/XA3/MN0/a_324_n18# 0 0.360407f
C190 SUNSAR_CAPT8B_CV_0/XC08/XA6/C 0 1.328497f
C191 SUNSAR_CAPT8B_CV_0/XC08/XA2/MN0/a_324_n18# 0 0.360407f
C192 SUNSAR_CAPT8B_CV_0/XC08/XA1/MN0/a_324_n18# 0 0.360407f
C193 SUNSAR_CAPT8B_CV_0/XC08/XA0/MN1/a_324_n18# 0 0.422415f
C194 SUNSAR_CAPT8B_CV_0/XE10/XA7/C 0 2.352415f
C195 SUNSAR_CAPT8B_CV_0/XE10/QN 0 0.966414f
C196 uo_out[4] 0 1.095506f
C197 SUNSAR_CAPT8B_CV_0/XE10/XA8/MN0/a_324_334# 0 0.422f
C198 SUNSAR_CAPT8B_CV_0/XE10/XA8/MN0/a_324_n18# 0 0.360407f
C199 SUNSAR_CAPT8B_CV_0/XE10/XA7/MN0/a_324_n18# 0 0.360407f
C200 SUNSAR_CAPT8B_CV_0/XE10/XA6/MN0/a_324_n18# 0 0.360407f
C201 SUNSAR_CAPT8B_CV_0/XE10/XA5/A 0 0.896691f
C202 SUNSAR_CAPT8B_CV_0/XE10/XA6/A 0 1.098676f
C203 SUNSAR_CAPT8B_CV_0/XE10/XA5/MN0/a_324_n18# 0 0.360407f
C204 SUNSAR_CAPT8B_CV_0/XE10/XA4/MN0/a_324_n18# 0 0.360407f
C205 SUNSAR_CAPT8B_CV_0/XE10/XA3/MN0/a_324_n18# 0 0.360407f
C206 SUNSAR_CAPT8B_CV_0/XE10/XA6/C 0 1.328497f
C207 SUNSAR_CAPT8B_CV_0/XE10/XA2/MN0/a_324_n18# 0 0.360407f
C208 SUNSAR_CAPT8B_CV_0/XE10/XA1/MN0/a_324_n18# 0 0.360407f
C209 SUNSAR_CAPT8B_CV_0/XE10/XA0/MN1/a_324_n18# 0 0.422415f
C210 SUNSAR_CAPT8B_CV_0/XG12/XA7/C 0 2.352415f
C211 SUNSAR_CAPT8B_CV_0/XG12/QN 0 0.966414f
C212 uo_out[2] 0 1.120428f
C213 SUNSAR_CAPT8B_CV_0/XG12/XA8/MN0/a_324_334# 0 0.422f
C214 SUNSAR_CAPT8B_CV_0/XG12/XA8/MN0/a_324_n18# 0 0.360407f
C215 SUNSAR_CAPT8B_CV_0/XG12/XA7/MN0/a_324_n18# 0 0.360407f
C216 SUNSAR_CAPT8B_CV_0/XG12/XA6/MN0/a_324_n18# 0 0.360407f
C217 SUNSAR_CAPT8B_CV_0/XG12/XA5/A 0 0.896691f
C218 SUNSAR_CAPT8B_CV_0/XG12/XA6/A 0 1.098676f
C219 SUNSAR_CAPT8B_CV_0/XG12/XA5/MN0/a_324_n18# 0 0.360407f
C220 SUNSAR_CAPT8B_CV_0/XG12/XA4/MN0/a_324_n18# 0 0.360407f
C221 SUNSAR_CAPT8B_CV_0/XG12/XA3/MN0/a_324_n18# 0 0.360407f
C222 SUNSAR_CAPT8B_CV_0/XG12/XA6/C 0 1.328497f
C223 SUNSAR_CAPT8B_CV_0/XG12/XA2/MN0/a_324_n18# 0 0.360407f
C224 SUNSAR_CAPT8B_CV_0/XG12/XA1/MN0/a_324_n18# 0 0.360407f
C225 SUNSAR_CAPT8B_CV_0/XG12/XA0/MN1/a_324_n18# 0 0.422415f
C226 SUNSAR_CAPT8B_CV_0/XI14/XA7/C 0 2.352415f
C227 SUNSAR_CAPT8B_CV_0/XI14/QN 0 0.966414f
C228 uo_out[0] 0 1.493281f
C229 SUNSAR_CAPT8B_CV_0/XI14/XA8/MN0/a_324_334# 0 0.422f
C230 SUNSAR_CAPT8B_CV_0/XI14/XA8/MN0/a_324_n18# 0 0.360407f
C231 SUNSAR_CAPT8B_CV_0/XI14/XA7/MN0/a_324_n18# 0 0.360407f
C232 SUNSAR_CAPT8B_CV_0/XI14/XA6/MN0/a_324_n18# 0 0.360407f
C233 SUNSAR_CAPT8B_CV_0/XI14/XA5/A 0 0.896691f
C234 SUNSAR_CAPT8B_CV_0/XI14/XA6/A 0 1.098676f
C235 SUNSAR_CAPT8B_CV_0/XI14/XA5/MN0/a_324_n18# 0 0.360407f
C236 SUNSAR_CAPT8B_CV_0/XI14/XA4/MN0/a_324_n18# 0 0.360407f
C237 SUNSAR_CAPT8B_CV_0/XI14/XA3/MN0/a_324_n18# 0 0.360407f
C238 SUNSAR_CAPT8B_CV_0/XI14/XA6/C 0 1.328497f
C239 SUNSAR_CAPT8B_CV_0/XI14/XA2/MN0/a_324_n18# 0 0.360407f
C240 SUNSAR_CAPT8B_CV_0/XI14/XA1/MN0/a_324_n18# 0 0.360407f
C241 SUNSAR_CAPT8B_CV_0/XI14/XA0/MN1/a_324_n18# 0 0.422415f
C242 ui_in[0] 0 1.237376f
C243 SUNSAR_CAPT8B_CV_0/XA1/MN1/a_324_334# 0 0.359492f
C244 SUNSAR_CAPT8B_CV_0/XB07/XA7/C 0 2.352415f
C245 SUNSAR_CAPT8B_CV_0/XB07/QN 0 0.966414f
C246 uo_out[7] 0 1.986758f
C247 SUNSAR_CAPT8B_CV_0/XB07/XA8/MN0/a_324_334# 0 0.422f
C248 SUNSAR_CAPT8B_CV_0/XB07/XA8/MN0/a_324_n18# 0 0.360407f
C249 SUNSAR_CAPT8B_CV_0/XB07/XA7/MN0/a_324_n18# 0 0.360407f
C250 SUNSAR_CAPT8B_CV_0/XB07/XA6/MN0/a_324_n18# 0 0.360407f
C251 SUNSAR_CAPT8B_CV_0/XB07/XA5/A 0 0.896691f
C252 SUNSAR_CAPT8B_CV_0/XB07/XA6/A 0 1.098676f
C253 SUNSAR_CAPT8B_CV_0/XB07/XA5/MN0/a_324_n18# 0 0.360407f
C254 SUNSAR_CAPT8B_CV_0/XB07/XA4/MN0/a_324_n18# 0 0.360407f
C255 SUNSAR_CAPT8B_CV_0/XB07/XA3/MN0/a_324_n18# 0 0.360407f
C256 SUNSAR_CAPT8B_CV_0/XB07/XA6/C 0 1.328497f
C257 SUNSAR_CAPT8B_CV_0/XB07/XA2/MN0/a_324_n18# 0 0.360407f
C258 SUNSAR_SAR8B_CV_0/DONE 0 12.867176f
C259 SUNSAR_CAPT8B_CV_0/XB07/XA1/MN0/a_324_n18# 0 0.360407f
C260 SUNSAR_CAPT8B_CV_0/XB07/XA0/MN1/a_324_n18# 0 0.422415f
C261 SUNSAR_CAPT8B_CV_0/XD09/XA7/C 0 2.352415f
C262 SUNSAR_CAPT8B_CV_0/XD09/QN 0 0.966414f
C263 uo_out[5] 0 1.119996f
C264 SUNSAR_CAPT8B_CV_0/XD09/XA8/MN0/a_324_334# 0 0.422f
C265 SUNSAR_CAPT8B_CV_0/XD09/XA8/MN0/a_324_n18# 0 0.360407f
C266 SUNSAR_CAPT8B_CV_0/XD09/XA7/MN0/a_324_n18# 0 0.360407f
C267 SUNSAR_CAPT8B_CV_0/XD09/XA6/MN0/a_324_n18# 0 0.360407f
C268 SUNSAR_CAPT8B_CV_0/XD09/XA5/A 0 0.896691f
C269 SUNSAR_CAPT8B_CV_0/XD09/XA6/A 0 1.098676f
C270 SUNSAR_CAPT8B_CV_0/XD09/XA5/MN0/a_324_n18# 0 0.360407f
C271 SUNSAR_CAPT8B_CV_0/XD09/XA4/MN0/a_324_n18# 0 0.360407f
C272 SUNSAR_CAPT8B_CV_0/XD09/XA3/MN0/a_324_n18# 0 0.360407f
C273 SUNSAR_CAPT8B_CV_0/XD09/XA6/C 0 1.328497f
C274 SUNSAR_CAPT8B_CV_0/XD09/XA2/MN0/a_324_n18# 0 0.360407f
C275 SUNSAR_CAPT8B_CV_0/XD09/XA1/MN0/a_324_n18# 0 0.360407f
C276 SUNSAR_CAPT8B_CV_0/XD09/XA0/MN1/a_324_n18# 0 0.422415f
C277 SUNSAR_SAR8B_CV_0/XA7/XA9/MN1/a_324_334# 0 0.360407f
C278 SUNSAR_SAR8B_CV_0/XA7/XA9/MN0/a_324_n18# 0 0.360407f
C279 SUNSAR_SAR8B_CV_0/XA7/XA9/A 0 1.250075f
C280 SUNSAR_SAR8B_CV_0/XA7/XA7/MN0/a_324_n18# 0 0.360407f
C281 SUNSAR_SAR8B_CV_0/XA7/XA8/MN0/a_324_n18# 0 0.360407f
C282 SUNSAR_SAR8B_CV_0/XA7/XA9/B 0 1.158058f
C283 SUNSAR_SAR8B_CV_0/XA7/XA6/MN0/a_324_n18# 0 0.360407f
C284 SUNSAR_SAR8B_CV_0/XA7/XA4/A 0 2.621765f
C285 SUNSAR_SAR8B_CV_0/XA7/XA4/MN0/a_324_n18# 0 0.360407f
C286 SUNSAR_SAR8B_CV_0/XA7/CP0 0 2.4163f
C287 SUNSAR_SAR8B_CV_0/XA7/CN0 0 0.312365f
C288 SUNSAR_SAR8B_CV_0/XA7/XA5/MN0/a_324_n18# 0 0.360407f
C289 SUNSAR_SAR8B_CV_0/XA7/CN1 0 2.428168f
C290 SUNSAR_SAR8B_CV_0/D<0> 0 1.87393f
C291 SUNSAR_SAR8B_CV_0/XA7/XA3/MN0/a_324_n18# 0 0.360407f
C292 SUNSAR_SAR8B_CV_0/XA7/XA2/A 0 2.030764f
C293 SUNSAR_SAR8B_CV_0/XA7/XA2/MN0/a_324_n18# 0 0.360407f
C294 SUNSAR_SAR8B_CV_0/XA7/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C295 SUNSAR_SAR8B_CV_0/XA7/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C296 SUNSAR_SAR8B_CV_0/XA7/XA1/XA2/Y 0 1.060197f
C297 SUNSAR_SAR8B_CV_0/XA7/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C298 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C299 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C300 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C301 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MP3/G 0 0.827484f
C302 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN2/S 0 0.200627f
C303 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C304 SUNSAR_SAR8B_CV_0/XA7/ENO 0 1.582724f
C305 SUNSAR_SAR8B_CV_0/XA7/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C306 SUNSAR_SAR8B_CV_0/XA7/XA13/MN1/a_324_334# 0 0.422f
C307 SUNSAR_SAR8B_CV_0/XA7/XA12/MN0/a_324_n18# 0 0.360407f
C308 SUNSAR_SAR8B_CV_0/XA7/XA13/MN1/a_324_n18# 0 0.360407f
C309 SUNSAR_SAR8B_CV_0/XA7/XA12/A 0 0.755669f
C310 SUNSAR_SAR8B_CV_0/XA7/XA11/MN0/a_324_n18# 0 0.360407f
C311 SUNSAR_SAR8B_CV_0/XA6/CEO 0 1.009021f
C312 SUNSAR_SAR8B_CV_0/XA7/XA11/A 0 0.662715f
C313 SUNSAR_SAR8B_CV_0/XA7/XA9/Y 0 0.718246f
C314 SUNSAR_SAR8B_CV_0/XA6/XA9/MN1/a_324_334# 0 0.360407f
C315 SUNSAR_SAR8B_CV_0/XA6/XA9/MN0/a_324_n18# 0 0.360407f
C316 SUNSAR_SAR8B_CV_0/XA6/XA9/A 0 1.250075f
C317 SUNSAR_SAR8B_CV_0/XA6/DONE 0 0.13094f
C318 SUNSAR_SAR8B_CV_0/XA6/XA7/MN0/a_324_n18# 0 0.360407f
C319 SUNSAR_SAR8B_CV_0/XA6/XA8/MN0/a_324_n18# 0 0.360407f
C320 SUNSAR_SAR8B_CV_0/XA6/XA9/B 0 1.158058f
C321 SUNSAR_SAR8B_CV_0/XA6/XA6/MN0/a_324_n18# 0 0.360407f
C322 SUNSAR_SAR8B_CV_0/XA6/XA4/A 0 2.621765f
C323 SUNSAR_SAR8B_CV_0/XA6/XA4/MN0/a_324_n18# 0 0.360407f
C324 SUNSAR_SAR8B_CV_0/XA6/CP0 0 2.4163f
C325 SUNSAR_SAR8B_CV_0/XA6/CN0 0 4.160099f
C326 SUNSAR_SAR8B_CV_0/XA6/XA5/MN0/a_324_n18# 0 0.360407f
C327 SUNSAR_SAR8B_CV_0/XA6/CN1 0 2.428168f
C328 SUNSAR_SAR8B_CV_0/D<1> 0 5.818007f
C329 SUNSAR_SAR8B_CV_0/XA6/XA3/MN0/a_324_n18# 0 0.360407f
C330 SUNSAR_SAR8B_CV_0/XA6/XA2/A 0 2.030764f
C331 SUNSAR_SAR8B_CV_0/XA6/XA2/MN0/a_324_n18# 0 0.360407f
C332 SUNSAR_SAR8B_CV_0/XA6/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C333 SUNSAR_SAR8B_CV_0/XA6/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C334 SUNSAR_SAR8B_CV_0/XA6/XA1/XA2/Y 0 1.060197f
C335 SUNSAR_SAR8B_CV_0/XA6/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C336 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C337 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C338 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C339 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MP3/G 0 0.827484f
C340 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN2/S 0 0.200627f
C341 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C342 SUNSAR_SAR8B_CV_0/XA7/EN 0 3.856368f
C343 SUNSAR_SAR8B_CV_0/XA6/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C344 SUNSAR_SAR8B_CV_0/XA6/XA13/MN1/a_324_334# 0 0.422f
C345 SUNSAR_SAR8B_CV_0/XA6/XA12/MN0/a_324_n18# 0 0.360407f
C346 SUNSAR_SAR8B_CV_0/XA6/XA13/MN1/a_324_n18# 0 0.360407f
C347 SUNSAR_SAR8B_CV_0/XA6/XA12/A 0 0.755669f
C348 SUNSAR_SAR8B_CV_0/XA6/XA11/MN0/a_324_n18# 0 0.360407f
C349 SUNSAR_SAR8B_CV_0/XA5/CEO 0 1.104751f
C350 SUNSAR_SAR8B_CV_0/XA6/XA11/A 0 0.662715f
C351 SUNSAR_SAR8B_CV_0/XA6/XA9/Y 0 0.718246f
C352 SUNSAR_SAR8B_CV_0/XA5/XA9/MN1/a_324_334# 0 0.360407f
C353 SUNSAR_SAR8B_CV_0/XA5/XA9/MN0/a_324_n18# 0 0.360407f
C354 SUNSAR_SAR8B_CV_0/XA5/XA9/A 0 1.250075f
C355 SUNSAR_SAR8B_CV_0/XA5/DONE 0 0.123486f
C356 SUNSAR_SAR8B_CV_0/XA5/XA7/MN0/a_324_n18# 0 0.360407f
C357 SUNSAR_SAR8B_CV_0/XA5/XA8/MN0/a_324_n18# 0 0.360407f
C358 SUNSAR_SAR8B_CV_0/XA5/XA9/B 0 1.158058f
C359 SUNSAR_SAR8B_CV_0/XA5/XA6/MN0/a_324_n18# 0 0.360407f
C360 SUNSAR_SAR8B_CV_0/XA5/XA4/A 0 2.621765f
C361 SUNSAR_SAR8B_CV_0/XA5/XA4/MN0/a_324_n18# 0 0.360407f
C362 SUNSAR_SAR8B_CV_0/XA5/CP0 0 2.4163f
C363 SUNSAR_SAR8B_CV_0/XA5/CN0 0 3.052303f
C364 SUNSAR_SAR8B_CV_0/XA5/XA5/MN0/a_324_n18# 0 0.360407f
C365 SUNSAR_SAR8B_CV_0/XA5/CN1 0 2.428168f
C366 SUNSAR_SAR8B_CV_0/D<2> 0 5.190204f
C367 SUNSAR_SAR8B_CV_0/XA5/XA3/MN0/a_324_n18# 0 0.360407f
C368 SUNSAR_SAR8B_CV_0/XA5/XA2/A 0 2.030764f
C369 SUNSAR_SAR8B_CV_0/XA5/XA2/MN0/a_324_n18# 0 0.360407f
C370 SUNSAR_SAR8B_CV_0/XA5/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C371 SUNSAR_SAR8B_CV_0/XA5/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C372 SUNSAR_SAR8B_CV_0/XA5/XA1/XA2/Y 0 1.060197f
C373 SUNSAR_SAR8B_CV_0/XA5/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C374 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C375 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C376 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C377 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MP3/G 0 0.827484f
C378 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN2/S 0 0.200627f
C379 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C380 SUNSAR_SAR8B_CV_0/XA6/EN 0 3.679756f
C381 SUNSAR_SAR8B_CV_0/XA5/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C382 SUNSAR_SAR8B_CV_0/XA5/XA13/MN1/a_324_334# 0 0.422f
C383 SUNSAR_SAR8B_CV_0/XA5/XA12/MN0/a_324_n18# 0 0.360407f
C384 SUNSAR_SAR8B_CV_0/XA5/XA13/MN1/a_324_n18# 0 0.360407f
C385 SUNSAR_SAR8B_CV_0/XA5/XA12/A 0 0.755669f
C386 SUNSAR_SAR8B_CV_0/XA5/XA11/MN0/a_324_n18# 0 0.360407f
C387 SUNSAR_SAR8B_CV_0/XA4/CEO 0 1.086041f
C388 SUNSAR_SAR8B_CV_0/XA5/XA11/A 0 0.662715f
C389 SUNSAR_SAR8B_CV_0/XA5/XA9/Y 0 0.718246f
C390 SUNSAR_SAR8B_CV_0/XA4/XA9/MN1/a_324_334# 0 0.360407f
C391 SUNSAR_SAR8B_CV_0/XA4/XA9/MN0/a_324_n18# 0 0.360407f
C392 SUNSAR_SAR8B_CV_0/XA4/XA9/A 0 1.250075f
C393 SUNSAR_SAR8B_CV_0/XA4/DONE 0 0.13094f
C394 SUNSAR_SAR8B_CV_0/XA4/XA7/MN0/a_324_n18# 0 0.360407f
C395 SUNSAR_SAR8B_CV_0/XA4/XA8/MN0/a_324_n18# 0 0.360407f
C396 SUNSAR_SAR8B_CV_0/XA4/XA9/B 0 1.158058f
C397 SUNSAR_SAR8B_CV_0/XA4/XA6/MN0/a_324_n18# 0 0.360407f
C398 SUNSAR_SAR8B_CV_0/XA4/XA4/A 0 2.621765f
C399 SUNSAR_SAR8B_CV_0/XA4/XA4/MN0/a_324_n18# 0 0.360407f
C400 SUNSAR_SAR8B_CV_0/XA4/CP0 0 2.4163f
C401 SUNSAR_SAR8B_CV_0/XA4/CN0 0 2.237548f
C402 SUNSAR_SAR8B_CV_0/XA4/XA5/MN0/a_324_n18# 0 0.360407f
C403 SUNSAR_SAR8B_CV_0/XA4/CN1 0 2.428168f
C404 SUNSAR_SAR8B_CV_0/D<3> 0 4.013408f
C405 SUNSAR_SAR8B_CV_0/XA4/XA3/MN0/a_324_n18# 0 0.360407f
C406 SUNSAR_SAR8B_CV_0/XA4/XA2/A 0 2.030764f
C407 SUNSAR_SAR8B_CV_0/XA4/XA2/MN0/a_324_n18# 0 0.360407f
C408 SUNSAR_SAR8B_CV_0/XA4/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C409 SUNSAR_SAR8B_CV_0/XA4/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C410 SUNSAR_SAR8B_CV_0/XA4/XA1/XA2/Y 0 1.060197f
C411 SUNSAR_SAR8B_CV_0/XA4/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C412 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C413 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C414 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C415 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MP3/G 0 0.827484f
C416 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN2/S 0 0.200627f
C417 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C418 SUNSAR_SAR8B_CV_0/XA5/EN 0 3.635208f
C419 SUNSAR_SAR8B_CV_0/XA4/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C420 SUNSAR_SAR8B_CV_0/XA4/XA13/MN1/a_324_334# 0 0.422f
C421 SUNSAR_SAR8B_CV_0/XA4/XA12/MN0/a_324_n18# 0 0.360407f
C422 SUNSAR_SAR8B_CV_0/XA4/XA13/MN1/a_324_n18# 0 0.360407f
C423 SUNSAR_SAR8B_CV_0/XA4/XA12/A 0 0.755669f
C424 SUNSAR_SAR8B_CV_0/XA4/XA11/MN0/a_324_n18# 0 0.360407f
C425 SUNSAR_SAR8B_CV_0/XA3/CEO 0 1.107611f
C426 SUNSAR_SAR8B_CV_0/XA4/XA11/A 0 0.662715f
C427 SUNSAR_SAR8B_CV_0/XA4/XA9/Y 0 0.718246f
C428 SUNSAR_SAR8B_CV_0/XA3/XA9/MN1/a_324_334# 0 0.360407f
C429 SUNSAR_SAR8B_CV_0/XA3/XA9/MN0/a_324_n18# 0 0.360407f
C430 SUNSAR_SAR8B_CV_0/XA3/XA9/A 0 1.250075f
C431 SUNSAR_SAR8B_CV_0/XA3/DONE 0 0.123486f
C432 SUNSAR_SAR8B_CV_0/XA3/XA7/MN0/a_324_n18# 0 0.360407f
C433 SUNSAR_SAR8B_CV_0/XA3/XA8/MN0/a_324_n18# 0 0.360407f
C434 SUNSAR_SAR8B_CV_0/XA3/XA9/B 0 1.158058f
C435 SUNSAR_SAR8B_CV_0/XA3/XA6/MN0/a_324_n18# 0 0.360407f
C436 SUNSAR_SAR8B_CV_0/XA3/XA4/A 0 2.621765f
C437 SUNSAR_SAR8B_CV_0/XA3/XA4/MN0/a_324_n18# 0 0.360407f
C438 SUNSAR_SAR8B_CV_0/XA3/CP0 0 2.4163f
C439 SUNSAR_SAR8B_CV_0/XA3/CN0 0 3.224855f
C440 SUNSAR_SAR8B_CV_0/XA3/XA5/MN0/a_324_n18# 0 0.360407f
C441 SUNSAR_SAR8B_CV_0/XA3/CN1 0 2.428168f
C442 SUNSAR_SAR8B_CV_0/D<4> 0 4.549352f
C443 SUNSAR_SAR8B_CV_0/XA3/XA3/MN0/a_324_n18# 0 0.360407f
C444 SUNSAR_SAR8B_CV_0/XA3/XA2/A 0 2.030764f
C445 SUNSAR_SAR8B_CV_0/XA3/XA2/MN0/a_324_n18# 0 0.360407f
C446 SUNSAR_SAR8B_CV_0/XA3/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C447 SUNSAR_SAR8B_CV_0/XA3/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C448 SUNSAR_SAR8B_CV_0/XA3/XA1/XA2/Y 0 1.060197f
C449 SUNSAR_SAR8B_CV_0/XA3/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C450 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C451 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C452 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C453 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MP3/G 0 0.827484f
C454 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN2/S 0 0.200627f
C455 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C456 SUNSAR_SAR8B_CV_0/XA4/EN 0 3.720665f
C457 SUNSAR_SAR8B_CV_0/XA3/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C458 SUNSAR_SAR8B_CV_0/XA3/XA13/MN1/a_324_334# 0 0.422f
C459 SUNSAR_SAR8B_CV_0/XA3/XA12/MN0/a_324_n18# 0 0.360407f
C460 SUNSAR_SAR8B_CV_0/XA3/XA13/MN1/a_324_n18# 0 0.360407f
C461 SUNSAR_SAR8B_CV_0/XA3/XA12/A 0 0.755669f
C462 SUNSAR_SAR8B_CV_0/XA3/XA11/MN0/a_324_n18# 0 0.360407f
C463 SUNSAR_SAR8B_CV_0/XA2/CEO 0 1.085281f
C464 SUNSAR_SAR8B_CV_0/XA3/XA11/A 0 0.662715f
C465 SUNSAR_SAR8B_CV_0/XA3/XA9/Y 0 0.718246f
C466 SUNSAR_SAR8B_CV_0/XA2/XA9/MN1/a_324_334# 0 0.360407f
C467 SUNSAR_SAR8B_CV_0/XA2/XA9/MN0/a_324_n18# 0 0.360407f
C468 SUNSAR_SAR8B_CV_0/XA2/XA9/A 0 1.250075f
C469 SUNSAR_SAR8B_CV_0/XA2/DONE 0 0.13094f
C470 SUNSAR_SAR8B_CV_0/XA2/XA7/MN0/a_324_n18# 0 0.360407f
C471 SUNSAR_SAR8B_CV_0/XA2/XA8/MN0/a_324_n18# 0 0.360407f
C472 SUNSAR_SAR8B_CV_0/XA2/XA9/B 0 1.158058f
C473 SUNSAR_SAR8B_CV_0/XA2/XA6/MN0/a_324_n18# 0 0.360407f
C474 SUNSAR_SAR8B_CV_0/XA2/XA4/A 0 2.621765f
C475 SUNSAR_SAR8B_CV_0/XA2/XA4/MN0/a_324_n18# 0 0.360407f
C476 SUNSAR_SAR8B_CV_0/XA2/CP0 0 4.49437f
C477 SUNSAR_SAR8B_CV_0/XA2/CN0 0 2.820252f
C478 SUNSAR_SAR8B_CV_0/XA2/XA5/MN0/a_324_n18# 0 0.360407f
C479 SUNSAR_SAR8B_CV_0/XA2/CN1 0 6.112935f
C480 SUNSAR_SAR8B_CV_0/XA2/XA3/MN0/a_324_n18# 0 0.360407f
C481 SUNSAR_SAR8B_CV_0/XA2/XA2/A 0 2.030764f
C482 SUNSAR_SAR8B_CV_0/XA2/XA2/MN0/a_324_n18# 0 0.360407f
C483 SUNSAR_SAR8B_CV_0/XA2/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C484 SUNSAR_SAR8B_CV_0/XA2/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C485 SUNSAR_SAR8B_CV_0/XA2/XA1/XA2/Y 0 1.060197f
C486 SUNSAR_SAR8B_CV_0/XA2/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C487 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C488 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C489 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C490 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MP3/G 0 0.827484f
C491 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN2/S 0 0.200627f
C492 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C493 SUNSAR_SAR8B_CV_0/XA3/EN 0 3.784028f
C494 SUNSAR_SAR8B_CV_0/XA2/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C495 SUNSAR_SAR8B_CV_0/XA2/XA13/MN1/a_324_334# 0 0.422f
C496 SUNSAR_SAR8B_CV_0/XA2/XA12/MN0/a_324_n18# 0 0.360407f
C497 SUNSAR_SAR8B_CV_0/XA2/XA13/MN1/a_324_n18# 0 0.360407f
C498 SUNSAR_SAR8B_CV_0/XA2/XA12/A 0 0.755669f
C499 SUNSAR_SAR8B_CV_0/XA2/XA11/MN0/a_324_n18# 0 0.360407f
C500 SUNSAR_SAR8B_CV_0/XA1/CEO 0 1.104751f
C501 SUNSAR_SAR8B_CV_0/XA2/XA11/A 0 0.662715f
C502 SUNSAR_SAR8B_CV_0/XA2/XA9/Y 0 0.718246f
C503 SUNSAR_SAR8B_CV_0/XA1/XA9/MN1/a_324_334# 0 0.360407f
C504 SUNSAR_SAR8B_CV_0/XA1/XA9/MN0/a_324_n18# 0 0.360407f
C505 SUNSAR_SAR8B_CV_0/XA1/XA9/A 0 1.250075f
C506 SUNSAR_SAR8B_CV_0/XA1/DONE 0 0.123486f
C507 SUNSAR_SAR8B_CV_0/XA1/XA7/MN0/a_324_n18# 0 0.360407f
C508 SUNSAR_SAR8B_CV_0/XA1/XA8/MN0/a_324_n18# 0 0.360407f
C509 SUNSAR_SAR8B_CV_0/XA1/XA9/B 0 1.158058f
C510 SUNSAR_SAR8B_CV_0/XA1/XA6/MN0/a_324_n18# 0 0.360407f
C511 SUNSAR_SAR8B_CV_0/XA1/XA4/A 0 2.621765f
C512 SUNSAR_SAR8B_CV_0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C513 SUNSAR_SAR8B_CV_0/XA1/CP0 0 4.486094f
C514 SUNSAR_SAR8B_CV_0/XA1/CN0 0 2.798774f
C515 SUNSAR_SAR8B_CV_0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C516 SUNSAR_SAR8B_CV_0/XA1/CN1 0 4.70217f
C517 SUNSAR_SAR8B_CV_0/D<6> 0 4.492109f
C518 SUNSAR_SAR8B_CV_0/XA1/XA3/MN0/a_324_n18# 0 0.360407f
C519 SUNSAR_SAR8B_CV_0/XA1/XA2/A 0 2.030764f
C520 SUNSAR_SAR8B_CV_0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C521 SUNSAR_SAR8B_CV_0/XA1/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C522 SUNSAR_SAR8B_CV_0/XA1/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C523 SUNSAR_SAR8B_CV_0/XA1/XA1/XA2/Y 0 1.060197f
C524 SUNSAR_SAR8B_CV_0/XA1/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C525 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C526 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C527 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C528 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MP3/G 0 0.827484f
C529 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN2/S 0 0.200627f
C530 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C531 SUNSAR_SAR8B_CV_0/XA2/EN 0 3.720665f
C532 SUNSAR_SAR8B_CV_0/XA1/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C533 SUNSAR_SAR8B_CV_0/XA1/XA13/MN1/a_324_334# 0 0.422f
C534 SUNSAR_SAR8B_CV_0/XA1/XA12/MN0/a_324_n18# 0 0.360407f
C535 SUNSAR_SAR8B_CV_0/XA1/XA13/MN1/a_324_n18# 0 0.360407f
C536 SUNSAR_SAR8B_CV_0/XA1/XA12/A 0 0.755669f
C537 SUNSAR_SAR8B_CV_0/XA1/XA11/MN0/a_324_n18# 0 0.360407f
C538 SUNSAR_SAR8B_CV_0/XA0/CEO 0 1.083361f
C539 SUNSAR_SAR8B_CV_0/XA1/XA11/A 0 0.662715f
C540 SUNSAR_SAR8B_CV_0/XA1/XA9/Y 0 0.718246f
C541 SUNSAR_SAR8B_CV_0/XB2/XA7/MN1/a_324_n18# 0 0.359583f
C542 SUNSAR_SAR8B_CV_0/XB2/XA5b/MN1/a_324_n18# 0 0.422415f
C543 SUNSAR_SAR8B_CV_0/XB2/XA1/Y 0 0.690197f
C544 SUNSAR_SAR8B_CV_0/XB2/CKN 0 1.768971f
C545 SUNSAR_SAR8B_CV_0/XB2/XA4/MN0/a_324_n18# 0 0.359583f
C546 SUNSAR_SAR8B_CV_0/XB2/XA5/MN1/a_324_334# 0 0.422f
C547 SUNSAR_SAR8B_CV_0/XB2/XA3/MP0/S 0 0.743486f
C548 SUNSAR_SAR8B_CV_0/XB2/XA3/MN0/a_324_n18# 0 0.359583f
C549 SUNSAR_SAR8B_CV_0/XB2/XA2/MP0/G 0 0.708335f
C550 SUNSAR_SAR8B_CV_0/XB2/XA7/MN1/a_324_334# 0 0.359583f
C551 SUNSAR_SAR8B_CV_0/XB2/XA5/MN1/a_324_n18# 0 0.360407f
C552 SUNSAR_SAR8B_CV_0/XB2/XA1/MP0/G 0 0.788614f
C553 SUNSAR_SAR8B_CV_0/XB2/XA4/MN1/a_324_334# 0 0.359583f
C554 SUNSAR_SAR8B_CV_0/XB2/XA0/MN0/a_324_n18# 0 0.359583f
C555 SUNSAR_SAR8B_CV_0/XB2/M8/a_324_n18# 0 0.356977f
C556 SUNSAR_SAR8B_CV_0/XB2/M8/a_324_334# 0 0.422f
C557 SUNSAR_SAR8B_CV_0/XB2/M6/a_324_n18# 0 0.356977f
C558 SUNSAR_SAR8B_CV_0/XB2/M7/a_324_n18# 0 0.356977f
C559 SUNSAR_SAR8B_CV_0/XB2/XA3/B 0 54.41209f
C560 SUNSAR_SAR8B_CV_0/XB2/XA4/GNG 0 53.065117f
C561 SUNSAR_SAR8B_CV_0/XB2/M5/a_324_n18# 0 0.356977f
C562 SUNSAR_SAR8B_CV_0/XB2/M3/a_324_n18# 0 0.356977f
C563 SUNSAR_SAR8B_CV_0/XB2/M4/a_324_n18# 0 0.356977f
C564 SUNSAR_SAR8B_CV_0/XB2/M4/G 0 2.475647f
C565 ua[0] 0 2.335287f
C566 SUNSAR_SAR8B_CV_0/XB2/M1/a_324_n18# 0 0.422415f
C567 SUNSAR_SAR8B_CV_0/XB2/M2/a_324_n18# 0 0.356977f
C568 SUNSAR_SAR8B_CV_0/XA0/XA9/MN1/a_324_334# 0 0.360407f
C569 SUNSAR_SAR8B_CV_0/XA0/XA9/MN0/a_324_n18# 0 0.360407f
C570 SUNSAR_SAR8B_CV_0/XA0/XA9/A 0 1.250075f
C571 SUNSAR_SAR8B_CV_0/XA0/DONE 0 0.134046f
C572 SUNSAR_SAR8B_CV_0/XA0/XA7/MN0/a_324_n18# 0 0.360407f
C573 SUNSAR_SAR8B_CV_0/XA0/XA8/MN0/a_324_n18# 0 0.360407f
C574 SUNSAR_SAR8B_CV_0/XA0/XA9/B 0 1.158058f
C575 SUNSAR_SAR8B_CV_0/CK_SAMPLE 0 17.082773f
C576 SUNSAR_SAR8B_CV_0/XA0/XA6/MN0/a_324_n18# 0 0.360407f
C577 SUNSAR_SAR8B_CV_0/XA0/XA4/A 0 2.621765f
C578 SUNSAR_SAR8B_CV_0/XA0/XA4/MN0/a_324_n18# 0 0.360407f
C579 SUNSAR_SAR8B_CV_0/XA0/CP0 0 8.48089f
C580 SUNSAR_SAR8B_CV_0/XA0/XA5/MN0/a_324_n18# 0 0.360407f
C581 SUNSAR_SAR8B_CV_0/D<7> 0 9.577809f
C582 SUNSAR_SAR8B_CV_0/XA0/XA3/MN0/a_324_n18# 0 0.360407f
C583 SUNSAR_SAR8B_CV_0/XA0/XA2/A 0 2.030764f
C584 SUNSAR_SAR8B_CV_0/XA0/XA2/MN0/a_324_n18# 0 0.360407f
C585 SUNSAR_SAR8B_CV_0/XA20/CNO 0 12.667546f
C586 SUNSAR_SAR8B_CV_0/XA0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C587 SUNSAR_SAR8B_CV_0/EN 0 5.988511f
C588 SUNSAR_SAR8B_CV_0/XA0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C589 SUNSAR_SAR8B_CV_0/XA0/XA1/XA2/Y 0 1.060197f
C590 SUNSAR_SAR8B_CV_0/XA0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C591 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C592 SUNSAR_SAR8B_CV_0/XA20/CPO 0 11.091676f
C593 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C594 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C595 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MP3/G 0 0.827484f
C596 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN2/S 0 0.200627f
C597 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C598 SUNSAR_SAR8B_CV_0/XA1/EN 0 3.794638f
C599 SUNSAR_SAR8B_CV_0/XA0/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C600 VPWR 0 0.724262p
C601 SUNSAR_SAR8B_CV_0/XA0/XA13/MN1/a_324_334# 0 0.422f
C602 SUNSAR_SAR8B_CV_0/XA0/XA12/MN0/a_324_n18# 0 0.360407f
C603 SUNSAR_SAR8B_CV_0/XA0/XA13/MN1/a_324_n18# 0 0.360407f
C604 SUNSAR_SAR8B_CV_0/XA0/XA12/A 0 0.755669f
C605 SUNSAR_SAR8B_CV_0/XA0/XA11/MN0/a_324_n18# 0 0.360407f
C606 SUNSAR_SAR8B_CV_0/XA0/XA11/A 0 0.662715f
C607 SUNSAR_SAR8B_CV_0/XA0/XA9/Y 0 0.718246f
C608 SUNSAR_SAR8B_CV_0/XB1/XA7/MN1/a_324_n18# 0 0.359583f
C609 VGND 0 0.219536p
C610 SUNSAR_SAR8B_CV_0/XB1/XA5b/MN1/a_324_n18# 0 0.422415f
C611 SUNSAR_SAR8B_CV_0/XB1/XA1/Y 0 0.690197f
C612 SUNSAR_SAR8B_CV_0/XB1/CKN 0 1.768971f
C613 SUNSAR_SAR8B_CV_0/XB1/XA4/MN0/a_324_n18# 0 0.359583f
C614 SUNSAR_SAR8B_CV_0/XB1/XA5/MN1/a_324_334# 0 0.422f
C615 SUNSAR_SAR8B_CV_0/XB1/XA3/MP0/S 0 0.743486f
C616 SUNSAR_SAR8B_CV_0/XB1/XA3/MN0/a_324_n18# 0 0.359583f
C617 SUNSAR_SAR8B_CV_0/XB1/XA2/MP0/G 0 0.708335f
C618 SUNSAR_SAR8B_CV_0/XB1/XA7/MN1/a_324_334# 0 0.359583f
C619 SUNSAR_SAR8B_CV_0/XB1/XA5/MN1/a_324_n18# 0 0.360407f
C620 SUNSAR_SAR8B_CV_0/XB1/XA1/MP0/G 0 0.788614f
C621 SUNSAR_SAR8B_CV_0/XB1/XA4/MN1/a_324_334# 0 0.359583f
C622 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0 6.475628f
C623 SUNSAR_SAR8B_CV_0/XB1/XA0/MN0/a_324_n18# 0 0.359583f
C624 SUNSAR_SAR8B_CV_0/XB1/M8/a_324_n18# 0 0.356977f
C625 SUNSAR_SAR8B_CV_0/XB1/M8/a_324_334# 0 0.422f
C626 SUNSAR_SAR8B_CV_0/XB1/M6/a_324_n18# 0 0.356977f
C627 SUNSAR_SAR8B_CV_0/XB1/M7/a_324_n18# 0 0.356977f
C628 SUNSAR_SAR8B_CV_0/XB1/XA3/B 0 54.41209f
C629 SUNSAR_SAR8B_CV_0/XB1/XA4/GNG 0 53.065117f
C630 SUNSAR_SAR8B_CV_0/XA0/CEIN 0 19.901903f
C631 SUNSAR_SAR8B_CV_0/XB1/M5/a_324_n18# 0 0.356977f
C632 SUNSAR_SAR8B_CV_0/XB1/M3/a_324_n18# 0 0.356977f
C633 SUNSAR_SAR8B_CV_0/XB1/M4/a_324_n18# 0 0.356977f
C634 SUNSAR_SAR8B_CV_0/XB1/M4/G 0 2.475647f
C635 ua[1] 0 3.007717f
C636 SUNSAR_SAR8B_CV_0/XB1/M1/a_324_n18# 0 0.422415f
C637 SUNSAR_SAR8B_CV_0/XB1/M2/a_324_n18# 0 0.356977f
C638 SUNSAR_SAR8B_CV_0/XA20/XA9/MN0/a_324_n18# 0 0.360407f
C639 SUNSAR_SAR8B_CV_0/XA20/XA3/CO 0 2.703497f
C640 SUNSAR_SAR8B_CV_0/XA20/XA2/MN6/a_324_334# 0 0.360407f
C641 SUNSAR_SAR8B_CV_0/XA20/XA3a/A 0 2.536943f
C642 SUNSAR_SAR8B_CV_0/XA20/XA3/MN0/a_324_n18# 0 0.360407f
C643 SUNSAR_SAR8B_CV_0/XA20/XA3a/MN0/a_324_n18# 0 0.360407f
C644 SUNSAR_SAR8B_CV_0/XA20/XA4/MN0/a_324_n18# 0 0.360407f
C645 SUNSAR_SAR8B_CV_0/XA20/XA4/MP0/S 0 0.397005f
C646 SUNSAR_SAR8B_CV_0/SARN 0 30.043571f
C647 SUNSAR_SAR8B_CV_0/XA20/XA3/N2 0 0.234927f
C648 SUNSAR_SAR8B_CV_0/XA20/XA9/Y 0 3.176436f
C649 SUNSAR_SAR8B_CV_0/XA20/XA2/N2 0 0.234927f
C650 SUNSAR_SAR8B_CV_0/XA20/XA2/MN0/a_324_n18# 0 0.360407f
C651 SUNSAR_SAR8B_CV_0/XA20/XA3/N1 0 0.905385f
C652 SUNSAR_SAR8B_CV_0/SARP 0 30.653925f
C653 SUNSAR_SAR8B_CV_0/XA20/XA1/MN0/a_324_n18# 0 0.360407f
C654 SUNSAR_SAR8B_CV_0/XA20/XA1/MP0/S 0 0.397005f
C655 SUNSAR_SAR8B_CV_0/XA20/XA9/A 0 3.508213f
C656 SUNSAR_SAR8B_CV_0/XA20/XA0/MN1/a_324_n18# 0 0.422415f
C657 SUNSAR_SAR8B_CV_0/XA20/XA13/MN1/a_324_n18# 0 0.360407f
C658 SUNSAR_SAR8B_CV_0/XA20/XA13/MN1/a_324_334# 0 0.422f
C659 SUNSAR_SAR8B_CV_0/XA7/CEO 0 1.316615f
C660 SUNSAR_SAR8B_CV_0/XA20/XA12/MN0/a_324_n18# 0 0.360407f
C661 SUNSAR_SAR8B_CV_0/XA20/XA11/MN0/a_324_n18# 0 0.360407f
C662 SUNSAR_SAR8B_CV_0/XA20/XA9/MN0/a_324_334# 0 0.360407f
C663 SUNSAR_SAR8B_CV_0/XA20/XA12/Y 0 0.623343f
C664 SUNSAR_SAR8B_CV_0/XA20/XA11/Y 0 0.759616f
C665 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES2/B 0 3.1129f
C666 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES4/B 0 3.516117f
C667 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES8/B 0 3.933522f
C668 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES16/B 0 4.664508f
C669 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES1B/B 0 2.892833f
C670 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES1A/B 0 1.735354f
C671 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES2/B 0 3.1129f
C672 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES4/B 0 3.516117f
C673 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES8/B 0 3.933522f
C674 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES16/B 0 4.664508f
C675 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES1B/B 0 2.892833f
C676 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES1A/B 0 1.735354f
C677 SUNSAR_SAR8B_CV_0/XA0/CN0 0 6.776559f
C678 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES2/B 0 3.1129f
C679 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES4/B 0 3.516117f
C680 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES8/B 0 3.933522f
C681 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES16/B 0 4.664508f
C682 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES1B/B 0 2.892833f
C683 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES1A/B 0 1.735354f
C684 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES2/B 0 3.1129f
C685 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES4/B 0 3.516117f
C686 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES8/B 0 3.933522f
C687 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES16/B 0 4.664508f
C688 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES1B/B 0 2.892833f
C689 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES1A/B 0 1.735354f
C690 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES2/B 0 3.1129f
C691 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES4/B 0 3.516117f
C692 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES8/B 0 3.933522f
C693 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES16/B 0 4.664508f
C694 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES1B/B 0 2.892833f
C695 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES1A/B 0 1.735354f
C696 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES2/B 0 3.1129f
C697 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES4/B 0 3.516117f
C698 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES8/B 0 3.933522f
C699 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES16/B 0 4.664508f
C700 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES1B/B 0 2.892833f
C701 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES1A/B 0 1.735354f
C702 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES2/B 0 3.1129f
C703 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES4/B 0 3.516117f
C704 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES8/B 0 3.933522f
C705 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES16/B 0 4.664508f
C706 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES1B/B 0 2.892833f
C707 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES1A/B 0 1.735354f
C708 SUNSAR_SAR8B_CV_0/D<5> 0 5.830972f
C709 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES2/B 0 3.1129f
C710 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES4/B 0 3.516117f
C711 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES8/B 0 3.933522f
C712 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES16/B 0 4.664508f
C713 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES1B/B 0 2.892833f
C714 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES1A/B 0 1.735354f
C715 SUNSAR_SAR8B_CV_0/XA0/CP1 0 4.930175f
C716 tt_um_TT06_SAR_done_0/x5/MN1/a_324_334# 0 0.422f
C717 tt_um_TT06_SAR_done_0/x4/MP0/G 0 0.782647f
C718 tt_um_TT06_SAR_done_0/x5/MN1/a_324_n18# 0 0.360407f
C719 uio_oe[0] 0 1.630684f
C720 uio_out[0] 0 1.156269f
C721 tt_um_TT06_SAR_done_0/x3/MN1/a_324_n18# 0 0.355196f
C722 tt_um_TT06_SAR_done_0/x4/MN0/a_324_n18# 0 0.360407f
C723 tt_um_TT06_SAR_done_0/x3/MP1/G 0 0.95314f
C724 tt_um_TT06_SAR_done_0/x3/MN0/a_324_n18# 0 0.422415f
.ends

