* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

.subckt TT06SAR_NDIO a_n147_n147# a_n45_n45#
D0 a_n147_n147# a_n45_n45# sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
C0 a_n45_n45# a_n147_n147# 0.450369f
.ends

.subckt SUNTR_PCHDL D G S B 0 a_216_n18# a_216_334#
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 B G 0.33939f
C1 a_216_n18# G 0.067434f
C2 a_216_334# G 0.065834f
C3 a_216_n18# B 0.330729f
C4 a_216_334# B 0.331144f
C5 G 0 0.072524f
C6 B 0 2.80592f
C7 a_216_n18# 0 0.091271f
C8 a_216_334# 0 0.091271f
.ends

.subckt SUNTR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 a_324_334# G 0.067434f
C1 a_324_n18# G 0.065834f
C2 S B 0.06295f
C3 G B 0.411913f
C4 D B 0.06295f
C5 a_324_n18# B 0.422415f
C6 a_324_334# B 0.422f
.ends

.subckt SUNTR_BFX1_CV Y AVDD AVSS MP1/B MN1/a_324_334# MP1/G A 0 MP1/a_216_334#
XMP0 AVDD A MP1/G MP1/B 0 MP0/a_216_n18# MP1/a_216_n18# SUNTR_PCHDL
XMP1 Y MP1/G AVDD MP1/B 0 MP1/a_216_n18# MP1/a_216_334# SUNTR_PCHDL
XMN0 AVSS A MP1/G 0 MN0/a_324_n18# MN1/a_324_n18# SUNTR_NCHDL
XMN1 Y MP1/G AVSS 0 MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 AVDD MP1/B 0.181063f
C1 Y MP1/B 0.063474f
C2 AVSS AVDD 0.10499f
C3 MP1/G MP1/B 0.178777f
C4 A MP1/B 0.109691f
C5 MP1/G AVDD 0.062148f
C6 MP1/G AVSS 0.120067f
C7 MP1/G Y 0.07318f
C8 A MP1/G 0.156853f
C9 MP1/B MP1/a_216_n18# -0.310513f
C10 AVDD 0 0.276075f
C11 AVSS 0 0.45436f
C12 Y 0 0.218882f
C13 MN1/a_324_n18# 0 0.351938f
C14 MN1/a_324_334# 0 0.422f
C15 MP1/G 0 0.969276f
C16 A 0 0.55997f
C17 MN0/a_324_n18# 0 0.422415f
C18 MP1/a_216_334# 0 0.091338f
C19 MP1/B 0 4.386796f
C20 MP0/a_216_n18# 0 0.091338f
.ends

.subckt SUNTR_TIEH_CV Y AVDD AVSS MP0/B MP0/G 0 MP0/a_216_334# MP0/a_216_n18# MN0/a_324_n18#
+ MN0/a_324_334#
XMP0 Y MP0/G AVDD MP0/B 0 MP0/a_216_n18# MP0/a_216_334# SUNTR_PCHDL
XMN0 MP0/G MP0/G AVSS 0 MN0/a_324_n18# MN0/a_324_334# SUNTR_NCHDL
C0 AVSS AVDD 0.052497f
C1 AVSS MP0/G 0.060387f
C2 AVDD MP0/B 0.112171f
C3 MP0/B MP0/G 0.112479f
C4 AVDD 0 0.260853f
C5 AVSS 0 0.382267f
C6 MP0/G 0 0.78444f
C7 MN0/a_324_n18# 0 0.422415f
C8 MN0/a_324_334# 0 0.422f
C9 MP0/B 0 2.80738f
C10 MP0/a_216_n18# 0 0.091338f
C11 MP0/a_216_334# 0 0.091338f
.ends

.subckt SUNTR_TAPCELLB_CV AVDD AVSS MN1/a_324_n18# MP1/a_216_n18#
XMP1 AVDD AVDD AVDD AVDD AVSS MP1/a_216_n18# MP1/a_216_334# SUNTR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNTR_NCHDL
C0 AVDD AVSS 0.107602f
C1 AVSS 0 1.064147f
C2 MN1/a_324_n18# 0 0.422415f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.146627f
C5 MP1/a_216_n18# 0 0.091271f
C6 MP1/a_216_334# 0 0.091271f
.ends

.subckt tt_um_TT06_SAR_done DONE uio_out<0> uio_oe<0> VPWR VGND
Xx3 uio_out<0> VPWR VGND VPWR x4/MN0/a_324_n18# x3/MP1/G DONE VGND x4/MP0/a_216_n18#
+ SUNTR_BFX1_CV
Xx4 uio_oe<0> VPWR VGND VPWR x4/MP0/G VGND x5/MP1/a_216_n18# x4/MP0/a_216_n18# x4/MN0/a_324_n18#
+ x5/MN1/a_324_n18# SUNTR_TIEH_CV
Xx5 VPWR VGND x5/MN1/a_324_n18# x5/MP1/a_216_n18# SUNTR_TAPCELLB_CV
C0 uio_oe<0> VPWR 0.524617f
C1 x3/MP1/G x4/MP0/G 0.071481f
C2 x3/MP1/G uio_out<0> 0.07263f
C3 DONE uio_out<0> 0.05692f
C4 DONE VGND 0.094224f
C5 VGND x4/MP0/G 0.114893f
C6 VGND uio_out<0> 0.294473f
C7 x4/MP0/a_216_n18# VPWR -0.31151f
C8 VPWR uio_out<0> 0.077974f
C9 VPWR x5/MP1/a_216_n18# -0.314359f
C10 uio_oe<0> x4/MP0/G 0.055797f
C11 VGND 0 0.898244f
C12 x5/MN1/a_324_334# 0 0.422f
C13 VPWR 0 7.717914f
C14 x5/MP1/a_216_334# 0 0.091271f
C15 x4/MP0/G 0 0.782647f
C16 x5/MN1/a_324_n18# 0 0.360407f
C17 uio_oe<0> 0 0.133144f
C18 uio_out<0> 0 0.357519f
C19 x3/MN1/a_324_n18# 0 0.355196f
C20 x4/MN0/a_324_n18# 0 0.360407f
C21 x3/MP1/G 0 0.95314f
C22 DONE 0 0.720744f
C23 x3/MN0/a_324_n18# 0 0.422415f
C24 x3/MP0/a_216_n18# 0 0.091271f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_XS736D c1_n1946_n17480# m3_n1986_n17520# 0
X0 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X1 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X2 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X3 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X4 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X5 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X6 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X7 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X8 c1_n1946_n17480# m3_n1986_n17520# sky130_fd_pr__cap_mim_m3_1 l=18 w=18
C0 c1_n1946_n17480# m3_n1986_n17520# 0.265161p
C1 c1_n1946_n17480# 0 9.109429f
C2 m3_n1986_n17520# 0 65.3375f
.ends

.subckt SUNSAR_RM1 A B 0
R0 A B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
.ends

.subckt SUNSAR_CAP32C_CV C1B C2 C4 C16 CTOP AVSS C1A XRES1A/B C8 0 XRES1B/B
XXRES16 C16 XRES16/B 0 SUNSAR_RM1
XXRES2 C2 XRES2/B 0 SUNSAR_RM1
XXRES1A C1A XRES1A/B 0 SUNSAR_RM1
XXRES4 C4 XRES4/B 0 SUNSAR_RM1
XXRES1B C1B XRES1B/B 0 SUNSAR_RM1
XXRES8 C8 XRES8/B 0 SUNSAR_RM1
C0 XRES1A/B CTOP 3.552515f
C1 XRES8/B XRES2/B 0.419738f
C2 XRES8/B XRES4/B 0.449585f
C3 XRES16/B XRES2/B 0.441867f
C4 AVSS XRES2/B 4.083764f
C5 XRES16/B XRES4/B 0.058243f
C6 AVSS XRES4/B 4.927044f
C7 XRES16/B XRES8/B 0.098257f
C8 AVSS XRES8/B 6.541971f
C9 AVSS XRES16/B 9.801106f
C10 XRES1B/B XRES4/B 0.40569f
C11 XRES1B/B AVSS 3.75982f
C12 XRES2/B CTOP 6.866754f
C13 XRES4/B CTOP 13.651895f
C14 XRES1A/B XRES16/B 0.437694f
C15 XRES8/B CTOP 27.161474f
C16 XRES1A/B AVSS 3.7558f
C17 XRES16/B CTOP 54.216488f
C18 AVSS CTOP 9.918657f
C19 XRES1B/B CTOP 3.552515f
C20 CTOP 0 7.76011f
C21 XRES2/B 0 3.1129f
C22 XRES4/B 0 3.516117f
C23 XRES8/B 0 3.933522f
C24 XRES16/B 0 4.664508f
C25 AVSS 0 15.179144f
C26 C8 0 0.101745f
C27 XRES1B/B 0 2.892833f
C28 C1B 0 0.116997f
C29 C4 0 0.101745f
C30 XRES1A/B 0 1.735354f
C31 C1A 0 0.116997f
C32 C2 0 0.101745f
C33 C16 0 0.101745f
.ends

.subckt SUNSAR_CDAC7_CV CP<9> CP<8> CP<7> CP<6> CP<5> CP<4> CP<3> CP<2> CP<1> CP<0>
+ CTOP 0 AVSS
XX16ab CP<5> CP<5> CP<5> CP<6> CTOP AVSS CP<5> X16ab/XRES1A/B CP<4> 0 X16ab/XRES1B/B
+ SUNSAR_CAP32C_CV
XXC0 CP<9> CP<9> CP<9> CP<9> CTOP AVSS CP<9> XC0/XRES1A/B CP<9> 0 XC0/XRES1B/B SUNSAR_CAP32C_CV
XXC1 CP<8> CP<8> CP<8> CP<8> CTOP AVSS CP<8> XC1/XRES1A/B CP<8> 0 XC1/XRES1B/B SUNSAR_CAP32C_CV
XXC32a<0> CP<0> CP<1> CP<2> CP<7> CTOP AVSS AVSS XC32a<0>/XRES1A/B CP<3> 0 XC32a<0>/XRES1B/B
+ SUNSAR_CAP32C_CV
C0 CP<6> CP<5> 2.020583f
C1 CP<2> CP<0> 0.24075f
C2 XC32a<0>/XRES1A/B AVSS 0.082248f
C3 CP<1> CP<7> 0.188755f
C4 CP<8> AVSS 0.71211f
C5 CP<0> CP<8> 0.088104f
C6 CP<2> CP<8> 0.089552f
C7 CP<9> CTOP 0.074555f
C8 CP<1> CP<3> 0.220707f
C9 CP<9> CP<5> 0.103206f
C10 XC1/XRES1B/B AVSS 0.082248f
C11 XC1/XRES1B/B XC32a<0>/XRES1A/B 0.635098f
C12 X16ab/XRES1B/B XC0/XRES1A/B 0.635098f
C13 CP<0> CP<7> 0.081678f
C14 AVSS CTOP -1.633715f
C15 CP<5> AVSS 0.068641f
C16 CP<5> CP<0> 0.20259f
C17 CP<2> CP<7> 0.083155f
C18 CP<4> CP<8> 0.089689f
C19 CP<7> CP<8> 2.575701f
C20 CP<0> CP<3> 0.084671f
C21 X16ab/XRES1B/B AVSS 0.082248f
C22 CP<8> CTOP 0.122672f
C23 CP<5> CP<8> 0.359484f
C24 CP<2> CP<3> 2.212231f
C25 CP<0> CP<1> 1.909476f
C26 CP<3> CP<8> 0.0896f
C27 X16ab/XRES1A/B XC32a<0>/XRES1B/B 0.635098f
C28 X16ab/XRES1A/B AVSS 0.082248f
C29 CP<6> CP<8> 0.090483f
C30 CP<2> CP<1> 1.995553f
C31 CP<4> CP<7> 0.07877f
C32 XC0/XRES1A/B AVSS 0.082248f
C33 CP<5> CP<4> 1.57931f
C34 CP<5> CP<7> 0.394951f
C35 CP<9> AVSS 0.343312f
C36 CP<1> CP<8> 0.089524f
C37 CP<4> CP<3> 1.263888f
C38 CP<3> CP<7> 0.178438f
C39 CP<6> CP<4> 0.07931f
C40 XC32a<0>/XRES1B/B AVSS 0.082248f
C41 CP<6> CP<7> 1.652261f
C42 CP<5> CP<3> 0.229397f
C43 CP<9> CP<8> 0.889573f
C44 XC32a<0>/XRES2/B 0 3.1129f
C45 XC32a<0>/XRES4/B 0 3.516117f
C46 XC32a<0>/XRES8/B 0 3.933522f
C47 XC32a<0>/XRES16/B 0 4.664508f
C48 CP<3> 0 1.126461f
C49 XC32a<0>/XRES1B/B 0 2.892833f
C50 CP<0> 0 1.167979f
C51 CP<2> 0 0.834649f
C52 XC32a<0>/XRES1A/B 0 1.735354f
C53 CP<1> 0 1.392542f
C54 CP<7> 0 1.060384f
C55 CTOP 0 20.24516f
C56 XC1/XRES2/B 0 3.1129f
C57 XC1/XRES4/B 0 3.516117f
C58 XC1/XRES8/B 0 3.933522f
C59 XC1/XRES16/B 0 4.664508f
C60 AVSS 0 51.996902f
C61 XC1/XRES1B/B 0 2.892833f
C62 XC1/XRES1A/B 0 1.735354f
C63 CP<8> 0 3.823549f
C64 XC0/XRES2/B 0 3.1129f
C65 XC0/XRES4/B 0 3.516117f
C66 XC0/XRES8/B 0 3.933522f
C67 XC0/XRES16/B 0 4.664508f
C68 XC0/XRES1B/B 0 2.892833f
C69 XC0/XRES1A/B 0 1.735354f
C70 CP<5> 0 2.378288f
C71 X16ab/XRES2/B 0 3.1129f
C72 X16ab/XRES4/B 0 3.516117f
C73 X16ab/XRES8/B 0 3.933522f
C74 X16ab/XRES16/B 0 4.664508f
C75 CP<4> 0 0.757332f
C76 X16ab/XRES1B/B 0 2.892833f
C77 X16ab/XRES1A/B 0 1.735354f
C78 CP<6> 0 0.645761f
C79 CP<9> 0 2.290488f
.ends

.subckt SUNSAR_PCHDL D G S B 0 a_216_n18# a_216_334#
X0 D G S B sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 D S 0.050207f
C1 B G 0.341895f
C2 a_216_n18# G 0.067588f
C3 a_216_334# G 0.066018f
C4 a_216_n18# B 0.330729f
C5 a_216_334# B 0.331144f
C6 G 0 0.073301f
C7 B 0 2.80584f
C8 a_216_n18# 0 0.091271f
C9 a_216_334# 0 0.091271f
.ends

.subckt SUNSAR_NCHDL D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 D S 0.050207f
C1 a_324_n18# G 0.066018f
C2 a_324_334# G 0.067588f
C3 S B 0.06638f
C4 G B 0.415197f
C5 D B 0.06638f
C6 a_324_n18# B 0.422415f
C7 a_324_334# B 0.422f
.ends

.subckt SUNSAR_NDX1_CV Y AVDD AVSS MN1/a_324_334# B A BULKP BULKN MP0/a_216_n18# MN1/S
+ MP1/a_216_334# MN0/a_324_n18#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# B SUNSAR_PCHDL
XMP1 AVDD B Y BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 MN1/S A AVSS BULKN MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 Y B MN1/S BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 B Y 0.059989f
C1 BULKP B -0.247362f
C2 A BULKP -0.246413f
C3 AVDD AVSS 0.070991f
C4 Y AVDD 0.077947f
C5 BULKP AVDD 0.154562f
C6 AVSS BULKN 0.392705f
C7 MN1/a_324_334# BULKN 0.422f
C8 AVDD BULKN 0.326781f
C9 MN0/a_324_n18# BULKN 0.422415f
C10 Y BULKN 0.252959f
C11 B BULKN 0.538316f
C12 BULKP BULKN 3.595959f
C13 A BULKN 0.53919f
C14 MP1/a_216_334# BULKN 0.091338f
C15 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_NRX1_CV AVDD AVSS MN1/a_324_334# B BULKP BULKN MP0/a_216_n18# Y MP1/a_216_334#
+ A MN0/a_324_n18#
XMP0 MP1/S A AVDD BULKP BULKN MP0/a_216_n18# B SUNSAR_PCHDL
XMP1 Y B MP1/S BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# B SUNSAR_NCHDL
XMN1 AVSS B Y BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.122023f
C1 BULKP B -0.247362f
C2 A BULKP -0.246413f
C3 Y AVSS 0.112939f
C4 AVDD AVSS 0.071423f
C5 B Y 0.059989f
C6 BULKP Y 0.076318f
C7 AVSS BULKN 0.506278f
C8 Y BULKN 0.247181f
C9 MN1/a_324_334# BULKN 0.422f
C10 MN0/a_324_n18# BULKN 0.422415f
C11 AVDD BULKN 0.25764f
C12 B BULKN 0.538314f
C13 BULKP BULKN 3.595964f
C14 MP1/a_216_334# BULKN 0.091338f
C15 A BULKN 0.539194f
C16 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_IVX1_CV BULKP AVSS Y BULKN MP0/a_216_n18# MP0/a_216_334# AVDD A MN0/a_324_n18#
+ MN0/a_324_334#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.051104f
C1 BULKP A 0.109299f
C2 BULKP Y 0.061437f
C3 BULKP AVDD 0.103136f
C4 AVSS BULKN 0.367376f
C5 A BULKN 0.631634f
C6 Y BULKN 0.268384f
C7 MN0/a_324_n18# BULKN 0.422415f
C8 MN0/a_324_334# BULKN 0.422f
C9 AVDD BULKN 0.246592f
C10 BULKP BULKN 2.80697f
C11 MP0/a_216_n18# BULKN 0.091338f
C12 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TAPCELLB_CV AVDD MN1/a_324_n18# MN1/a_324_334# AVSS MP1/a_216_334#
+ MP1/a_216_n18#
XMP1 AVDD AVDD AVDD AVDD AVSS MP1/a_216_n18# MP1/a_216_334# SUNSAR_PCHDL
XMN1 AVSS AVSS AVSS AVSS MN1/a_324_n18# MN1/a_324_334# SUNSAR_NCHDL
C0 AVDD AVSS 0.104949f
C1 AVSS 0 1.048908f
C2 MN1/a_324_n18# 0 0.422415f
C3 MN1/a_324_334# 0 0.422f
C4 AVDD 0 3.134387f
C5 MP1/a_216_n18# 0 0.091271f
C6 MP1/a_216_334# 0 0.091271f
.ends

.subckt SUNSAR_SARKICKHX1_CV CI BULKP AVDD AVSS MP6_DMY/a_216_334# MN6/a_324_334#
+ MP0/S CKN MP0/a_216_n18# CK BULKN MN0/a_324_n18#
XMP1_DMY AVDD AVDD AVDD BULKP BULKN CKN AVDD SUNSAR_PCHDL
XMP4_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP0 AVDD CKN MP0/S BULKP BULKN MP0/a_216_n18# AVDD SUNSAR_PCHDL
XMN0 MP0/S CKN AVSS BULKN MN0/a_324_n18# CI SUNSAR_NCHDL
XMN1 MP0/S CI MP0/S BULKN CKN CI SUNSAR_NCHDL
XMN2 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN3 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN4 MP0/S CI MP0/S BULKN CI CI SUNSAR_NCHDL
XMN6 AVDD CK MP0/S BULKN CI MN6/a_324_334# SUNSAR_NCHDL
XMN5 MP0/S CI MP0/S BULKN CI CK SUNSAR_NCHDL
XMP3_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP6_DMY AVDD AVDD AVDD BULKP BULKN AVDD MP6_DMY/a_216_334# SUNSAR_PCHDL
XMP2_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
XMP5_DMY AVDD AVDD AVDD BULKP BULKN AVDD AVDD SUNSAR_PCHDL
C0 AVSS AVDD 0.180248f
C1 CKN MP0/S 0.058228f
C2 MP0/S AVDD 0.104608f
C3 MP0/S BULKP 0.11694f
C4 AVSS CI 0.05309f
C5 CKN BULKP -0.227092f
C6 BULKP AVDD -3.515122f
C7 MP0/S CI -0.056784f
C8 MP0/S AVSS 0.208328f
C9 MP6_DMY/a_216_334# BULKN 0.091338f
C10 AVDD BULKN 0.74157f
C11 BULKP BULKN 7.544365f
C12 CK BULKN 0.372036f
C13 MN6/a_324_334# BULKN 0.422f
C14 CI BULKN 1.791641f
C15 AVSS BULKN 0.555322f
C16 MN0/a_324_n18# BULKN 0.422415f
C17 MP0/S BULKN 0.370985f
C18 MP0/a_216_n18# BULKN 0.091338f
C19 CKN BULKN 0.56349f
.ends

.subckt SUNSAR_SARCMPHX1_CV CI CK VMR N2 AVDD AVSS MP6/a_216_334# MN6/a_324_334# BULKP
+ MP0/a_216_n18# CO BULKN MN0/a_324_n18# N1
XMP0 AVDD CK N1 BULKP BULKN MP0/a_216_n18# CK SUNSAR_PCHDL
XMP1 N2 CK AVDD BULKP BULKN CK AVDD SUNSAR_PCHDL
XMN0 N1 CK AVSS BULKN MN0/a_324_n18# CI SUNSAR_NCHDL
XMP2 AVDD AVDD N2 BULKP BULKN CK CK SUNSAR_PCHDL
XMN1 N2 CI N1 BULKN CK CI SUNSAR_NCHDL
XMP3 CO CK AVDD BULKP BULKN AVDD VMR SUNSAR_PCHDL
XMP4 AVDD VMR CO BULKP BULKN CK VMR SUNSAR_PCHDL
XMN2 N1 CI N2 BULKN CI CI SUNSAR_NCHDL
XMP5 CO VMR AVDD BULKP BULKN VMR VMR SUNSAR_PCHDL
XMN3 N2 CI N1 BULKN CI CI SUNSAR_NCHDL
XMN4 N1 CI N2 BULKN CI CI SUNSAR_NCHDL
XMP6 AVDD VMR CO BULKP BULKN VMR MP6/a_216_334# SUNSAR_PCHDL
XMN5 N2 CI N1 BULKN CI VMR SUNSAR_NCHDL
XMN6 CO VMR N2 BULKN CI MN6/a_324_334# SUNSAR_NCHDL
C0 N1 AVDD 0.059184f
C1 BULKP CK -1.349649f
C2 BULKP CO 0.063159f
C3 N1 CI 0.175052f
C4 N2 CO 0.076147f
C5 N2 BULKP 0.063625f
C6 N2 AVSS 0.095751f
C7 CO VMR 0.076819f
C8 BULKP VMR -1.552184f
C9 AVDD CK 0.06305f
C10 AVDD CO 0.222193f
C11 AVDD BULKP -0.442314f
C12 AVDD AVSS 0.157463f
C13 N1 CK 0.072917f
C14 N1 BULKP 0.069686f
C15 N1 AVSS 0.158948f
C16 AVDD N2 0.080721f
C17 CI AVSS 0.057076f
C18 N1 N2 0.189549f
C19 AVDD VMR 0.050722f
C20 AVSS BULKN 0.533831f
C21 MN6/a_324_334# BULKN 0.422f
C22 VMR BULKN 0.606867f
C23 MP6/a_216_334# BULKN 0.091338f
C24 CI BULKN 1.771056f
C25 CK BULKN 0.626869f
C26 CO BULKN 0.213838f
C27 BULKP BULKN 7.544966f
C28 N2 BULKN 0.221339f
C29 MN0/a_324_n18# BULKN 0.422415f
C30 AVDD BULKN 0.609607f
C31 N1 BULKN 0.369132f
C32 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_IVX4_CV AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18#
+ Y BULKN A MN0/a_324_n18#
XMP0 Y A AVDD BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 AVDD A Y BULKP BULKN A A SUNSAR_PCHDL
XMP2 Y A AVDD BULKP BULKN A A SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 AVDD A Y BULKP BULKN A MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS A Y BULKN A A SUNSAR_NCHDL
XMN2 Y A AVSS BULKN A A SUNSAR_NCHDL
XMN3 AVSS A Y BULKN A MN3/a_324_334# SUNSAR_NCHDL
C0 Y A 0.147008f
C1 AVDD A 0.064966f
C2 BULKP AVDD 0.166303f
C3 Y AVSS 0.174863f
C4 BULKP A -1.606473f
C5 AVDD AVSS 0.131604f
C6 AVSS A 0.064848f
C7 AVDD Y 0.146264f
C8 A BULKN 2.062361f
C9 AVSS BULKN 0.622587f
C10 MN3/a_324_334# BULKN 0.422f
C11 MP3/a_216_334# BULKN 0.091338f
C12 Y BULKN 0.278637f
C13 MN0/a_324_n18# BULKN 0.422415f
C14 AVDD BULKN 0.372455f
C15 BULKP BULKN 5.176431f
C16 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARCMPX1_CV CPI CNI CK_CMP XA3a/A CK_SAMPLE DONE XA9/A CPO XA4/MP0/S
+ AVDD CNO AVSS
XXA10 XA9/A AVDD AVSS XA11/MN0/a_324_n18# XA12/Y XA11/Y AVDD AVSS XA9/MP0/a_216_334#
+ XA10/MN1/S XA11/MP0/a_216_n18# XA9/MN0/a_324_334# SUNSAR_NDX1_CV
XXA11 AVDD AVSS XA12/MN0/a_324_n18# DONE AVDD AVSS XA11/MP0/a_216_n18# XA11/Y XA12/MP0/a_216_n18#
+ CK_SAMPLE XA11/MN0/a_324_n18# SUNSAR_NRX1_CV
XXA12 AVDD AVSS XA12/Y AVSS XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD CK_CMP XA12/MN0/a_324_n18#
+ XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVDD XA13/MN1/a_324_n18# XA13/MN1/a_324_334# AVSS XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# AVSS XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA1 CPI AVDD AVDD AVSS XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# XA1/MP0/S XA9/A XA1/MP0/a_216_n18#
+ XA9/Y AVSS XA1/MN0/a_324_n18# SUNSAR_SARKICKHX1_CV
XXA2 CPI XA9/Y XA3/CO XA2/N2 AVDD AVSS XA2/MP6/a_216_334# XA2/MN6/a_324_334# AVDD
+ XA2/MP0/a_216_n18# XA3a/A AVSS XA2/MN0/a_324_n18# XA3/N1 SUNSAR_SARCMPHX1_CV
XXA3 CNI XA9/Y XA3a/A XA3/N2 AVDD AVSS XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVDD
+ XA3/MP0/a_216_n18# XA3/CO AVSS XA3/MN0/a_324_n18# XA3/N1 SUNSAR_SARCMPHX1_CV
XXA4 CNI AVDD AVDD AVSS XA9/MP0/a_216_n18# XA9/MN0/a_324_n18# XA4/MP0/S XA9/A XA4/MP0/a_216_n18#
+ XA9/Y AVSS XA4/MN0/a_324_n18# SUNSAR_SARKICKHX1_CV
XXA3a AVDD AVSS XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVDD XA3a/MP0/a_216_n18# CNO
+ AVSS XA3a/A XA3a/MN0/a_324_n18# SUNSAR_IVX4_CV
XXA2a AVDD AVSS XA3a/MP0/a_216_n18# XA3a/MN0/a_324_n18# AVDD XA2/MP6/a_216_334# CPO
+ AVSS XA3/CO XA2/MN6/a_324_334# SUNSAR_IVX4_CV
XXA9 AVDD AVSS XA9/Y AVSS XA9/MP0/a_216_n18# XA9/MP0/a_216_334# AVDD XA9/A XA9/MN0/a_324_n18#
+ XA9/MN0/a_324_334# SUNSAR_IVX1_CV
C0 XA9/Y AVDD 0.164728f
C1 XA13/MP1/a_216_n18# AVDD -0.311986f
C2 XA3/CO XA9/A 0.141462f
C3 XA12/Y CK_CMP 0.05138f
C4 XA3a/MP0/a_216_n18# AVDD -0.312264f
C5 AVDD XA4/MP0/a_216_n18# -0.311987f
C6 AVDD XA2/MP6/a_216_334# -0.313518f
C7 XA9/MP0/a_216_334# AVDD -0.311309f
C8 XA3/CO XA3/N1 0.289212f
C9 XA11/MP0/a_216_n18# AVDD -0.312939f
C10 XA3/CO AVDD 1.166637f
C11 XA3/N1 CNO 0.113873f
C12 DONE CK_CMP 0.058881f
C13 XA3a/A CPO 0.108133f
C14 XA3a/A XA9/Y 0.391167f
C15 XA1/MP0/S AVDD 0.073122f
C16 CNI XA9/Y 0.382485f
C17 XA1/MP0/a_216_n18# AVDD -0.311986f
C18 XA9/MP0/a_216_n18# AVDD -0.311986f
C19 XA3a/A XA3/CO 1.092423f
C20 XA9/A AVDD 0.189383f
C21 XA9/Y CPI 0.27081f
C22 XA12/Y CK_SAMPLE 0.106092f
C23 XA3/N1 AVDD 0.195531f
C24 XA2/MP0/a_216_n18# AVDD -0.311986f
C25 XA11/Y CK_SAMPLE 0.050093f
C26 XA11/Y XA12/Y 0.130476f
C27 XA3a/A XA9/A 0.136678f
C28 CNI XA9/A 0.362147f
C29 XA3a/A XA3/N1 0.309118f
C30 XA3a/A AVDD 0.912932f
C31 XA3/CO XA4/MP0/S 0.095491f
C32 XA9/A CPI 0.297822f
C33 XA3/CO XA9/Y 0.24121f
C34 XA12/MP0/a_216_n18# AVDD -0.312799f
C35 XA3/N1 CPI 0.115376f
C36 XA11/Y XA9/A 0.268591f
C37 AVDD XA3/MP0/a_216_n18# -0.313369f
C38 XA9/A XA9/Y 1.524979f
C39 XA12/Y AVDD 0.490048f
C40 XA3/N1 CPO 0.068565f
C41 XA3/N1 XA9/Y 0.106124f
C42 XA11/Y AVDD 0.055244f
C43 XA9/MN0/a_324_n18# AVSS 0.355152f
C44 XA3/CO AVSS 2.700073f
C45 CPO AVSS 0.178234f
C46 XA2/MN6/a_324_334# AVSS 0.353692f
C47 XA3a/A AVSS 2.521704f
C48 XA3/MN0/a_324_n18# AVSS 0.353692f
C49 CNO AVSS 0.179699f
C50 XA3a/MN0/a_324_n18# AVSS 0.353692f
C51 XA4/MN0/a_324_n18# AVSS 0.3537f
C52 XA4/MP0/S AVSS 0.414246f
C53 CNI AVSS 3.621781f
C54 XA3/N2 AVSS 0.246915f
C55 XA9/Y AVSS 4.611301f
C56 XA2/N2 AVSS 0.246915f
C57 XA2/MN0/a_324_n18# AVSS 0.353761f
C58 XA3/N1 AVSS 1.207811f
C59 AVDD AVSS 46.225956f
C60 CPI AVSS 3.746344f
C61 XA1/MN0/a_324_n18# AVSS 0.356268f
C62 XA1/MP0/S AVSS 0.422681f
C63 XA9/A AVSS 4.708538f
C64 XA0/MN1/a_324_n18# AVSS 0.422415f
C65 XA0/MP1/a_216_n18# AVSS 0.091271f
C66 XA13/MN1/a_324_n18# AVSS 0.356268f
C67 XA13/MN1/a_324_334# AVSS 0.422f
C68 XA13/MP1/a_216_334# AVSS 0.091271f
C69 CK_CMP AVSS 0.538462f
C70 XA12/MN0/a_324_n18# AVSS 0.356976f
C71 XA11/MN0/a_324_n18# AVSS 0.354241f
C72 DONE AVSS 0.474555f
C73 CK_SAMPLE AVSS 0.470196f
C74 XA9/MN0/a_324_334# AVSS 0.355744f
C75 XA12/Y AVSS 0.688419f
C76 XA11/Y AVSS 0.835235f
.ends

.subckt SUNSAR_NCHDLR D G S B a_324_n18# a_324_334#
X0 D G S B sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 D S 0.050207f
C1 a_324_n18# G 0.066018f
C2 a_324_334# G 0.067588f
C3 S B 0.06638f
C4 G B 0.415197f
C5 D B 0.06638f
C6 a_324_n18# B 0.422415f
C7 a_324_334# B 0.422f
.ends

.subckt SUNSAR_CAP_BSSW_CV A B 0
R0 A m3_6948_120# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R1 m3_252_280# B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
C0 A B 65.019196f
C1 m3_6948_120# B 0.172147f
C2 m3_6876_120# B 0.0666f
C3 m3_324_280# A 0.0666f
C4 m3_252_280# A 0.105547f
C5 B 0 13.2906f
C6 A 0 13.2887f
.ends

.subckt SUNSAR_CAP_BSSW5_CV B 0 A
XXCAPB0 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB1 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB2 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB3 A B 0 SUNSAR_CAP_BSSW_CV
XXCAPB4 A B 0 SUNSAR_CAP_BSSW_CV
C0 A B 54.004265f
C1 B 0 54.06679f
C2 A 0 55.079098f
.ends

.subckt SUNSAR_TIEH_CV Y BULKP AVDD AVSS MP0/G BULKN MP0/a_216_n18# MP0/a_216_334#
+ MN0/a_324_n18# MN0/a_324_334#
XMP0 Y MP0/G AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 MP0/G MP0/G AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.106173f
C1 BULKP MP0/G 0.112786f
C2 AVSS AVDD 0.051104f
C3 MP0/G AVSS 0.057963f
C4 AVDD BULKN 0.24902f
C5 AVSS BULKN 0.367715f
C6 MP0/G BULKN 0.790179f
C7 MN0/a_324_n18# BULKN 0.422415f
C8 MN0/a_324_334# BULKN 0.422f
C9 BULKP BULKN 2.806854f
C10 MP0/a_216_n18# BULKN 0.091338f
C11 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TIEL_CV BULKP AVDD AVSS MP0/G Y BULKN MP0/a_216_n18# MP0/a_216_334#
+ MN0/a_324_n18# MN0/a_324_334#
XMP0 MP0/G MP0/G AVDD BULKP BULKN MP0/a_216_n18# MP0/a_216_334# SUNSAR_PCHDL
XMN0 Y MP0/G AVSS BULKN MN0/a_324_n18# MN0/a_324_334# SUNSAR_NCHDL
C0 BULKP AVDD 0.103703f
C1 BULKP MP0/G 0.161174f
C2 AVSS AVDD 0.051104f
C3 MP0/G AVDD 0.057965f
C4 AVDD BULKN 0.249049f
C5 AVSS BULKN 0.370369f
C6 MP0/G BULKN 0.708387f
C7 Y BULKN 0.05974f
C8 MN0/a_324_n18# BULKN 0.422415f
C9 MN0/a_324_334# BULKN 0.422f
C10 BULKP BULKN 2.806659f
C11 MP0/a_216_n18# BULKN 0.091338f
C12 MP0/a_216_334# BULKN 0.091338f
.ends

.subckt SUNSAR_TGPD_CV AVSS MP2/B MN2/a_324_334# MP0/S B MP0/a_216_n18# A 0 C MP2/a_216_334#
+ MN0/a_324_n18# AVDD
XMP1_DMY B AVDD AVDD MP2/B 0 C C SUNSAR_PCHDL
XMP0 AVDD C MP0/S MP2/B 0 MP0/a_216_n18# AVDD SUNSAR_PCHDL
XMN0 AVSS C MP0/S 0 MN0/a_324_n18# C SUNSAR_NCHDL
XMP2 A C B MP2/B 0 AVDD MP2/a_216_334# SUNSAR_PCHDL
XMN1 B C AVSS 0 C MP0/S SUNSAR_NCHDL
XMN2 A MP0/S B 0 C MN2/a_324_334# SUNSAR_NCHDL
C0 C MP2/B -0.388363f
C1 B MP0/S 0.056087f
C2 C MP0/S 0.148714f
C3 MP2/B AVDD -0.506518f
C4 MP0/S AVSS 0.094973f
C5 C AVDD 0.07024f
C6 AVSS AVDD 0.090372f
C7 B A 0.108f
C8 MP0/S MP2/B 0.064367f
C9 AVDD 0 0.478784f
C10 AVSS 0 0.352742f
C11 A 0 0.204323f
C12 MN2/a_324_334# 0 0.422f
C13 MP2/B 0 4.387254f
C14 MP2/a_216_334# 0 0.091338f
C15 MP0/S 0 0.747699f
C16 MN0/a_324_n18# 0 0.422415f
C17 MP0/a_216_n18# 0 0.091338f
C18 B 0 0.060014f
C19 C 0 0.995573f
.ends

.subckt SUNSAR_SARBSSWCTRL_CV GN GNG TIE_H BULKP AVDD AVSS MN1/a_324_334# C BULKN
+ MP0/a_216_n18# MP1/a_216_334# MN0/a_324_n18#
XMP0 GNG C GN BULKP BULKN MP0/a_216_n18# GN SUNSAR_PCHDL
XMP1 AVDD GN GNG BULKP BULKN C MP1/a_216_334# SUNSAR_PCHDL
XMN0 MN1/S C AVSS BULKN MN0/a_324_n18# TIE_H SUNSAR_NCHDL
XMN1 GN TIE_H MN1/S BULKN C MN1/a_324_334# SUNSAR_NCHDL
C0 BULKP GN -0.16538f
C1 BULKP C -0.234337f
C2 AVSS AVDD 0.059137f
C3 BULKP GNG -0.056171f
C4 GN AVDD 0.071443f
C5 GN AVSS 0.082479f
C6 C GN 0.105655f
C7 BULKP AVDD 0.119037f
C8 AVDD BULKN 0.263047f
C9 AVSS BULKN 0.384798f
C10 TIE_H BULKN 0.37082f
C11 GN BULKN 0.410388f
C12 MN1/a_324_334# BULKN 0.422f
C13 C BULKN 0.568156f
C14 MN0/a_324_n18# BULKN 0.422415f
C15 MP1/a_216_334# BULKN 0.091338f
C16 BULKP BULKN 3.595271f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARBSSW_CV VI CK TIE_L VO1 M4/G VO2 XA3/B CKN XA4/GNG AVDD AVSS
XM1 VI M4/G VO1 AVSS M1/a_324_n18# M2/a_324_n18# SUNSAR_NCHDLR
XM2 VI M4/G VO1 AVSS M2/a_324_n18# M3/a_324_n18# SUNSAR_NCHDLR
XM3 VI M4/G VO1 AVSS M3/a_324_n18# M4/a_324_n18# SUNSAR_NCHDLR
XM4 VI M4/G VO1 AVSS M4/a_324_n18# M5/a_324_n18# SUNSAR_NCHDLR
XM5 VI TIE_L VO2 AVSS M5/a_324_n18# M6/a_324_n18# SUNSAR_NCHDLR
XXCAPB1 XA3/B AVSS XA4/GNG SUNSAR_CAP_BSSW5_CV
XM6 VI TIE_L VO2 AVSS M6/a_324_n18# M7/a_324_n18# SUNSAR_NCHDLR
XM7 VI TIE_L VO2 AVSS M7/a_324_n18# M8/a_324_n18# SUNSAR_NCHDLR
XM8 VI TIE_L VO2 AVSS M8/a_324_n18# M8/a_324_334# SUNSAR_NCHDLR
XXA0 AVDD AVSS CKN AVSS XA0/MP0/a_216_n18# XA3/MP0/a_216_n18# AVDD CK XA0/MN0/a_324_n18#
+ XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA1 XA1/Y AVDD AVDD AVSS XA1/MP0/G AVSS XA4/MP1/a_216_334# XA7/MP1/a_216_n18# XA4/MN1/a_324_334#
+ XA7/MN1/a_324_n18# SUNSAR_TIEH_CV
XXA2 AVDD AVDD AVSS XA2/MP0/G TIE_L AVSS XA7/MP1/a_216_334# XA5/MP1/a_216_n18# XA7/MN1/a_324_334#
+ XA5/MN1/a_324_n18# SUNSAR_TIEL_CV
XXA3 AVSS AVDD XA4/MN0/a_324_n18# XA3/MP0/S XA3/B XA3/MP0/a_216_n18# VI AVSS CKN XA4/MP0/a_216_n18#
+ XA3/MN0/a_324_n18# AVDD SUNSAR_TGPD_CV
XXA5 AVDD XA5/MN1/a_324_n18# XA5/MN1/a_324_334# AVSS XA5/MP1/a_216_334# XA5/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA4 M4/G XA4/GNG XA1/Y AVDD AVDD AVSS XA4/MN1/a_324_334# CKN AVSS XA4/MP0/a_216_n18#
+ XA4/MP1/a_216_334# XA4/MN0/a_324_n18# SUNSAR_SARBSSWCTRL_CV
XXA5b AVDD XA5b/MN1/a_324_n18# XA0/MN0/a_324_n18# AVSS XA0/MP0/a_216_n18# XA5b/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA7 AVDD XA7/MN1/a_324_n18# XA7/MN1/a_324_334# AVSS XA7/MP1/a_216_334# XA7/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
C0 CK CKN 0.081692f
C1 AVDD AVSS 0.15268f
C2 AVDD XA1/Y 0.335195f
C3 TIE_L VO2 0.067503f
C4 XA1/MP0/G AVSS 0.086644f
C5 XA1/MP0/G XA1/Y 0.210055f
C6 M4/G XA4/GNG 0.159364f
C7 AVDD XA3/MP0/a_216_n18# -0.315912f
C8 AVSS CKN 0.456081f
C9 VO2 AVSS 0.115254f
C10 TIE_L AVSS 0.570893f
C11 XA1/Y CKN 0.083971f
C12 XA2/MP0/G AVDD 0.154505f
C13 M4/G CKN 0.164954f
C14 VI CKN 0.158203f
C15 VI VO2 0.402032f
C16 VI TIE_L 0.431895f
C17 XA4/MP0/a_216_n18# AVDD -0.315004f
C18 XA3/MP0/S CKN 0.35416f
C19 XA7/MP1/a_216_n18# AVDD -0.314016f
C20 XA3/B AVDD 1.133969f
C21 XA5/MP1/a_216_n18# AVDD -0.311986f
C22 XA4/GNG AVDD 2.405915f
C23 AVDD CKN 0.381615f
C24 VO1 AVSS 0.112136f
C25 XA1/Y AVSS 0.269286f
C26 M4/G AVSS 0.641192f
C27 VI AVSS 0.44414f
C28 XA4/MP1/a_216_334# AVDD -0.310882f
C29 M4/G VO1 0.121857f
C30 M4/G XA1/Y 0.191529f
C31 TIE_L XA2/MP0/G 0.062843f
C32 XA4/GNG XA3/B 0.074834f
C33 VI VO1 0.509495f
C34 VI M4/G 0.733023f
C35 XA7/MP1/a_216_334# AVDD -0.311812f
C36 XA0/MP0/a_216_n18# AVDD -0.310529f
C37 XA3/B CKN 0.220083f
C38 VI XA3/MP0/S 0.083601f
C39 XA4/GNG CKN 0.13356f
C40 XA7/MN1/a_324_n18# 0 0.359583f
C41 AVSS 0 2.93973f
C42 XA5b/MN1/a_324_n18# 0 0.422415f
C43 AVDD 0 16.012844f
C44 XA5b/MP1/a_216_n18# 0 0.091271f
C45 XA1/Y 0 0.690197f
C46 CKN 0 1.768971f
C47 XA4/MN0/a_324_n18# 0 0.359583f
C48 XA5/MN1/a_324_334# 0 0.422f
C49 XA5/MP1/a_216_334# 0 0.091271f
C50 XA3/MP0/S 0 0.743486f
C51 XA3/MN0/a_324_n18# 0 0.359583f
C52 XA2/MP0/G 0 0.708335f
C53 XA7/MN1/a_324_334# 0 0.359583f
C54 XA5/MN1/a_324_n18# 0 0.360407f
C55 XA1/MP0/G 0 0.788614f
C56 XA4/MN1/a_324_334# 0 0.359583f
C57 CK 0 0.513823f
C58 XA0/MN0/a_324_n18# 0 0.359583f
C59 M8/a_324_n18# 0 0.356977f
C60 M8/a_324_334# 0 0.422f
C61 M6/a_324_n18# 0 0.356977f
C62 M7/a_324_n18# 0 0.356977f
C63 XA3/B 0 54.41209f
C64 XA4/GNG 0 53.065117f
C65 VO2 0 0.317444f
C66 TIE_L 0 2.408263f
C67 M5/a_324_n18# 0 0.356977f
C68 M3/a_324_n18# 0 0.356977f
C69 M4/a_324_n18# 0 0.356977f
C70 VO1 0 0.370636f
C71 M4/G 0 2.475647f
C72 VI 0 1.254522f
C73 M1/a_324_n18# 0 0.422415f
C74 M2/a_324_n18# 0 0.356977f
.ends

.subckt SUNSAR_SAREMX1_CV B EN ENO AVDD MP3/a_216_334# MN3/a_324_334# MP3/G A MN2/S
+ BULKP MP0/a_216_n18# AVSS BULKN RST_N MN0/a_324_n18#
XMP0 AVDD RST_N MP3/G BULKP BULKN MP0/a_216_n18# MP1/a_216_n18# SUNSAR_PCHDL
XMP1 MP2/S B ENO BULKP BULKN MP1/a_216_n18# MP2/a_216_n18# SUNSAR_PCHDL
XMP2 MP3/S A MP2/S BULKP BULKN MP2/a_216_n18# MP3/a_216_n18# SUNSAR_PCHDL
XMN0 MN2/S EN MP3/G BULKN MN0/a_324_n18# MN1/a_324_n18# SUNSAR_NCHDL
XMP3 AVDD MP3/G MP3/S BULKP BULKN MP3/a_216_n18# MP3/a_216_334# SUNSAR_PCHDL
XMN1 MN2/S B AVSS BULKN MN1/a_324_n18# MN2/a_324_n18# SUNSAR_NCHDL
XMN2 AVSS A MN2/S BULKN MN2/a_324_n18# MN3/a_324_n18# SUNSAR_NCHDL
XMN3 ENO MP3/G AVSS BULKN MN3/a_324_n18# MN3/a_324_334# SUNSAR_NCHDL
C0 MP3/S AVDD 0.067256f
C1 MP2/S ENO 0.064105f
C2 B A 0.058881f
C3 BULKP MP2/a_216_n18# -0.311038f
C4 ENO AVDD 0.155663f
C5 ENO AVSS 0.064883f
C6 MP2/S AVDD 0.054398f
C7 BULKP ENO 0.182005f
C8 BULKP MP1/a_216_n18# -0.311038f
C9 AVSS AVDD 0.157524f
C10 MP3/G A 0.105132f
C11 BULKP AVDD 0.233317f
C12 BULKP AVSS 0.058487f
C13 BULKP A 0.108551f
C14 MP3/S MP3/G 0.063428f
C15 BULKP B 0.113772f
C16 ENO MP3/G 0.133485f
C17 MP2/S MP3/G 0.064105f
C18 MP3/G AVDD 0.124994f
C19 ENO MP3/S 0.064105f
C20 MP3/G AVSS 0.050803f
C21 BULKP MP3/a_216_n18# -0.311038f
C22 RST_N MP3/G 0.054556f
C23 MN2/S AVSS 0.206972f
C24 BULKP MP3/G 0.480172f
C25 AVDD BULKN 0.390025f
C26 AVSS BULKN 0.695296f
C27 MN3/a_324_n18# BULKN 0.35253f
C28 MN3/a_324_334# BULKN 0.422f
C29 A BULKN 0.498033f
C30 MN2/a_324_n18# BULKN 0.352522f
C31 B BULKN 0.513991f
C32 MN1/a_324_n18# BULKN 0.352522f
C33 MP3/a_216_334# BULKN 0.091338f
C34 MP3/G BULKN 0.827536f
C35 EN BULKN 0.386445f
C36 MN2/S BULKN 0.207484f
C37 MN0/a_324_n18# BULKN 0.422415f
C38 ENO BULKN 0.246284f
C39 BULKP BULKN 7.539519f
C40 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARLTX1_CV RST_N EN LCK_N AVDD AVSS MN2/a_324_334# A BULKP MP0/a_216_n18#
+ CHL BULKN MP2/a_216_334# MN0/a_324_n18#
XMP0 MP1/S RST_N AVDD BULKP BULKN MP0/a_216_n18# RST_N SUNSAR_PCHDL
XMP1 MP2/S RST_N MP1/S BULKP BULKN RST_N RST_N SUNSAR_PCHDL
XMN0 MN1/S A AVSS BULKN MN0/a_324_n18# LCK_N SUNSAR_NCHDL
XMP2 CHL RST_N MP2/S BULKP BULKN RST_N MP2/a_216_334# SUNSAR_PCHDL
XMN1 MN2/S LCK_N MN1/S BULKN A EN SUNSAR_NCHDL
XMN2 CHL EN MN2/S BULKN LCK_N MN2/a_324_334# SUNSAR_NCHDL
C0 BULKP MP2/S -0.050867f
C1 BULKP RST_N -1.319845f
C2 BULKP CHL 0.074842f
C3 AVDD AVSS 0.088964f
C4 AVDD BULKP 0.143379f
C5 MP1/S BULKP -0.050867f
C6 EN BULKN 0.372036f
C7 MN2/a_324_334# BULKN 0.422f
C8 LCK_N BULKN 0.335836f
C9 AVSS BULKN 0.428199f
C10 RST_N BULKN 0.123012f
C11 CHL BULKN 0.260933f
C12 BULKP BULKN 4.387078f
C13 MP2/a_216_334# BULKN 0.091338f
C14 A BULKN 0.372036f
C15 MN0/a_324_n18# BULKN 0.422415f
C16 AVDD BULKN 0.276832f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARMRYX1_CV CMP_OP CHL_OP CHL_ON XA1/MP3/G RST_N XA5/MP2/a_216_334#
+ ENO XA5/MN2/a_324_334# XA1/MN2/S CMP_ON AVDD AVSS XA2/Y EN
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# AVSS XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA1 CMP_ON EN ENO AVDD XA2/MP0/a_216_n18# XA2/MN0/a_324_n18# XA1/MP3/G CMP_OP XA1/MN2/S
+ AVDD XA1/MP0/a_216_n18# AVSS AVSS RST_N XA1/MN0/a_324_n18# SUNSAR_SAREMX1_CV
XXA2 AVDD AVSS XA2/Y AVSS XA2/MP0/a_216_n18# XA4/MP0/a_216_n18# AVDD ENO XA2/MN0/a_324_n18#
+ XA4/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA4 RST_N EN XA2/Y AVDD AVSS XA5/MN0/a_324_n18# CMP_OP AVDD XA4/MP0/a_216_n18# CHL_OP
+ AVSS XA5/MP0/a_216_n18# XA4/MN0/a_324_n18# SUNSAR_SARLTX1_CV
XXA5 RST_N EN XA2/Y AVDD AVSS XA5/MN2/a_324_334# CMP_ON AVDD XA5/MP0/a_216_n18# CHL_ON
+ AVSS XA5/MP2/a_216_334# XA5/MN0/a_324_n18# SUNSAR_SARLTX1_CV
C0 ENO XA2/Y 0.081815f
C1 ENO CMP_OP 0.15365f
C2 XA2/MP0/a_216_n18# AVDD -0.31403f
C3 XA1/MP0/a_216_n18# AVDD -0.311986f
C4 AVDD RST_N 1.195814f
C5 AVDD XA2/Y 0.086382f
C6 ENO XA1/MP3/G 0.074928f
C7 CMP_OP XA2/Y 0.183507f
C8 AVDD XA4/MP0/a_216_n18# -0.31403f
C9 CMP_ON XA2/Y 0.130187f
C10 CMP_ON CMP_OP 0.054599f
C11 XA1/MP3/G RST_N 0.080501f
C12 EN XA2/Y 0.114038f
C13 EN CMP_OP 0.196887f
C14 AVDD CHL_OP 0.069236f
C15 AVDD XA5/MP0/a_216_n18# -0.31403f
C16 EN CMP_ON 0.54292f
C17 XA5/MN2/a_324_334# AVSS 0.422f
C18 CHL_ON AVSS 0.232377f
C19 XA5/MP2/a_216_334# AVSS 0.091271f
C20 XA5/MN0/a_324_n18# AVSS 0.3537f
C21 RST_N AVSS 0.223373f
C22 CHL_OP AVSS 0.170032f
C23 XA4/MN0/a_324_n18# AVSS 0.3537f
C24 XA2/Y AVSS 1.191276f
C25 XA2/MN0/a_324_n18# AVSS 0.353715f
C26 XA1/MN3/a_324_n18# AVSS 0.352733f
C27 CMP_OP AVSS 1.302224f
C28 XA1/MN2/a_324_n18# AVSS 0.353381f
C29 CMP_ON AVSS 1.822119f
C30 XA1/MN1/a_324_n18# AVSS 0.358f
C31 XA1/MP3/G AVSS 0.885586f
C32 EN AVSS 2.425524f
C33 XA1/MN2/S AVSS 0.199983f
C34 XA1/MN0/a_324_n18# AVSS 0.356268f
C35 ENO AVSS 0.8336f
C36 XA0/MN1/a_324_n18# AVSS 0.422415f
C37 AVDD AVSS 17.159056f
C38 XA0/MP1/a_216_n18# AVSS 0.091271f
.ends

.subckt SUNSAR_SWX4_CV MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18# Y BULKN
+ AVSS A MN0/a_324_n18# VREF
XMP0 Y A VREF BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 VREF A Y BULKP BULKN A A SUNSAR_PCHDL
XMP2 Y A VREF BULKP BULKN A A SUNSAR_PCHDL
XMN0 Y A AVSS BULKN MN0/a_324_n18# A SUNSAR_NCHDL
XMP3 VREF A Y BULKP BULKN A MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS A Y BULKN A A SUNSAR_NCHDL
XMN2 Y A AVSS BULKN A A SUNSAR_NCHDL
XMN3 AVSS A Y BULKN A MN3/a_324_334# SUNSAR_NCHDL
C0 BULKP A -1.606473f
C1 VREF AVSS 0.05784f
C2 A AVSS 0.076196f
C3 Y AVSS 0.180645f
C4 BULKP AVSS 0.062361f
C5 A VREF 0.184236f
C6 Y VREF 0.133073f
C7 Y A 0.147007f
C8 BULKP VREF 0.281929f
C9 AVSS BULKN 0.66508f
C10 MN3/a_324_334# BULKN 0.422f
C11 MP3/a_216_334# BULKN 0.091338f
C12 VREF BULKN 0.501044f
C13 A BULKN 2.06236f
C14 Y BULKN 0.278638f
C15 MN0/a_324_n18# BULKN 0.422415f
C16 BULKP BULKN 5.176431f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARCEX1_CV B Y RST AVDD AVSS MP3/a_216_334# MN3/a_324_334# BULKP MP0/a_216_n18#
+ BULKN A MN0/a_324_n18#
XMP0 MP1/S A Y BULKP BULKN MP0/a_216_n18# A SUNSAR_PCHDL
XMP1 AVDD A MP1/S BULKP BULKN A B SUNSAR_PCHDL
XMP2 MP3/S B AVDD BULKP BULKN A B SUNSAR_PCHDL
XMN0 MN1/S RST AVSS BULKN MN0/a_324_n18# RST SUNSAR_NCHDL
XMP3 Y B MP3/S BULKP BULKN B MP3/a_216_334# SUNSAR_PCHDL
XMN1 AVSS RST MN1/S BULKN RST RST SUNSAR_NCHDL
XMN2 MN3/S RST AVSS BULKN RST RST SUNSAR_NCHDL
XMN3 Y RST MN3/S BULKN RST MN3/a_324_334# SUNSAR_NCHDL
C0 AVSS Y 0.129646f
C1 BULKP B -1.00547f
C2 BULKP MP3/S -0.050867f
C3 RST Y 0.072094f
C4 BULKP AVDD 0.114602f
C5 BULKP A -1.005062f
C6 BULKP MP1/S -0.050867f
C7 MN1/S AVSS 0.058507f
C8 Y AVDD 0.07728f
C9 BULKP Y 0.191403f
C10 AVSS AVDD 0.106506f
C11 AVDD BULKN 0.247044f
C12 Y BULKN 0.484249f
C13 MN3/a_324_334# BULKN 0.422f
C14 AVSS BULKN 0.495556f
C15 MP3/a_216_334# BULKN 0.091338f
C16 RST BULKN 1.501372f
C17 MN0/a_324_n18# BULKN 0.422415f
C18 B BULKN 0.072331f
C19 A BULKN 0.072331f
C20 BULKP BULKN 5.174408f
C21 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_SARDIGEX4_CV CMP_OP CMP_ON CP0 CN1 XA1/XA2/Y XA9/B DONE XA1/XA1/MP3/G
+ CN0 RST_N XA11/A CEO CKS XA2/A ENO XA1/XA1/MN2/S XA4/A CP1 EN VREF CEIN XA12/A AVSS
+ AVDD
XXA10 AVDD AVSS XA11/A AVSS XA9/MP1/a_216_334# XA11/MP0/a_216_n18# AVDD XA9/Y XA9/MN1/a_324_334#
+ XA11/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA11 AVDD AVSS XA12/MN0/a_324_n18# CEIN AVDD AVSS XA11/MP0/a_216_n18# XA12/A XA12/MP0/a_216_n18#
+ XA11/A XA11/MN0/a_324_n18# SUNSAR_NRX1_CV
XXA12 AVDD AVSS CEO AVSS XA12/MP0/a_216_n18# XA13/MP1/a_216_n18# AVDD XA12/A XA12/MN0/a_324_n18#
+ XA13/MN1/a_324_n18# SUNSAR_IVX1_CV
XXA13 AVDD XA13/MN1/a_324_n18# XA13/MN1/a_324_334# AVSS XA13/MP1/a_216_334# XA13/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA1 CMP_OP XA4/A XA2/A XA1/XA1/MP3/G RST_N XA2/MP0/a_216_n18# ENO XA2/MN0/a_324_n18#
+ XA1/XA1/MN2/S CMP_ON AVDD AVSS XA1/XA2/Y EN SUNSAR_SARMRYX1_CV
XXA2 XA3/MP0/a_216_n18# XA3/MN0/a_324_n18# AVDD XA2/MP0/a_216_n18# CN1 AVSS AVSS XA2/A
+ XA2/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA3 XA4/MP0/a_216_n18# XA4/MN0/a_324_n18# AVDD XA3/MP0/a_216_n18# CP1 AVSS AVSS CN1
+ XA3/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA5 XA6/MP0/a_216_n18# XA6/MN0/a_324_n18# AVDD XA5/MP0/a_216_n18# CN0 AVSS AVSS CP0
+ XA5/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA4 XA5/MP0/a_216_n18# XA5/MN0/a_324_n18# AVDD XA4/MP0/a_216_n18# CP0 AVSS AVSS XA4/A
+ XA4/MN0/a_324_n18# VREF SUNSAR_SWX4_CV
XXA6 CP1 XA9/B CKS AVDD AVSS XA7/MP0/a_216_n18# XA7/MN0/a_324_n18# AVDD XA6/MP0/a_216_n18#
+ AVSS CN0 XA6/MN0/a_324_n18# SUNSAR_SARCEX1_CV
XXA7 AVDD AVSS XA9/A AVSS XA7/MP0/a_216_n18# XA8/MP0/a_216_n18# AVDD ENO XA7/MN0/a_324_n18#
+ XA8/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA8 AVDD AVSS DONE AVSS XA8/MP0/a_216_n18# XA9/MP0/a_216_n18# AVDD XA9/A XA8/MN0/a_324_n18#
+ XA9/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA9 XA9/Y AVDD AVSS XA9/MN1/a_324_334# XA9/B XA9/A AVDD AVSS XA9/MP0/a_216_n18# XA9/MN1/S
+ XA9/MP1/a_216_334# XA9/MN0/a_324_n18# SUNSAR_NDX1_CV
C0 AVDD XA5/MP0/a_216_n18# -0.298676f
C1 ENO XA2/A 0.090499f
C2 ENO XA9/B 0.051732f
C3 VREF CP1 1.096312f
C4 XA9/Y XA11/A 0.134948f
C5 AVDD VREF 2.204398f
C6 CN1 XA4/A 0.466806f
C7 ENO CMP_ON 0.067952f
C8 AVDD XA7/MP0/a_216_n18# -0.311987f
C9 XA12/A AVDD 0.092687f
C10 XA9/A XA9/B 0.245863f
C11 EN XA4/A 0.118846f
C12 CN0 CP0 0.298273f
C13 AVDD XA2/A 0.202922f
C14 AVDD XA9/B 0.076392f
C15 ENO CN1 0.083894f
C16 AVDD XA2/MP0/a_216_n18# -0.306139f
C17 AVDD XA9/MP1/a_216_334# -0.311908f
C18 ENO XA1/XA1/MP3/G 0.086456f
C19 CEO AVDD 0.06867f
C20 CN0 CP1 0.319562f
C21 AVDD CN0 0.409213f
C22 XA2/A VREF 0.115624f
C23 ENO XA4/A 0.119578f
C24 VREF XA9/B 0.062419f
C25 XA12/MP0/a_216_n18# AVDD -0.311309f
C26 CN1 CP1 0.208539f
C27 CP0 XA4/A 0.350838f
C28 AVDD CN1 0.114213f
C29 CN0 VREF 0.089412f
C30 AVDD XA8/MP0/a_216_n18# -0.311987f
C31 XA11/A AVDD 0.076411f
C32 CP1 XA4/A 0.193274f
C33 AVDD XA4/A 0.106262f
C34 CEIN XA12/A 0.110841f
C35 ENO CP0 0.08098f
C36 CN0 XA9/B 0.069404f
C37 AVDD XA6/MP0/a_216_n18# -0.306081f
C38 ENO XA9/A 0.07744f
C39 XA11/MP0/a_216_n18# AVDD -0.311842f
C40 XA9/A DONE 0.063409f
C41 XA13/MP1/a_216_n18# AVDD -0.311986f
C42 XA11/A XA12/A 0.07223f
C43 ENO CP1 0.402013f
C44 AVDD XA4/MP0/a_216_n18# -0.298676f
C45 AVDD ENO 2.495094f
C46 CN1 XA2/A 0.327387f
C47 AVDD DONE 0.055168f
C48 AVDD XA3/MP0/a_216_n18# -0.298153f
C49 CP1 CP0 0.176643f
C50 XA9/Y XA9/B 0.108031f
C51 XA1/XA2/Y XA4/A 0.161989f
C52 AVDD CP0 0.163708f
C53 XA2/A XA4/A 0.111482f
C54 ENO VREF 0.694105f
C55 AVDD XA9/A 0.068695f
C56 ENO RST_N 0.661116f
C57 AVDD XA9/MP0/a_216_n18# -0.311986f
C58 AVDD CP1 0.743971f
C59 XA9/MN1/a_324_334# AVSS 0.355152f
C60 XA9/MN0/a_324_n18# AVSS 0.3539f
C61 XA9/A AVSS 1.385168f
C62 DONE AVSS 0.144639f
C63 XA7/MN0/a_324_n18# AVSS 0.354718f
C64 XA8/MN0/a_324_n18# AVSS 0.355152f
C65 XA9/B AVSS 1.502327f
C66 CKS AVSS 1.45158f
C67 XA6/MN0/a_324_n18# AVSS 0.356268f
C68 XA4/A AVSS 3.131355f
C69 XA4/MN0/a_324_n18# AVSS 0.355744f
C70 CP0 AVSS 2.560386f
C71 CN0 AVSS 0.340136f
C72 XA5/MN0/a_324_n18# AVSS 0.355152f
C73 VREF AVSS 0.8336f
C74 CN1 AVSS 2.510553f
C75 CP1 AVSS 0.513004f
C76 XA3/MN0/a_324_n18# AVSS 0.355152f
C77 XA2/A AVSS 2.066712f
C78 XA2/MN0/a_324_n18# AVSS 0.355744f
C79 XA1/XA5/MN0/a_324_n18# AVSS 0.359841f
C80 RST_N AVSS 0.189551f
C81 XA1/XA4/MN0/a_324_n18# AVSS 0.360407f
C82 XA1/XA2/Y AVSS 1.04564f
C83 XA1/XA2/MN0/a_324_n18# AVSS 0.360407f
C84 XA1/XA1/MN3/a_324_n18# AVSS 0.355196f
C85 CMP_OP AVSS 1.158538f
C86 XA1/XA1/MN2/a_324_n18# AVSS 0.355196f
C87 CMP_ON AVSS 1.344542f
C88 XA1/XA1/MN1/a_324_n18# AVSS 0.355196f
C89 XA1/XA1/MP3/G AVSS 0.827195f
C90 EN AVSS 2.11207f
C91 XA1/XA1/MN2/S AVSS 0.200627f
C92 XA1/XA1/MN0/a_324_n18# AVSS 0.360407f
C93 ENO AVSS 1.875766f
C94 XA1/XA0/MN1/a_324_n18# AVSS 0.422415f
C95 AVDD AVSS 49.971783f
C96 XA1/XA0/MP1/a_216_n18# AVSS 0.091271f
C97 XA13/MN1/a_324_334# AVSS 0.422f
C98 XA13/MP1/a_216_334# AVSS 0.091271f
C99 CEO AVSS 0.198916f
C100 XA12/MN0/a_324_n18# AVSS 0.355467f
C101 XA13/MN1/a_324_n18# AVSS 0.356268f
C102 XA12/A AVSS 0.87316f
C103 XA11/MN0/a_324_n18# AVSS 0.355152f
C104 CEIN AVSS 0.470391f
C105 XA11/A AVSS 0.773693f
C106 XA9/Y AVSS 0.833f
.ends

.subckt SUNSAR_SAR8B_CV SAR_IP SAR_IN DONE D<7> D<4> D<1> EN XA3/CEO XA6/CN0 XA6/CP0
+ XA3/CN0 XA20/XA9/A XA3/CP0 XA4/DONE XA0/XA9/B XA7/CEO XA0/CP0 XA4/CEO XA7/CN0 D<0>
+ XA1/CEO XA7/CP0 XA4/CN0 D<3> XA0/CEIN XA4/CP0 XA1/CN0 D<6> XA2/DONE XA1/CP0 XA5/CEO
+ XA20/XA4/MP0/S CK_SAMPLE XA2/CEO SARP CK_SAMPLE_BSSW XA5/CN0 D<2> XA0/CEO XA5/CP0
+ XA6/DONE XA0/XA4/A XA2/CN0 D<5> VREF XA2/CP0 SARN AVDD XA6/CEO AVSS
XXDAC1 XA0/CP1 XA0/CP0 D<6> XA1/CP0 D<5> XA2/CP0 D<4> D<3> D<2> D<1> SARP AVSS AVSS
+ SUNSAR_CDAC7_CV
XXDAC2 D<7> XA0/CN0 XA1/CN1 XA1/CN0 XA2/CN1 XA2/CN0 XA3/CN0 XA4/CN0 XA5/CN0 XA6/CN0
+ SARN AVSS AVSS SUNSAR_CDAC7_CV
XXA20 SARP SARN XA7/CEO XA20/XA3a/A CK_SAMPLE DONE XA20/XA9/A XA20/CPO XA20/XA4/MP0/S
+ AVDD XA20/CNO AVSS SUNSAR_SARCMPX1_CV
XXB1 SAR_IP CK_SAMPLE_BSSW XA0/CEIN SARP XB1/M4/G SARN XB1/XA3/B XB1/CKN XB1/XA4/GNG
+ AVDD AVSS SUNSAR_SARBSSW_CV
XXA0 XA20/CPO XA20/CNO XA0/CP0 D<7> XA0/XA1/XA2/Y XA0/XA9/B XA0/DONE XA0/XA1/XA1/MP3/G
+ XA0/CN0 EN XA0/XA11/A XA0/CEO CK_SAMPLE XA0/XA2/A XA1/EN XA0/XA1/XA1/MN2/S XA0/XA4/A
+ XA0/CP1 EN VREF XA0/CEIN XA0/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXB2 SAR_IN CK_SAMPLE_BSSW XA0/CEIN SARN XB2/M4/G SARP XB2/XA3/B XB2/CKN XB2/XA4/GNG
+ AVDD AVSS SUNSAR_SARBSSW_CV
XXA1 XA20/CPO XA20/CNO XA1/CP0 XA1/CN1 XA1/XA1/XA2/Y XA1/XA9/B XA1/DONE XA1/XA1/XA1/MP3/G
+ XA1/CN0 EN XA1/XA11/A XA1/CEO CK_SAMPLE XA1/XA2/A XA2/EN XA1/XA1/XA1/MN2/S XA1/XA4/A
+ D<6> XA1/EN VREF XA0/CEO XA1/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA2 XA20/CPO XA20/CNO XA2/CP0 XA2/CN1 XA2/XA1/XA2/Y XA2/XA9/B XA2/DONE XA2/XA1/XA1/MP3/G
+ XA2/CN0 EN XA2/XA11/A XA2/CEO CK_SAMPLE XA2/XA2/A XA3/EN XA2/XA1/XA1/MN2/S XA2/XA4/A
+ D<5> XA2/EN VREF XA1/CEO XA2/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA3 XA20/CPO XA20/CNO XA3/CP0 XA3/CN1 XA3/XA1/XA2/Y XA3/XA9/B XA3/DONE XA3/XA1/XA1/MP3/G
+ XA3/CN0 EN XA3/XA11/A XA3/CEO CK_SAMPLE XA3/XA2/A XA4/EN XA3/XA1/XA1/MN2/S XA3/XA4/A
+ D<4> XA3/EN VREF XA2/CEO XA3/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA4 XA20/CPO XA20/CNO XA4/CP0 XA4/CN1 XA4/XA1/XA2/Y XA4/XA9/B XA4/DONE XA4/XA1/XA1/MP3/G
+ XA4/CN0 EN XA4/XA11/A XA4/CEO CK_SAMPLE XA4/XA2/A XA5/EN XA4/XA1/XA1/MN2/S XA4/XA4/A
+ D<3> XA4/EN VREF XA3/CEO XA4/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA5 XA20/CPO XA20/CNO XA5/CP0 XA5/CN1 XA5/XA1/XA2/Y XA5/XA9/B XA5/DONE XA5/XA1/XA1/MP3/G
+ XA5/CN0 EN XA5/XA11/A XA5/CEO CK_SAMPLE XA5/XA2/A XA6/EN XA5/XA1/XA1/MN2/S XA5/XA4/A
+ D<2> XA5/EN VREF XA4/CEO XA5/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA6 XA20/CPO XA20/CNO XA6/CP0 XA6/CN1 XA6/XA1/XA2/Y XA6/XA9/B XA6/DONE XA6/XA1/XA1/MP3/G
+ XA6/CN0 EN XA6/XA11/A XA6/CEO CK_SAMPLE XA6/XA2/A XA7/EN XA6/XA1/XA1/MN2/S XA6/XA4/A
+ D<1> XA6/EN VREF XA5/CEO XA6/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
XXA7 XA20/CPO XA20/CNO XA7/CP0 XA7/CN1 XA7/XA1/XA2/Y XA7/XA9/B DONE XA7/XA1/XA1/MP3/G
+ XA7/CN0 EN XA7/XA11/A XA7/CEO CK_SAMPLE XA7/XA2/A XA7/ENO XA7/XA1/XA1/MN2/S XA7/XA4/A
+ D<0> XA7/EN VREF XA6/CEO XA7/XA12/A AVSS AVDD SUNSAR_SARDIGEX4_CV
C0 XA5/CEO AVDD 0.342105f
C1 AVDD XA4/EN 0.11184f
C2 AVDD XA20/CNO 2.72258f
C3 D<4> XA1/CN0 0.070567f
C4 XA0/CP0 D<5> 0.306186f
C5 XA0/DONE AVSS 0.27339f
C6 XA20/CPO XA1/XA1/XA2/Y 0.078271f
C7 XA4/CN0 XA6/CN0 0.14269f
C8 XA7/XA12/A XA6/CEO 0.115411f
C9 VREF XA3/CN0 0.061066f
C10 XA2/CN0 XA1/CN0 2.065852f
C11 D<7> XA1/CP0 0.073351f
C12 XA1/CP0 XA0/CN0 0.398101f
C13 XA2/EN XA1/CN0 0.127391f
C14 XA0/CEIN XB2/CKN 0.100038f
C15 D<2> XA20/CNO 0.063406f
C16 XA7/CEO XA6/CEO 0.137785f
C17 XA6/EN AVSS 0.355405f
C18 D<7> XA0/CN0 0.494507f
C19 XA1/EN XA2/EN 1.263077f
C20 SARP SARN 5.1717f
C21 CK_SAMPLE XA0/XA9/B 0.07743f
C22 XA5/EN XA4/XA1/XA1/MP3/G 0.058161f
C23 XA4/CN0 AVSS 0.234489f
C24 XA5/DONE XA5/XA9/B 0.061581f
C25 XA20/CPO XA1/CP0 0.05767f
C26 AVSS XA7/CEO 0.539406f
C27 AVDD XA2/CEO 1.256112f
C28 CK_SAMPLE XA6/XA9/B 0.07743f
C29 XA20/CPO D<7> 0.239708f
C30 XA20/CPO XA0/CN0 0.06056f
C31 XA7/EN XA20/CPO 0.251284f
C32 XA1/CN1 XA1/CN0 0.608838f
C33 XA1/EN XA1/CN1 0.231611f
C34 D<7> XA3/CN0 0.073456f
C35 XA3/CN0 XA0/CN0 0.073103f
C36 CK_SAMPLE XA7/XA9/B 0.082731f
C37 D<6> XA1/CN0 0.099307f
C38 XA5/CN0 XA1/CN0 0.092052f
C39 XA1/EN D<6> 0.062843f
C40 D<4> XA2/CN1 0.098494f
C41 XA20/CPO XA3/CN0 0.068343f
C42 CK_SAMPLE XA3/XA9/B 0.078405f
C43 XA5/XA4/A XA6/XA4/A 0.082663f
C44 EN XA4/EN 0.235383f
C45 CK_SAMPLE D<5> 0.100705f
C46 XA20/CNO EN 2.032689f
C47 XA2/CN0 XA2/CN1 0.583006f
C48 XA20/CNO D<1> 0.063875f
C49 XA1/CN0 XA6/CN0 0.071338f
C50 XA2/EN XA2/CN1 0.336738f
C51 XA5/EN XA5/CN0 0.070138f
C52 XA0/CEIN SARP 0.431405f
C53 XA4/XA4/A XA3/XA4/A 0.082663f
C54 AVDD XA6/CP0 -0.052017f
C55 XA20/CNO XA2/CP0 0.054091f
C56 XA20/CNO XA1/XA4/A 0.286129f
C57 CK_SAMPLE XA3/EN 0.092446f
C58 XA1/CN0 AVSS 0.126506f
C59 VREF XA4/EN 0.175304f
C60 XA1/CN1 XA0/CP1 0.268769f
C61 AVDD XA2/CN0 2.508128f
C62 XA1/CN1 XA2/CN1 2.837019f
C63 XA0/XA4/A EN 0.080713f
C64 XA1/EN AVSS 0.167653f
C65 AVDD XA2/EN 0.11184f
C66 XA5/EN XA6/CN0 0.115359f
C67 D<6> XA0/CP1 1.561198f
C68 XA5/XA2/A EN 0.11418f
C69 D<6> XA2/CN1 0.199516f
C70 XA20/XA3a/A XA20/CNO 0.119511f
C71 XA5/CN0 XA2/CN1 0.073237f
C72 XA2/CEO XA3/XA12/A 0.084465f
C73 XA1/EN XA0/XA1/XA1/MP3/G 0.058161f
C74 D<2> XA2/CN0 0.077577f
C75 XA5/EN AVSS 0.218031f
C76 XA1/XA12/A XA1/CEO 0.264746f
C77 XA4/CEO XA5/XA12/A 0.084465f
C78 CK_SAMPLE D<0> 0.102094f
C79 XA7/EN XA7/XA1/XA1/MP3/G 0.096884f
C80 XB1/XA3/B AVDD 0.185337f
C81 VREF XA2/CEO 0.348781f
C82 XA20/CNO XA1/CP0 0.053078f
C83 CK_SAMPLE XA7/ENO 0.097331f
C84 XA2/CN1 XA6/CN0 0.077601f
C85 XA20/CNO D<7> 0.17726f
C86 XA20/CNO XA0/CN0 0.058198f
C87 XA5/CN0 AVDD 2.476604f
C88 XA7/EN XA20/CNO 0.39054f
C89 D<2> XA1/CN1 0.080525f
C90 XA20/XA9/A XA7/EN 0.291697f
C91 XA1/CEO AVSS 0.43736f
C92 XA20/CPO XA4/EN 0.378571f
C93 AVSS XA0/CP1 1.87901f
C94 XA4/CN1 XA4/CN0 0.051467f
C95 XA20/CNO XA20/CPO 6.984268f
C96 XA20/CNO XA2/XA4/A 0.212166f
C97 XA2/CN1 AVSS 1.031315f
C98 XA20/XA9/A XA20/CPO 0.365673f
C99 XA2/EN XA1/XA1/XA1/MN2/S 0.064012f
C100 XA5/DONE AVSS 0.267946f
C101 XA5/CN0 D<2> 1.58415f
C102 XA4/EN XA3/CN0 0.13801f
C103 EN D<4> 0.07107f
C104 AVDD XA6/CN0 2.589875f
C105 XA5/XA1/XA2/Y XA20/CPO 0.078271f
C106 XA0/XA4/A D<7> 0.06833f
C107 SARP XA0/CP0 0.107476f
C108 XA20/CNO XA3/CN0 0.064465f
C109 AVDD XA6/CEO 1.255434f
C110 EN XA2/CN0 0.066928f
C111 XA2/CN0 D<1> 0.075983f
C112 EN XA2/EN 0.235383f
C113 XA2/CP0 D<4> 0.835772f
C114 XA6/EN XA5/XA1/XA1/MN2/S 0.064012f
C115 AVDD AVSS 7.430067f
C116 D<2> XA6/CN0 0.155398f
C117 XB2/XA3/B AVSS 1.491395f
C118 XA1/CN0 D<5> 0.061568f
C119 XA2/CP0 XA2/CN0 3.180099f
C120 VREF D<4> 0.083402f
C121 XB1/M4/G SARN 0.156031f
C122 XB2/XA4/GNG AVSS 1.208553f
C123 XA20/XA3/N1 XA20/CPO 0.062971f
C124 D<2> AVSS 1.856228f
C125 EN XA1/CN1 0.09741f
C126 VREF XA2/CN0 0.061066f
C127 XA1/CN1 D<1> 0.070318f
C128 SAR_IP SARN 0.203945f
C129 VREF XA2/EN 0.175304f
C130 EN XA3/XA4/A 0.088236f
C131 EN D<6> 0.062969f
C132 XA2/CP0 XA1/CN1 0.065837f
C133 XA5/CN0 EN 0.073683f
C134 XA5/CN0 D<1> 0.07478f
C135 XA1/CN1 XA1/XA4/A 0.092747f
C136 D<4> XA1/CP0 0.174549f
C137 XA6/CN0 XA6/CN1 0.051467f
C138 D<7> D<4> 0.073464f
C139 D<4> XA0/CN0 0.077963f
C140 CK_SAMPLE XA1/XA9/B 0.078405f
C141 XA2/EN XA1/CP0 0.085659f
C142 XA3/CN1 XA3/CN0 0.051393f
C143 EN XA6/CN0 0.073805f
C144 XA6/CN0 D<1> 2.256405f
C145 VREF D<6> 0.083401f
C146 D<7> XA2/CN0 0.073503f
C147 XA2/CN0 XA0/CN0 0.07731f
C148 XA20/CPO D<4> 0.071873f
C149 XA5/CN0 VREF 0.061065f
C150 XB1/XA4/GNG XDAC1/XC1/XRES16/B 0.107427f
C151 XA2/CN1 D<5> 0.490947f
C152 XA0/CEIN XB1/M4/G 0.110451f
C153 XB1/XA4/GNG XDAC1/XC1/XRES1A/B 0.386137f
C154 XA5/EN XA5/XA1/XA1/MP3/G 0.095485f
C155 XA20/CNO XA4/EN 0.457818f
C156 XA20/CPO XA2/CN0 0.06056f
C157 EN AVSS 1.655709f
C158 XA20/CPO XA2/EN 0.378571f
C159 D<4> XA3/CN0 1.581234f
C160 AVSS D<1> 1.876198f
C161 XA1/CN1 XA1/CP0 0.174582f
C162 SARN AVDD 0.08218f
C163 XA20/XA9/A XA20/CNO 0.101825f
C164 XA0/CEIN SAR_IP 0.059924f
C165 VREF XA6/CN0 0.061065f
C166 D<7> XA1/CN1 2.492607f
C167 XA1/CN1 XA0/CN0 0.495948f
C168 XA2/CN0 XA3/CN0 2.194396f
C169 XA2/CP0 AVSS 0.193422f
C170 D<6> XA1/CP0 4.060233f
C171 VREF XA6/CEO 0.348791f
C172 XA20/CPO XA3/XA1/XA2/Y 0.078271f
C173 SARN XB2/XA4/GNG 1.624341f
C174 D<3> CK_SAMPLE 0.100705f
C175 D<7> D<6> 0.073624f
C176 XA20/CPO XA1/CN1 0.267213f
C177 D<6> XA0/CN0 0.058151f
C178 VREF AVSS 1.049192f
C179 DONE AVSS 0.493308f
C180 XA5/CN0 D<7> 0.073409f
C181 XA5/CN0 XA0/CN0 0.09322f
C182 XA0/XA4/A XA20/CNO 0.212166f
C183 XA4/DONE AVSS 0.2733f
C184 XA20/CPO D<6> 0.062597f
C185 XA1/CN1 XA3/CN0 0.066079f
C186 AVDD XA3/EN 0.79199f
C187 XA0/CEO XA1/XA12/A 0.084465f
C188 XA5/CN0 XA20/CPO 0.068343f
C189 D<7> XA6/CN0 0.077804f
C190 XA0/CN0 XA6/CN0 0.077861f
C191 XA7/EN XA6/CN0 0.056481f
C192 XA6/EN CK_SAMPLE 0.09249f
C193 XA5/CN0 XA3/CN0 0.095106f
C194 XA4/CN0 CK_SAMPLE 0.070685f
C195 XA1/CP0 AVSS 0.19218f
C196 XA20/CPO XA6/CN0 0.068386f
C197 XA0/CEIN AVDD 9.065545f
C198 D<7> AVSS 1.140293f
C199 AVSS XA0/CN0 0.144488f
C200 XA0/CEO AVSS 0.267201f
C201 XA7/EN AVSS 0.231176f
C202 D<3> XA4/CN0 1.470811f
C203 XA3/EN XA2/XA1/XA1/MP3/G 0.058161f
C204 XA6/XA1/XA2/Y XA20/CPO 0.069955f
C205 XA3/CN0 XA6/CN0 0.071838f
C206 XA20/CPO AVSS 1.94788f
C207 XA7/XA11/A XA6/CEO 0.097953f
C208 AVDD XA7/ENO 0.076028f
C209 D<4> XA4/EN 0.094074f
C210 EN XA2/XA2/A 0.11426f
C211 XA4/CN0 XA4/CP0 0.125928f
C212 DONE XA7/XA9/A 0.052108f
C213 XA20/CNO D<4> 0.063433f
C214 EN D<5> 0.06282f
C215 XA3/CN0 AVSS 0.25506f
C216 XA7/CEO XA7/XA12/A 0.069744f
C217 DONE XA7/XA9/B 0.27523f
C218 XA5/XA4/A EN 0.088236f
C219 XA20/CNO XA2/CN0 0.058198f
C220 XA20/CNO XA2/EN 0.457819f
C221 XA2/CP0 D<5> 3.965242f
C222 XB2/XA4/GNG XDAC2/XC1/XRES1A/B 0.386137f
C223 SARP XB1/M4/G 0.144008f
C224 EN XA3/EN 0.311923f
C225 VREF D<5> 0.083365f
C226 XA0/CP0 XA0/CP1 4.153562f
C227 CK_SAMPLE_BSSW AVSS 0.75049f
C228 SARP SAR_IP 0.279047f
C229 XA0/CP0 XA2/CN1 0.144778f
C230 CK_SAMPLE XA1/CN0 0.071036f
C231 XA5/CEO XA5/XA11/A 0.13078f
C232 XA20/CNO XA1/CN1 0.19102f
C233 XA1/EN CK_SAMPLE 0.092446f
C234 D<3> XA1/CN0 0.07156f
C235 VREF XA3/EN 0.175304f
C236 XA20/CNO XA3/XA4/A 0.286128f
C237 XA20/CNO D<6> 0.054548f
C238 SARN D<7> 0.059383f
C239 SARN XA0/CN0 0.109275f
C240 XA5/CN0 XA20/CNO 0.064438f
C241 XA3/XA11/A XA2/CEO 0.068277f
C242 XA1/CP0 D<5> 0.762697f
C243 XA5/EN CK_SAMPLE 0.092446f
C244 SARN XA20/CPO 0.096247f
C245 D<7> D<5> 0.073518f
C246 EN XA7/ENO 0.096521f
C247 XA0/CN0 D<5> 0.058768f
C248 XA5/CP0 AVDD -0.052017f
C249 XA0/XA1/XA2/Y XA20/CPO 0.069784f
C250 XA0/CEIN VREF 0.054033f
C251 XA4/CEO AVDD 1.256112f
C252 XA20/CNO XA6/CN0 0.066819f
C253 XA20/CPO D<5> 0.061883f
C254 XA3/XA1/XA1/MP3/G XA3/EN 0.095485f
C255 VREF D<0> 0.078578f
C256 XA4/CN0 XA1/CN0 0.066599f
C257 XA5/CEO AVSS 0.43736f
C258 XA4/EN AVSS 0.355405f
C259 SARP AVDD 0.073696f
C260 VREF XA7/ENO 0.175304f
C261 CK_SAMPLE XA0/CP1 0.100695f
C262 XA20/CNO AVSS 2.172184f
C263 XA2/CN0 D<4> 0.070556f
C264 XA20/CPO XA3/EN 0.251162f
C265 XA5/EN XA6/EN 1.263077f
C266 XA5/EN XA4/CN0 0.056535f
C267 D<3> XA2/CN1 0.105016f
C268 EN XA3/XA2/A 0.11418f
C269 XA3/EN XA3/CN0 0.070743f
C270 XA2/CEO AVSS 0.266939f
C271 AVDD CK_SAMPLE 4.279234f
C272 D<4> XA1/CN1 0.066004f
C273 EN XA0/CP0 0.060919f
C274 AVDD XA3/CEO 0.342105f
C275 XA7/EN XA7/ENO 0.779051f
C276 XA1/XA11/A XA1/CEO 0.13078f
C277 XA2/CN0 XA1/CN1 0.066278f
C278 XA1/CN1 XA2/EN 0.107883f
C279 D<2> CK_SAMPLE 0.1008f
C280 XA4/CN0 XA2/CN1 0.073436f
C281 XA20/XA9/Y CK_SAMPLE 0.069412f
C282 XA20/CPO XA7/ENO 0.092502f
C283 D<3> D<2> 0.983626f
C284 D<6> XA2/EN 0.081832f
C285 XA5/CN0 XA2/CN0 0.084337f
C286 XA4/CP0 AVDD -0.052017f
C287 EN XA1/XA2/A 0.11418f
C288 XA1/EN XA1/CN0 0.061773f
C289 XA0/CEIN XB1/CKN 0.100039f
C290 XA6/EN AVDD 0.11184f
C291 XA6/CP0 XA6/CN0 0.125928f
C292 XA0/CEIN CK_SAMPLE_BSSW 6.834396f
C293 XA4/CN0 AVDD 2.483943f
C294 AVDD XA7/CEO 0.348014f
C295 SARN XA20/CNO 0.092221f
C296 XA20/XA3/CO XA20/CPO 0.104539f
C297 SARN XB2/M4/G 0.24502f
C298 XA2/CN0 XA6/CN0 0.071524f
C299 XA20/XA9/A SARN 0.113134f
C300 XA4/CEO VREF 0.348781f
C301 D<6> XA1/CN1 0.616721f
C302 XA5/CN0 XA1/CN1 0.065942f
C303 D<4> AVSS 1.856228f
C304 XA6/EN D<2> 0.094074f
C305 XA20/CNO D<5> 0.054559f
C306 CK_SAMPLE XA7/CN0 0.071036f
C307 EN XA6/XA4/A 0.088464f
C308 XA4/CN0 D<2> 0.073269f
C309 SARN SAR_IN 0.271831f
C310 XA0/CP0 XA1/CP0 1.795396f
C311 XA1/DONE AVSS 0.267946f
C312 XA2/CN0 AVSS 0.127755f
C313 XA2/EN AVSS 0.296958f
C314 XA5/XA4/A XA20/CNO 0.286129f
C315 D<7> XA0/CP0 0.111006f
C316 XA0/CP0 XA0/CN0 3.564213f
C317 CK_SAMPLE D<1> 0.100705f
C318 XA1/CN1 XA6/CN0 0.070367f
C319 XA4/EN XA3/EN 1.263078f
C320 D<3> EN 0.070973f
C321 XA20/CNO XA3/EN 0.302924f
C322 D<3> D<1> 0.181155f
C323 XA20/CPO XA0/CP0 0.057707f
C324 XA1/CN0 XA2/CN1 0.547507f
C325 XA20/XA3/N1 SARN 0.135724f
C326 XA5/CN0 XA6/CN0 1.883929f
C327 XA1/CN1 AVSS 1.316495f
C328 XB1/XA3/B AVSS 1.491396f
C329 XA3/XA12/A XA3/CEO 0.264747f
C330 CK_SAMPLE DONE 0.086955f
C331 VREF CK_SAMPLE 1.866437f
C332 XA20/CNO XA7/XA4/A 0.304482f
C333 SARP D<7> 0.187721f
C334 XA20/XA9/A XA7/XA4/A 0.11382f
C335 D<6> AVSS 1.853472f
C336 D<3> VREF 0.083365f
C337 XB1/XA4/GNG AVSS 1.208553f
C338 XA5/CN0 AVSS 0.234223f
C339 CK_SAMPLE XA2/XA9/B 0.07743f
C340 XA0/CEIN XB2/M4/G 0.111673f
C341 AVDD XA1/CN0 2.473342f
C342 XA6/EN EN 0.235384f
C343 SARP XA20/CPO 0.054401f
C344 XA4/CN0 EN 0.073779f
C345 XA4/CN0 D<1> 0.072622f
C346 AVDD XA1/EN 0.791991f
C347 XA0/CEIN SAR_IN 0.064238f
C348 XA20/CNO XA7/ENO 0.088037f
C349 AVSS XA6/CN0 0.279681f
C350 D<2> XA1/CN0 0.082802f
C351 XA5/EN AVDD 0.791989f
C352 CK_SAMPLE XA0/CN0 0.070685f
C353 XA7/EN CK_SAMPLE 0.092446f
C354 XA6/EN VREF 0.175304f
C355 AVSS XA6/CEO 0.276115f
C356 XA4/CN0 VREF 0.061065f
C357 XA2/CN1 XA0/CP1 1.265362f
C358 D<3> D<7> 0.073432f
C359 D<4> D<5> 0.356702f
C360 D<3> XA0/CN0 0.08508f
C361 DONE XA7/CEO 0.119439f
C362 XA5/CEO XA5/XA12/A 0.264747f
C363 XA1/EN XA1/XA1/XA1/MP3/G 0.095485f
C364 XB2/XA4/GNG XDAC2/XC1/XRES16/B 0.107427f
C365 XA0/XA2/A EN 0.11426f
C366 XA5/EN D<2> 0.070574f
C367 D<3> XA20/CPO 0.071226f
C368 AVDD XA1/CEO 0.342105f
C369 CK_SAMPLE XA3/CN0 0.071036f
C370 D<4> XA3/EN 0.070945f
C371 D<3> XA3/CN0 0.081287f
C372 XA2/CN0 XA3/EN 0.052744f
C373 XA4/CN0 D<7> 0.073427f
C374 XA4/CN0 XA0/CN0 0.072808f
C375 XA1/XA11/A XA0/CEO 0.068277f
C376 XA1/CN1 D<5> 0.06654f
C377 EN XA1/CN0 0.066764f
C378 XA1/CN0 D<1> 0.079158f
C379 XA5/CN1 XA5/CN0 0.051393f
C380 XA20/CNO XA0/CP0 0.054091f
C381 XA6/EN XA20/CPO 0.378571f
C382 D<2> XA2/CN1 0.137975f
C383 XA1/EN EN 0.315013f
C384 XA4/CN0 XA20/CPO 0.068386f
C385 D<6> D<5> 1.055163f
C386 XA2/CP0 XA1/CN0 0.063884f
C387 XA5/CEO XA4/CEO 0.431793f
C388 AVDD XB2/XA3/B 0.185337f
C389 XA4/CN0 XA3/CN0 1.410099f
C390 XA5/EN EN 0.311923f
C391 VREF XA1/CN0 0.061065f
C392 XA1/EN VREF 0.175304f
C393 XA4/XA4/A EN 0.088464f
C394 XA20/XA9/A SARP 0.092582f
C395 SARN AVSS 3.513515f
C396 AVDD XA3/CP0 -0.052017f
C397 XA4/XA2/A EN 0.11426f
C398 SARP SAR_IN 0.091622f
C399 XA5/EN VREF 0.175304f
C400 AVSS D<5> 1.873407f
C401 EN XA0/CP1 0.068097f
C402 XA20/CNO XA6/XA4/A 0.212166f
C403 XA1/CN0 XA1/CP0 3.345594f
C404 EN XA2/CN1 0.099756f
C405 XA20/CPO XA2/XA1/XA2/Y 0.069955f
C406 XA2/CN1 D<1> 0.077649f
C407 CK_SAMPLE XA4/EN 0.09249f
C408 D<7> XA1/CN0 0.073792f
C409 XA1/EN XA1/CP0 0.05876f
C410 XA1/CN0 XA0/CN0 2.961017f
C411 XA2/DONE AVSS 0.2733f
C412 XA20/XA9/A CK_SAMPLE 0.169353f
C413 XA1/EN XA0/CN0 0.052744f
C414 XA3/EN AVSS 0.214912f
C415 XA2/CP0 XA2/CN1 0.110086f
C416 D<3> XA20/CNO 0.063902f
C417 XA20/CPO XA1/CN0 0.060404f
C418 VREF XA0/CP1 0.083365f
C419 EN XA6/XA2/A 0.11426f
C420 AVDD EN 2.755226f
C421 XA1/EN XA20/CPO 0.251162f
C422 XA0/CP0 D<4> 0.207798f
C423 XA1/CN0 XA3/CN0 0.06759f
C424 XA3/DONE AVSS 0.267946f
C425 XA0/CEIN AVSS 2.00975f
C426 XA5/EN XA20/CPO 0.251162f
C427 D<2> EN 0.07107f
C428 D<2> D<1> 1.784246f
C429 XA2/CEO XA3/CEO 0.431793f
C430 XA6/EN XA20/CNO 0.457818f
C431 AVDD VREF 15.778251f
C432 XA4/CN0 XA20/CNO 0.066024f
C433 XA5/XA9/B CK_SAMPLE 0.078405f
C434 XA0/CEO XA1/CEO 0.431792f
C435 XA1/CP0 XA2/CN1 0.143675f
C436 D<7> XA0/CP1 0.831597f
C437 D<7> XA2/CN1 0.074905f
C438 XA2/CN1 XA0/CN0 0.0725f
C439 XA0/CP0 XA1/CN1 0.139477f
C440 D<2> VREF 0.083401f
C441 XA1/DONE XA1/XA9/B 0.061581f
C442 XA3/XA1/XA1/MN2/S XA4/EN 0.064012f
C443 XA20/CPO XA0/CP1 0.061883f
C444 XA20/CPO XA2/CN1 0.255235f
C445 XA2/CN1 XA2/XA4/A 0.06833f
C446 XA0/CP0 D<6> 0.81476f
C447 XA20/XA3/CO AVSS 0.073081f
C448 AVDD XA0/CN0 2.477148f
C449 AVDD XA0/CEO 1.256112f
C450 XA7/EN AVDD 0.809492f
C451 XA4/XA1/XA2/Y XA20/CPO 0.069955f
C452 XA4/CEO XA5/XA11/A 0.068277f
C453 XA2/CN1 XA3/CN0 0.074031f
C454 XA5/CN0 XA5/CP0 0.125928f
C455 CK_SAMPLE D<4> 0.1008f
C456 SARP XA1/CN1 0.062345f
C457 EN D<1> 0.070973f
C458 AVDD XA20/CPO 2.513656f
C459 D<3> D<4> 0.665607f
C460 CK_SAMPLE XA2/CN0 0.070685f
C461 CK_SAMPLE XA2/EN 0.09249f
C462 D<2> D<7> 0.086175f
C463 D<2> XA0/CN0 0.099255f
C464 SARP XB1/XA4/GNG 1.624342f
C465 EN XA2/CP0 0.058498f
C466 D<3> XA2/CN0 0.073287f
C467 XA0/CEIN SARN 0.265285f
C468 XA20/CNO XA7/XA2/A 0.076673f
C469 AVDD XA3/CN0 2.477465f
C470 EN XA1/XA4/A 0.088236f
C471 XA0/CP0 AVSS 0.207167f
C472 XA20/CNO XA1/CN0 0.056881f
C473 XA3/DONE XA3/XA9/B 0.061581f
C474 D<2> XA20/CPO 0.071873f
C475 VREF EN 0.66498f
C476 VREF D<1> 0.083365f
C477 XA1/EN XA20/CNO 0.302765f
C478 XA3/XA11/A XA3/CEO 0.13078f
C479 D<2> XA3/CN0 0.073198f
C480 XA4/CEO AVSS 0.266939f
C481 D<3> XA1/CN1 0.06595f
C482 CK_SAMPLE_BSSW AVDD 14.874317f
C483 XA7/EN XA6/XA1/XA1/MP3/G 0.058161f
C484 CK_SAMPLE D<6> 0.1008f
C485 XA3/CN0 XA3/CP0 0.125928f
C486 XA5/EN XA20/CNO 0.302925f
C487 XA5/CN0 CK_SAMPLE 0.071036f
C488 XA4/CN0 XA2/CN0 0.068184f
C489 SARP AVSS 0.540564f
C490 XA4/XA4/A XA20/CNO 0.212166f
C491 AVSS XA6/DONE 0.2733f
C492 EN XA1/CP0 0.058341f
C493 D<7> EN 0.334727f
C494 EN XA0/CN0 0.068738f
C495 XA4/XA9/B CK_SAMPLE 0.07743f
C496 XA7/EN EN 0.173811f
C497 D<7> D<1> 0.077821f
C498 XA0/CN0 D<1> 0.232115f
C499 CK_SAMPLE XA6/CN0 0.070685f
C500 XA2/CP0 XA1/CP0 1.213936f
C501 XA4/CN0 XA1/CN1 0.06599f
C502 XA20/CPO EN 0.728023f
C503 XA20/CNO XA0/CP1 0.054559f
C504 XA20/CPO XA7/XA1/XA2/Y 0.081064f
C505 D<7> XA2/CP0 0.073351f
C506 XA2/CP0 XA0/CN0 1.220085f
C507 EN XA2/XA4/A 0.088464f
C508 XA20/CPO D<1> 0.071226f
C509 XA20/CNO XA2/CN1 0.188581f
C510 CK_SAMPLE AVSS 2.799086f
C511 XA6/EN XA5/CN0 0.13801f
C512 VREF XA0/CN0 0.061065f
C513 VREF XA0/CEO 0.348781f
C514 XA20/CPO XA2/CP0 0.057707f
C515 XA7/EN VREF 0.175304f
C516 EN XA3/CN0 0.073639f
C517 XA4/CN0 XA5/CN0 1.362054f
C518 XA3/CN0 D<1> 0.072559f
C519 D<3> AVSS 1.876198f
C520 XA3/CEO AVSS 0.437359f
C521 XA1/XA4/A XA2/XA4/A 0.082663f
C522 XA7/XA9/MN1/a_324_334# 0 0.360407f
C523 XA7/XA9/MN0/a_324_n18# 0 0.360407f
C524 XA7/XA9/A 0 1.250071f
C525 XA7/XA7/MN0/a_324_n18# 0 0.360407f
C526 XA7/XA8/MN0/a_324_n18# 0 0.360407f
C527 XA7/XA9/B 0 1.15806f
C528 XA7/XA6/MN0/a_324_n18# 0 0.360407f
C529 XA7/XA4/A 0 2.621765f
C530 XA7/XA4/MN0/a_324_n18# 0 0.360407f
C531 XA7/CP0 0 2.4163f
C532 XA7/CN0 0 0.312365f
C533 XA7/XA5/MN0/a_324_n18# 0 0.360407f
C534 XA7/CN1 0 2.428168f
C535 D<0> 0 0.412798f
C536 XA7/XA3/MN0/a_324_n18# 0 0.360407f
C537 XA7/XA2/A 0 2.030764f
C538 XA7/XA2/MN0/a_324_n18# 0 0.360407f
C539 XA7/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C540 XA7/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C541 XA7/XA1/XA2/Y 0 1.060197f
C542 XA7/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C543 XA7/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C544 XA7/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C545 XA7/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C546 XA7/XA1/XA1/MP3/G 0 0.827484f
C547 XA7/XA1/XA1/MN2/S 0 0.200627f
C548 XA7/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C549 XA7/ENO 0 1.582724f
C550 XA7/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C551 XA7/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C552 XA7/XA13/MN1/a_324_334# 0 0.422f
C553 XA7/XA13/MP1/a_216_334# 0 0.091271f
C554 XA7/CEO 0 1.316615f
C555 XA7/XA12/MN0/a_324_n18# 0 0.360407f
C556 XA7/XA13/MN1/a_324_n18# 0 0.360407f
C557 XA7/XA12/A 0 0.755669f
C558 XA7/XA11/MN0/a_324_n18# 0 0.360407f
C559 XA6/CEO 0 1.009021f
C560 XA7/XA11/A 0 0.662715f
C561 XA7/XA9/Y 0 0.718246f
C562 XA6/XA9/MN1/a_324_334# 0 0.360407f
C563 XA6/XA9/MN0/a_324_n18# 0 0.360407f
C564 XA6/XA9/A 0 1.250071f
C565 XA6/DONE 0 0.13094f
C566 XA6/XA7/MN0/a_324_n18# 0 0.360407f
C567 XA6/XA8/MN0/a_324_n18# 0 0.360407f
C568 XA6/XA9/B 0 1.15806f
C569 XA6/XA6/MN0/a_324_n18# 0 0.360407f
C570 XA6/XA4/A 0 2.621765f
C571 XA6/XA4/MN0/a_324_n18# 0 0.360407f
C572 XA6/CP0 0 2.4163f
C573 XA6/CN0 0 4.160099f
C574 XA6/XA5/MN0/a_324_n18# 0 0.360407f
C575 XA6/CN1 0 2.428168f
C576 D<1> 0 4.424545f
C577 XA6/XA3/MN0/a_324_n18# 0 0.360407f
C578 XA6/XA2/A 0 2.030764f
C579 XA6/XA2/MN0/a_324_n18# 0 0.360407f
C580 XA6/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C581 XA6/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C582 XA6/XA1/XA2/Y 0 1.060197f
C583 XA6/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C584 XA6/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C585 XA6/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C586 XA6/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C587 XA6/XA1/XA1/MP3/G 0 0.827484f
C588 XA6/XA1/XA1/MN2/S 0 0.200627f
C589 XA6/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C590 XA7/EN 0 3.856368f
C591 XA6/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C592 XA6/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C593 XA6/XA13/MN1/a_324_334# 0 0.422f
C594 XA6/XA13/MP1/a_216_334# 0 0.091271f
C595 XA6/XA12/MN0/a_324_n18# 0 0.360407f
C596 XA6/XA13/MN1/a_324_n18# 0 0.360407f
C597 XA6/XA12/A 0 0.755669f
C598 XA6/XA11/MN0/a_324_n18# 0 0.360407f
C599 XA5/CEO 0 1.104751f
C600 XA6/XA11/A 0 0.662715f
C601 XA6/XA9/Y 0 0.718246f
C602 XA5/XA9/MN1/a_324_334# 0 0.360407f
C603 XA5/XA9/MN0/a_324_n18# 0 0.360407f
C604 XA5/XA9/A 0 1.250071f
C605 XA5/DONE 0 0.123486f
C606 XA5/XA7/MN0/a_324_n18# 0 0.360407f
C607 XA5/XA8/MN0/a_324_n18# 0 0.360407f
C608 XA5/XA9/B 0 1.15806f
C609 XA5/XA6/MN0/a_324_n18# 0 0.360407f
C610 XA5/XA4/A 0 2.621765f
C611 XA5/XA4/MN0/a_324_n18# 0 0.360407f
C612 XA5/CP0 0 2.4163f
C613 XA5/CN0 0 3.052303f
C614 XA5/XA5/MN0/a_324_n18# 0 0.360407f
C615 XA5/CN1 0 2.428168f
C616 D<2> 0 3.706573f
C617 XA5/XA3/MN0/a_324_n18# 0 0.360407f
C618 XA5/XA2/A 0 2.030764f
C619 XA5/XA2/MN0/a_324_n18# 0 0.360407f
C620 XA5/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C621 XA5/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C622 XA5/XA1/XA2/Y 0 1.060197f
C623 XA5/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C624 XA5/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C625 XA5/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C626 XA5/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C627 XA5/XA1/XA1/MP3/G 0 0.827484f
C628 XA5/XA1/XA1/MN2/S 0 0.200627f
C629 XA5/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C630 XA6/EN 0 3.679756f
C631 XA5/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C632 XA5/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C633 XA5/XA13/MN1/a_324_334# 0 0.422f
C634 XA5/XA13/MP1/a_216_334# 0 0.091271f
C635 XA5/XA12/MN0/a_324_n18# 0 0.360407f
C636 XA5/XA13/MN1/a_324_n18# 0 0.360407f
C637 XA5/XA12/A 0 0.755669f
C638 XA5/XA11/MN0/a_324_n18# 0 0.360407f
C639 XA4/CEO 0 1.086041f
C640 XA5/XA11/A 0 0.662715f
C641 XA5/XA9/Y 0 0.718246f
C642 XA4/XA9/MN1/a_324_334# 0 0.360407f
C643 XA4/XA9/MN0/a_324_n18# 0 0.360407f
C644 XA4/XA9/A 0 1.250071f
C645 XA4/DONE 0 0.13094f
C646 XA4/XA7/MN0/a_324_n18# 0 0.360407f
C647 XA4/XA8/MN0/a_324_n18# 0 0.360407f
C648 XA4/XA9/B 0 1.15806f
C649 XA4/XA6/MN0/a_324_n18# 0 0.360407f
C650 XA4/XA4/A 0 2.621765f
C651 XA4/XA4/MN0/a_324_n18# 0 0.360407f
C652 XA4/CP0 0 2.4163f
C653 XA4/CN0 0 2.237548f
C654 XA4/XA5/MN0/a_324_n18# 0 0.360407f
C655 XA4/CN1 0 2.428168f
C656 D<3> 0 2.560026f
C657 XA4/XA3/MN0/a_324_n18# 0 0.360407f
C658 XA4/XA2/A 0 2.030764f
C659 XA4/XA2/MN0/a_324_n18# 0 0.360407f
C660 XA4/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C661 XA4/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C662 XA4/XA1/XA2/Y 0 1.060197f
C663 XA4/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C664 XA4/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C665 XA4/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C666 XA4/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C667 XA4/XA1/XA1/MP3/G 0 0.827484f
C668 XA4/XA1/XA1/MN2/S 0 0.200627f
C669 XA4/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C670 XA5/EN 0 3.635208f
C671 XA4/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C672 XA4/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C673 XA4/XA13/MN1/a_324_334# 0 0.422f
C674 XA4/XA13/MP1/a_216_334# 0 0.091271f
C675 XA4/XA12/MN0/a_324_n18# 0 0.360407f
C676 XA4/XA13/MN1/a_324_n18# 0 0.360407f
C677 XA4/XA12/A 0 0.755669f
C678 XA4/XA11/MN0/a_324_n18# 0 0.360407f
C679 XA3/CEO 0 1.107611f
C680 XA4/XA11/A 0 0.662715f
C681 XA4/XA9/Y 0 0.718246f
C682 XA3/XA9/MN1/a_324_334# 0 0.360407f
C683 XA3/XA9/MN0/a_324_n18# 0 0.360407f
C684 XA3/XA9/A 0 1.250071f
C685 XA3/DONE 0 0.123486f
C686 XA3/XA7/MN0/a_324_n18# 0 0.360407f
C687 XA3/XA8/MN0/a_324_n18# 0 0.360407f
C688 XA3/XA9/B 0 1.15806f
C689 XA3/XA6/MN0/a_324_n18# 0 0.360407f
C690 XA3/XA4/A 0 2.621765f
C691 XA3/XA4/MN0/a_324_n18# 0 0.360407f
C692 XA3/CP0 0 2.4163f
C693 XA3/CN0 0 3.224855f
C694 XA3/XA5/MN0/a_324_n18# 0 0.360407f
C695 XA3/CN1 0 2.428168f
C696 D<4> 0 3.08566f
C697 XA3/XA3/MN0/a_324_n18# 0 0.360407f
C698 XA3/XA2/A 0 2.030764f
C699 XA3/XA2/MN0/a_324_n18# 0 0.360407f
C700 XA3/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C701 XA3/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C702 XA3/XA1/XA2/Y 0 1.060197f
C703 XA3/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C704 XA3/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C705 XA3/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C706 XA3/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C707 XA3/XA1/XA1/MP3/G 0 0.827484f
C708 XA3/XA1/XA1/MN2/S 0 0.200627f
C709 XA3/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C710 XA4/EN 0 3.720665f
C711 XA3/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C712 XA3/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C713 XA3/XA13/MN1/a_324_334# 0 0.422f
C714 XA3/XA13/MP1/a_216_334# 0 0.091271f
C715 XA3/XA12/MN0/a_324_n18# 0 0.360407f
C716 XA3/XA13/MN1/a_324_n18# 0 0.360407f
C717 XA3/XA12/A 0 0.755669f
C718 XA3/XA11/MN0/a_324_n18# 0 0.360407f
C719 XA2/CEO 0 1.085281f
C720 XA3/XA11/A 0 0.662715f
C721 XA3/XA9/Y 0 0.718246f
C722 XA2/XA9/MN1/a_324_334# 0 0.360407f
C723 XA2/XA9/MN0/a_324_n18# 0 0.360407f
C724 XA2/XA9/A 0 1.250071f
C725 XA2/DONE 0 0.13094f
C726 XA2/XA7/MN0/a_324_n18# 0 0.360407f
C727 XA2/XA8/MN0/a_324_n18# 0 0.360407f
C728 XA2/XA9/B 0 1.15806f
C729 XA2/XA6/MN0/a_324_n18# 0 0.360407f
C730 XA2/XA4/A 0 2.621765f
C731 XA2/XA4/MN0/a_324_n18# 0 0.360407f
C732 XA2/CP0 0 4.49437f
C733 XA2/CN0 0 2.820252f
C734 XA2/XA5/MN0/a_324_n18# 0 0.360407f
C735 XA2/CN1 0 6.112935f
C736 XA2/XA3/MN0/a_324_n18# 0 0.360407f
C737 XA2/XA2/A 0 2.030764f
C738 XA2/XA2/MN0/a_324_n18# 0 0.360407f
C739 XA2/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C740 XA2/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C741 XA2/XA1/XA2/Y 0 1.060197f
C742 XA2/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C743 XA2/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C744 XA2/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C745 XA2/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C746 XA2/XA1/XA1/MP3/G 0 0.827484f
C747 XA2/XA1/XA1/MN2/S 0 0.200627f
C748 XA2/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C749 XA3/EN 0 3.784028f
C750 XA2/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C751 XA2/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C752 XA2/XA13/MN1/a_324_334# 0 0.422f
C753 XA2/XA13/MP1/a_216_334# 0 0.091271f
C754 XA2/XA12/MN0/a_324_n18# 0 0.360407f
C755 XA2/XA13/MN1/a_324_n18# 0 0.360407f
C756 XA2/XA12/A 0 0.755669f
C757 XA2/XA11/MN0/a_324_n18# 0 0.360407f
C758 XA1/CEO 0 1.104751f
C759 XA2/XA11/A 0 0.662715f
C760 XA2/XA9/Y 0 0.718246f
C761 XA1/XA9/MN1/a_324_334# 0 0.360407f
C762 XA1/XA9/MN0/a_324_n18# 0 0.360407f
C763 XA1/XA9/A 0 1.250071f
C764 XA1/DONE 0 0.123486f
C765 XA1/XA7/MN0/a_324_n18# 0 0.360407f
C766 XA1/XA8/MN0/a_324_n18# 0 0.360407f
C767 XA1/XA9/B 0 1.15806f
C768 XA1/XA6/MN0/a_324_n18# 0 0.360407f
C769 XA1/XA4/A 0 2.621765f
C770 XA1/XA4/MN0/a_324_n18# 0 0.360407f
C771 XA1/CP0 0 4.486094f
C772 XA1/CN0 0 2.798774f
C773 XA1/XA5/MN0/a_324_n18# 0 0.360407f
C774 XA1/CN1 0 4.70217f
C775 D<6> 0 2.989828f
C776 XA1/XA3/MN0/a_324_n18# 0 0.360407f
C777 XA1/XA2/A 0 2.030764f
C778 XA1/XA2/MN0/a_324_n18# 0 0.360407f
C779 XA1/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C780 XA1/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C781 XA1/XA1/XA2/Y 0 1.060197f
C782 XA1/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C783 XA1/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C784 XA1/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C785 XA1/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C786 XA1/XA1/XA1/MP3/G 0 0.827484f
C787 XA1/XA1/XA1/MN2/S 0 0.200627f
C788 XA1/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C789 XA2/EN 0 3.720665f
C790 XA1/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C791 XA1/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C792 XA1/XA13/MN1/a_324_334# 0 0.422f
C793 XA1/XA13/MP1/a_216_334# 0 0.091271f
C794 XA1/XA12/MN0/a_324_n18# 0 0.360407f
C795 XA1/XA13/MN1/a_324_n18# 0 0.360407f
C796 XA1/XA12/A 0 0.755669f
C797 XA1/XA11/MN0/a_324_n18# 0 0.360407f
C798 XA0/CEO 0 1.083361f
C799 XA1/XA11/A 0 0.662715f
C800 XA1/XA9/Y 0 0.718246f
C801 XB2/XA7/MN1/a_324_n18# 0 0.359583f
C802 XB2/XA5b/MN1/a_324_n18# 0 0.422415f
C803 XB2/XA5b/MP1/a_216_n18# 0 0.091271f
C804 XB2/XA1/Y 0 0.690197f
C805 XB2/CKN 0 1.768971f
C806 XB2/XA4/MN0/a_324_n18# 0 0.359583f
C807 XB2/XA5/MN1/a_324_334# 0 0.422f
C808 XB2/XA5/MP1/a_216_334# 0 0.091271f
C809 XB2/XA3/MP0/S 0 0.743486f
C810 XB2/XA3/MN0/a_324_n18# 0 0.359583f
C811 XB2/XA2/MP0/G 0 0.708335f
C812 XB2/XA7/MN1/a_324_334# 0 0.359583f
C813 XB2/XA5/MN1/a_324_n18# 0 0.360407f
C814 XB2/XA1/MP0/G 0 0.788614f
C815 XB2/XA4/MN1/a_324_334# 0 0.359583f
C816 XB2/XA0/MN0/a_324_n18# 0 0.359583f
C817 XB2/M8/a_324_n18# 0 0.356977f
C818 XB2/M8/a_324_334# 0 0.422f
C819 XB2/M6/a_324_n18# 0 0.356977f
C820 XB2/M7/a_324_n18# 0 0.356977f
C821 XB2/XA3/B 0 54.41209f
C822 XB2/XA4/GNG 0 53.065117f
C823 XB2/M5/a_324_n18# 0 0.356977f
C824 XB2/M3/a_324_n18# 0 0.356977f
C825 XB2/M4/a_324_n18# 0 0.356977f
C826 XB2/M4/G 0 2.475647f
C827 SAR_IN 0 1.184896f
C828 XB2/M1/a_324_n18# 0 0.422415f
C829 XB2/M2/a_324_n18# 0 0.356977f
C830 XA0/XA9/MN1/a_324_334# 0 0.360407f
C831 XA0/XA9/MN0/a_324_n18# 0 0.360407f
C832 XA0/XA9/A 0 1.250071f
C833 XA0/DONE 0 0.134046f
C834 XA0/XA7/MN0/a_324_n18# 0 0.360407f
C835 XA0/XA8/MN0/a_324_n18# 0 0.360407f
C836 XA0/XA9/B 0 1.15806f
C837 CK_SAMPLE 0 15.793598f
C838 XA0/XA6/MN0/a_324_n18# 0 0.360407f
C839 XA0/XA4/A 0 2.621765f
C840 XA0/XA4/MN0/a_324_n18# 0 0.360407f
C841 XA0/CP0 0 8.48089f
C842 XA0/XA5/MN0/a_324_n18# 0 0.360407f
C843 VREF 0 27.717136f
C844 D<7> 0 7.541619f
C845 XA0/XA3/MN0/a_324_n18# 0 0.360407f
C846 XA0/XA2/A 0 2.030764f
C847 XA0/XA2/MN0/a_324_n18# 0 0.360407f
C848 XA0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C849 EN 0 4.718864f
C850 XA0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C851 XA0/XA1/XA2/Y 0 1.060197f
C852 XA0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C853 XA0/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C854 XA20/CPO 0 11.091676f
C855 XA0/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C856 XA20/CNO 0 12.667546f
C857 XA0/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C858 XA0/XA1/XA1/MP3/G 0 0.827484f
C859 XA0/XA1/XA1/MN2/S 0 0.200627f
C860 XA0/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C861 XA1/EN 0 3.794638f
C862 XA0/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C863 AVDD 0 0.517971p
C864 XA0/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C865 XA0/XA13/MN1/a_324_334# 0 0.422f
C866 XA0/XA13/MP1/a_216_334# 0 0.091271f
C867 XA0/XA12/MN0/a_324_n18# 0 0.360407f
C868 XA0/XA13/MN1/a_324_n18# 0 0.360407f
C869 XA0/XA12/A 0 0.755669f
C870 XA0/XA11/MN0/a_324_n18# 0 0.360407f
C871 XA0/XA11/A 0 0.662715f
C872 XA0/XA9/Y 0 0.718246f
C873 XB1/XA7/MN1/a_324_n18# 0 0.359583f
C874 AVSS 0 0.14072p
C875 XB1/XA5b/MN1/a_324_n18# 0 0.422415f
C876 XB1/XA5b/MP1/a_216_n18# 0 0.091271f
C877 XB1/XA1/Y 0 0.690197f
C878 XB1/CKN 0 1.768971f
C879 XB1/XA4/MN0/a_324_n18# 0 0.359583f
C880 XB1/XA5/MN1/a_324_334# 0 0.422f
C881 XB1/XA5/MP1/a_216_334# 0 0.091271f
C882 XB1/XA3/MP0/S 0 0.743486f
C883 XB1/XA3/MN0/a_324_n18# 0 0.359583f
C884 XB1/XA2/MP0/G 0 0.708335f
C885 XB1/XA7/MN1/a_324_334# 0 0.359583f
C886 XB1/XA5/MN1/a_324_n18# 0 0.360407f
C887 XB1/XA1/MP0/G 0 0.788614f
C888 XB1/XA4/MN1/a_324_334# 0 0.359583f
C889 CK_SAMPLE_BSSW 0 3.70264f
C890 XB1/XA0/MN0/a_324_n18# 0 0.359583f
C891 XB1/M8/a_324_n18# 0 0.356977f
C892 XB1/M8/a_324_334# 0 0.422f
C893 XB1/M6/a_324_n18# 0 0.356977f
C894 XB1/M7/a_324_n18# 0 0.356977f
C895 XB1/XA3/B 0 54.41209f
C896 XB1/XA4/GNG 0 53.065117f
C897 XA0/CEIN 0 19.901903f
C898 XB1/M5/a_324_n18# 0 0.356977f
C899 XB1/M3/a_324_n18# 0 0.356977f
C900 XB1/M4/a_324_n18# 0 0.356977f
C901 XB1/M4/G 0 2.475647f
C902 SAR_IP 0 1.184896f
C903 XB1/M1/a_324_n18# 0 0.422415f
C904 XB1/M2/a_324_n18# 0 0.356977f
C905 XA20/XA9/MN0/a_324_n18# 0 0.360407f
C906 XA20/XA3/CO 0 2.703497f
C907 XA20/XA2/MN6/a_324_334# 0 0.360407f
C908 XA20/XA3a/A 0 2.536943f
C909 XA20/XA3/MN0/a_324_n18# 0 0.360407f
C910 XA20/XA3a/MN0/a_324_n18# 0 0.360407f
C911 XA20/XA4/MN0/a_324_n18# 0 0.360407f
C912 XA20/XA4/MP0/S 0 0.397005f
C913 SARN 0 29.964926f
C914 XA20/XA3/N2 0 0.234927f
C915 XA20/XA9/Y 0 3.176436f
C916 XA20/XA2/N2 0 0.234927f
C917 XA20/XA2/MN0/a_324_n18# 0 0.360407f
C918 XA20/XA3/N1 0 0.905385f
C919 SARP 0 30.549707f
C920 XA20/XA1/MN0/a_324_n18# 0 0.360407f
C921 XA20/XA1/MP0/S 0 0.397005f
C922 XA20/XA9/A 0 3.508213f
C923 XA20/XA0/MN1/a_324_n18# 0 0.422415f
C924 XA20/XA0/MP1/a_216_n18# 0 0.091271f
C925 XA20/XA13/MN1/a_324_n18# 0 0.360407f
C926 XA20/XA13/MN1/a_324_334# 0 0.422f
C927 XA20/XA13/MP1/a_216_334# 0 0.091271f
C928 XA20/XA12/MN0/a_324_n18# 0 0.360407f
C929 XA20/XA11/MN0/a_324_n18# 0 0.360407f
C930 DONE 0 0.902344f
C931 XA20/XA9/MN0/a_324_334# 0 0.360407f
C932 XA20/XA12/Y 0 0.623344f
C933 XA20/XA11/Y 0 0.759612f
C934 XDAC2/XC32a<0>/XRES2/B 0 3.1129f
C935 XDAC2/XC32a<0>/XRES4/B 0 3.516117f
C936 XDAC2/XC32a<0>/XRES8/B 0 3.933522f
C937 XDAC2/XC32a<0>/XRES16/B 0 4.664508f
C938 XDAC2/XC32a<0>/XRES1B/B 0 2.892833f
C939 XDAC2/XC32a<0>/XRES1A/B 0 1.735354f
C940 XDAC2/XC1/XRES2/B 0 3.1129f
C941 XDAC2/XC1/XRES4/B 0 3.516117f
C942 XDAC2/XC1/XRES8/B 0 3.933522f
C943 XDAC2/XC1/XRES16/B 0 4.664508f
C944 XDAC2/XC1/XRES1B/B 0 2.892833f
C945 XDAC2/XC1/XRES1A/B 0 1.735354f
C946 XA0/CN0 0 6.776559f
C947 XDAC2/XC0/XRES2/B 0 3.1129f
C948 XDAC2/XC0/XRES4/B 0 3.516117f
C949 XDAC2/XC0/XRES8/B 0 3.933522f
C950 XDAC2/XC0/XRES16/B 0 4.664508f
C951 XDAC2/XC0/XRES1B/B 0 2.892833f
C952 XDAC2/XC0/XRES1A/B 0 1.735354f
C953 XDAC2/X16ab/XRES2/B 0 3.1129f
C954 XDAC2/X16ab/XRES4/B 0 3.516117f
C955 XDAC2/X16ab/XRES8/B 0 3.933522f
C956 XDAC2/X16ab/XRES16/B 0 4.664508f
C957 XDAC2/X16ab/XRES1B/B 0 2.892833f
C958 XDAC2/X16ab/XRES1A/B 0 1.735354f
C959 XDAC1/XC32a<0>/XRES2/B 0 3.1129f
C960 XDAC1/XC32a<0>/XRES4/B 0 3.516117f
C961 XDAC1/XC32a<0>/XRES8/B 0 3.933522f
C962 XDAC1/XC32a<0>/XRES16/B 0 4.664508f
C963 XDAC1/XC32a<0>/XRES1B/B 0 2.892833f
C964 XDAC1/XC32a<0>/XRES1A/B 0 1.735354f
C965 XDAC1/XC1/XRES2/B 0 3.1129f
C966 XDAC1/XC1/XRES4/B 0 3.516117f
C967 XDAC1/XC1/XRES8/B 0 3.933522f
C968 XDAC1/XC1/XRES16/B 0 4.664508f
C969 XDAC1/XC1/XRES1B/B 0 2.892833f
C970 XDAC1/XC1/XRES1A/B 0 1.735354f
C971 XDAC1/XC0/XRES2/B 0 3.1129f
C972 XDAC1/XC0/XRES4/B 0 3.516117f
C973 XDAC1/XC0/XRES8/B 0 3.933522f
C974 XDAC1/XC0/XRES16/B 0 4.664508f
C975 XDAC1/XC0/XRES1B/B 0 2.892833f
C976 XDAC1/XC0/XRES1A/B 0 1.735354f
C977 D<5> 0 4.36517f
C978 XDAC1/X16ab/XRES2/B 0 3.1129f
C979 XDAC1/X16ab/XRES4/B 0 3.516117f
C980 XDAC1/X16ab/XRES8/B 0 3.933522f
C981 XDAC1/X16ab/XRES16/B 0 4.664508f
C982 XDAC1/X16ab/XRES1B/B 0 2.892833f
C983 XDAC1/X16ab/XRES1A/B 0 1.735354f
C984 XA0/CP1 0 4.930175f
.ends

.subckt SUNSAR_IVTRIX1_CV CN AVDD AVSS MN1/a_324_334# C Y BULKP BULKN MP0/a_216_n18#
+ MP1/a_216_334# A MN0/a_324_n18#
XMP0 MP1/S A AVDD BULKP BULKN MP0/a_216_n18# CN SUNSAR_PCHDL
XMP1 Y CN MP1/S BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 MN1/S A AVSS BULKN MN0/a_324_n18# C SUNSAR_NCHDL
XMN1 Y C MN1/S BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 CN BULKP -0.345553f
C1 AVSS AVDD 0.070034f
C2 BULKP AVDD 0.123213f
C3 BULKP Y 0.069031f
C4 A BULKP -0.231483f
C5 AVDD BULKN 0.259844f
C6 AVSS BULKN 0.395374f
C7 C BULKN 0.372036f
C8 Y BULKN 0.262859f
C9 MN1/a_324_334# BULKN 0.422f
C10 A BULKN 0.569283f
C11 MN0/a_324_n18# BULKN 0.422415f
C12 MP1/a_216_334# BULKN 0.091338f
C13 BULKP BULKN 3.597147f
C14 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_DFQNX1_CV Q QN XA7/C CK D AVDD AVSS
XXA0 AVDD XA0/MN1/a_324_n18# XA1/MN0/a_324_n18# AVSS XA1/MP0/a_216_n18# XA0/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA1 AVDD AVSS XA7/C AVSS XA1/MP0/a_216_n18# XA2/MP0/a_216_n18# AVDD CK XA1/MN0/a_324_n18#
+ XA2/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA2 AVDD AVSS XA6/C AVSS XA2/MP0/a_216_n18# XA3/MP0/a_216_n18# AVDD XA7/C XA2/MN0/a_324_n18#
+ XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA3 XA6/C AVDD AVSS XA4/MN0/a_324_n18# XA7/C XA5/A AVDD AVSS XA3/MP0/a_216_n18# XA4/MP0/a_216_n18#
+ D XA3/MN0/a_324_n18# SUNSAR_IVTRIX1_CV
XXA4 XA7/C AVDD AVSS XA5/MN0/a_324_n18# XA6/C XA5/A AVDD AVSS XA4/MP0/a_216_n18# XA5/MP0/a_216_n18#
+ XA6/A XA4/MN0/a_324_n18# SUNSAR_IVTRIX1_CV
XXA5 AVDD AVSS XA6/A AVSS XA5/MP0/a_216_n18# XA6/MP0/a_216_n18# AVDD XA5/A XA5/MN0/a_324_n18#
+ XA6/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA6 XA7/C AVDD AVSS XA7/MN0/a_324_n18# XA6/C QN AVDD AVSS XA6/MP0/a_216_n18# XA7/MP0/a_216_n18#
+ XA6/A XA6/MN0/a_324_n18# SUNSAR_IVTRIX1_CV
XXA7 XA6/C AVDD AVSS XA8/MN0/a_324_n18# XA7/C QN AVDD AVSS XA7/MP0/a_216_n18# XA8/MP0/a_216_n18#
+ Q XA7/MN0/a_324_n18# SUNSAR_IVTRIX1_CV
XXA8 AVDD AVSS Q AVSS XA8/MP0/a_216_n18# XA8/MP0/a_216_334# AVDD QN XA8/MN0/a_324_n18#
+ XA8/MN0/a_324_334# SUNSAR_IVX1_CV
C0 XA8/MP0/a_216_n18# AVDD -0.312509f
C1 XA5/MP0/a_216_n18# AVDD -0.313035f
C2 XA6/C AVDD 0.894074f
C3 XA7/C XA2/MP0/a_216_n18# 0.066871f
C4 XA3/MP0/a_216_n18# AVDD -0.313035f
C5 AVSS QN 0.208618f
C6 XA7/C CK 0.13667f
C7 XA5/A AVSS 0.31114f
C8 XA6/A AVSS 0.060481f
C9 XA7/C AVSS 0.523585f
C10 XA6/MP0/a_216_n18# AVDD -0.315634f
C11 XA6/C QN 0.060794f
C12 XA5/A XA6/C 0.400241f
C13 XA6/C Q 0.188983f
C14 XA6/A XA6/C 0.511866f
C15 XA6/C D 0.110712f
C16 XA7/C XA6/C 0.555229f
C17 AVDD XA1/MP0/a_216_n18# -0.311986f
C18 AVDD XA4/MP0/a_216_n18# -0.313035f
C19 AVSS XA6/C 0.2601f
C20 XA7/MP0/a_216_n18# AVDD -0.314611f
C21 QN AVDD 0.152707f
C22 XA5/A AVDD 0.149071f
C23 Q AVDD 0.337452f
C24 XA6/A AVDD 0.50597f
C25 XA7/C AVDD 1.562268f
C26 XA2/MP0/a_216_n18# AVDD -0.31496f
C27 Q QN 0.164289f
C28 XA6/A XA5/A 0.225387f
C29 XA7/C QN 0.28651f
C30 XA7/C XA5/A 0.090185f
C31 XA7/C Q 0.128539f
C32 XA7/C XA6/A 0.41755f
C33 XA7/C D 0.117769f
C34 XA7/C 0 2.352415f
C35 QN 0 0.966414f
C36 Q 0 0.838602f
C37 XA8/MN0/a_324_334# 0 0.422f
C38 XA8/MP0/a_216_334# 0 0.091271f
C39 XA8/MN0/a_324_n18# 0 0.360407f
C40 XA7/MN0/a_324_n18# 0 0.360407f
C41 XA6/MN0/a_324_n18# 0 0.360407f
C42 XA5/A 0 0.896691f
C43 XA6/A 0 1.098676f
C44 XA5/MN0/a_324_n18# 0 0.360407f
C45 XA4/MN0/a_324_n18# 0 0.360407f
C46 D 0 0.487386f
C47 XA3/MN0/a_324_n18# 0 0.360407f
C48 XA6/C 0 1.328497f
C49 XA2/MN0/a_324_n18# 0 0.360407f
C50 CK 0 0.515118f
C51 XA1/MN0/a_324_n18# 0 0.360407f
C52 AVSS 0 -0.115052f
C53 XA0/MN1/a_324_n18# 0 0.422415f
C54 AVDD 0 18.699612f
C55 XA0/MP1/a_216_n18# 0 0.091271f
.ends

.subckt SUNSAR_ORX1_CV AVDD AVSS B XA1/MP0/a_216_n18# XA2/A XA1/MN0/a_324_n18# XA2/MP0/a_216_334#
+ A BULKP XA2/MN0/a_324_334# BULKN Y
XXA1 AVDD AVSS XA2/MN0/a_324_n18# B BULKP BULKN XA1/MP0/a_216_n18# XA2/A XA2/MP0/a_216_n18#
+ A XA1/MN0/a_324_n18# SUNSAR_NRX1_CV
XXA2 BULKP AVSS Y BULKN XA2/MP0/a_216_n18# XA2/MP0/a_216_334# AVDD XA2/A XA2/MN0/a_324_n18#
+ XA2/MN0/a_324_334# SUNSAR_IVX1_CV
C0 BULKP XA2/MP0/a_216_n18# -0.310513f
C1 AVSS XA2/A 0.063933f
C2 AVDD XA2/A 0.062592f
C3 B XA2/A 0.110841f
C4 Y BULKN 0.217477f
C5 XA2/MN0/a_324_n18# BULKN 0.357149f
C6 XA2/MN0/a_324_334# BULKN 0.422f
C7 AVDD BULKN 0.321354f
C8 XA2/MP0/a_216_334# BULKN 0.091271f
C9 AVSS BULKN 0.551073f
C10 XA2/A BULKN 0.902459f
C11 XA1/MN0/a_324_n18# BULKN 0.422415f
C12 B BULKN 0.472321f
C13 BULKP BULKN 5.173117f
C14 A BULKN 0.541859f
C15 XA1/MP0/a_216_n18# BULKN 0.091271f
.ends

.subckt SUNSAR_BFX1_CV Y AVDD AVSS MN1/a_324_334# MP1/G A BULKP BULKN MP0/a_216_n18#
+ MP1/a_216_334# MN0/a_324_n18#
XMP0 AVDD A MP1/G BULKP BULKN MP0/a_216_n18# MP1/G SUNSAR_PCHDL
XMP1 Y MP1/G AVDD BULKP BULKN A MP1/a_216_334# SUNSAR_PCHDL
XMN0 AVSS A MP1/G BULKN MN0/a_324_n18# MP1/G SUNSAR_NCHDL
XMN1 Y MP1/G AVSS BULKN A MN1/a_324_334# SUNSAR_NCHDL
C0 MP1/G A 0.120372f
C1 BULKP Y 0.054823f
C2 BULKP AVDD 0.074098f
C3 BULKP A -0.246947f
C4 AVDD AVSS 0.070127f
C5 BULKP MP1/G -0.189656f
C6 MP1/G Y 0.094089f
C7 MP1/G AVSS 0.079416f
C8 AVSS BULKN 0.330762f
C9 Y BULKN 0.213901f
C10 MN1/a_324_334# BULKN 0.422f
C11 AVDD BULKN 0.225252f
C12 MN0/a_324_n18# BULKN 0.422415f
C13 MP1/G BULKN 0.888781f
C14 BULKP BULKN 3.596797f
C15 A BULKN 0.536396f
C16 MP1/a_216_334# BULKN 0.091338f
C17 MP0/a_216_n18# BULKN 0.091338f
.ends

.subckt SUNSAR_ANX1_CV B XA1/MP0/a_216_n18# XA2/A XA1/MN0/a_324_n18# XA2/MP0/a_216_334#
+ A BULKP XA2/MN0/a_324_334# AVDD AVSS BULKN Y XA1/MN1/S
XXA1 XA2/A AVDD AVSS XA2/MN0/a_324_n18# B A BULKP BULKN XA1/MP0/a_216_n18# XA1/MN1/S
+ XA2/MP0/a_216_n18# XA1/MN0/a_324_n18# SUNSAR_NDX1_CV
XXA2 BULKP AVSS Y BULKN XA2/MP0/a_216_n18# XA2/MP0/a_216_334# AVDD XA2/A XA2/MN0/a_324_n18#
+ XA2/MN0/a_324_334# SUNSAR_IVX1_CV
C0 B XA2/A 0.072536f
C1 BULKP XA2/MP0/a_216_n18# -0.310513f
C2 XA2/A AVSS 0.096305f
C3 Y BULKN 0.219919f
C4 XA2/MN0/a_324_n18# BULKN 0.357149f
C5 XA2/MN0/a_324_334# BULKN 0.422f
C6 XA2/MP0/a_216_334# BULKN 0.091271f
C7 AVSS BULKN 0.513075f
C8 AVDD BULKN 0.340245f
C9 XA1/MN0/a_324_n18# BULKN 0.422415f
C10 XA2/A BULKN 0.881652f
C11 B BULKN 0.474447f
C12 BULKP BULKN 5.173112f
C13 A BULKN 0.541856f
C14 XA1/MP0/a_216_n18# BULKN 0.091271f
.ends

.subckt SUNSAR_CAPT8B_CV CKS ENABLE CK_SAMPLE CK_SAMPLE_BSSW EN D<7> D<6> D<5> D<4>
+ D<3> D<2> D<1> D<0> DO<7> DO<6> DO<5> DO<4> DO<3> DO<2> DO<1> DO<0> TIE_L DONE AVSS
+ AVDD
XXD09 DO<5> XD09/QN XD09/XA7/C DONE D<5> AVDD AVSS SUNSAR_DFQNX1_CV
XXB07 DO<7> XB07/QN XB07/XA7/C DONE D<7> AVDD AVSS SUNSAR_DFQNX1_CV
XSUNSAR_IVX1_CV_0 AVDD AVSS XA5/B AVSS XA1/MP1/a_216_334# XA3/MP0/a_216_n18# AVDD
+ ENABLE XA1/MN1/a_324_334# XA3/MN0/a_324_n18# SUNSAR_IVX1_CV
XXI14 DO<0> XI14/QN XI14/XA7/C DONE D<0> AVDD AVSS SUNSAR_DFQNX1_CV
XXG12 DO<2> XG12/QN XG12/XA7/C DONE D<2> AVDD AVSS SUNSAR_DFQNX1_CV
XXE10 DO<4> XE10/QN XE10/XA7/C DONE D<4> AVDD AVSS SUNSAR_DFQNX1_CV
XXC08 DO<6> XC08/QN XC08/XA7/C DONE D<6> AVDD AVSS SUNSAR_DFQNX1_CV
XXA1 AVDD XA1/MN1/a_324_n18# XA1/MN1/a_324_334# AVSS XA1/MP1/a_216_334# XA1/MP1/a_216_n18#
+ SUNSAR_TAPCELLB_CV
XXA2 AVDD AVDD AVSS XA2/MP0/G TIE_L AVSS XA2/MP0/a_216_n18# XA2/MP0/a_216_334# XA2/MN0/a_324_n18#
+ XA2/MN0/a_324_334# SUNSAR_TIEL_CV
XXA5a AVDD AVSS EN AVSS XA5a/MP0/a_216_n18# XA5a/MP0/a_216_334# AVDD CK_SAMPLE XA5a/MN0/a_324_n18#
+ XA5a/MN0/a_324_334# SUNSAR_IVX1_CV
XXA3 AVDD AVSS XA6/B AVSS XA3/MP0/a_216_n18# XA4/MP0/a_216_n18# AVDD XA5/B XA3/MN0/a_324_n18#
+ XA4/MN0/a_324_n18# SUNSAR_IVX1_CV
XXA5 AVDD AVSS XA5/B XA4/MP1/a_216_334# XA5/XA2/A XA4/MN1/a_324_334# XA5a/MP0/a_216_n18#
+ XA6/A AVDD XA5a/MN0/a_324_n18# AVSS CK_SAMPLE SUNSAR_ORX1_CV
XXA4 XA6/A AVDD AVSS XA4/MN1/a_324_334# XA4/MP1/G CKS AVDD AVSS XA4/MP0/a_216_n18#
+ XA4/MP1/a_216_334# XA4/MN0/a_324_n18# SUNSAR_BFX1_CV
XXH13 DO<1> XH13/QN XH13/XA7/C DONE D<1> AVDD AVSS SUNSAR_DFQNX1_CV
XXA6 XA6/B XA5a/MP0/a_216_334# XA6/XA2/A XA5a/MN0/a_324_334# XA2/MP0/a_216_n18# XA6/A
+ AVDD XA2/MN0/a_324_n18# AVDD AVSS AVSS CK_SAMPLE_BSSW XA6/XA1/MN1/S SUNSAR_ANX1_CV
XXF11 DO<3> XF11/QN XF11/XA7/C DONE D<3> AVDD AVSS SUNSAR_DFQNX1_CV
C0 XA6/A CK_SAMPLE 0.103062f
C1 DONE D<3> 0.295113f
C2 DONE D<4> 0.295113f
C3 AVDD DONE 2.494628f
C4 TIE_L AVSS 0.167035f
C5 D<0> AVSS 0.32707f
C6 D<2> XG12/XA7/C 0.159126f
C7 AVDD XA2/MP0/a_216_n18# -0.313603f
C8 XA6/B XA4/MP1/G 0.300066f
C9 AVDD D<2> 0.137402f
C10 XE10/XA7/C XF11/XA7/C 0.060807f
C11 DONE AVSS 7.136208f
C12 AVDD D<5> 0.137402f
C13 XA6/XA2/A EN 0.058309f
C14 D<7> XB07/XA7/C 0.159126f
C15 D<6> XC08/XA7/C 0.159126f
C16 XA6/B XA5/XA2/A 0.134182f
C17 AVDD D<6> 0.137402f
C18 XD09/XA7/C XC08/XA7/C 0.060807f
C19 AVDD CK_SAMPLE 0.496932f
C20 XA6/XA2/A XA2/MP0/G 0.060853f
C21 CK_SAMPLE XA6/B 0.199415f
C22 D<2> AVSS 0.301985f
C23 AVDD XA6/A 0.089821f
C24 D<5> AVSS 0.301985f
C25 XA6/A XA6/B 0.223197f
C26 XB07/XA7/C XC08/XA7/C 0.233892f
C27 AVSS D<6> 0.301985f
C28 AVDD XA1/MP1/a_216_334# -0.311986f
C29 AVDD XA5a/MP0/a_216_334# -0.313603f
C30 CK_SAMPLE AVSS 0.395202f
C31 D<7> AVDD 0.129858f
C32 XA6/A AVSS 0.540389f
C33 D<1> XH13/XA7/C 0.159126f
C34 AVDD ENABLE 0.145509f
C35 AVDD CK_SAMPLE_BSSW 0.508937f
C36 XA5/B XA4/MP1/G 0.138434f
C37 DO<3> AVSS 0.187665f
C38 D<3> D<4> 0.12805f
C39 DONE D<1> 0.295113f
C40 D<7> AVSS 0.290141f
C41 AVDD D<3> 0.137402f
C42 AVDD D<4> 0.137402f
C43 AVDD XA3/MP0/a_216_n18# -0.311309f
C44 ENABLE AVSS 0.410372f
C45 AVDD XA6/B 0.218203f
C46 XA5/B XA5/XA2/A 0.08845f
C47 AVSS DO<1> 0.187666f
C48 AVSS CK_SAMPLE_BSSW 0.339545f
C49 D<2> D<1> 0.12805f
C50 XF11/XA7/C XG12/XA7/C 0.233892f
C51 XA6/A CKS 0.198582f
C52 AVSS D<3> 0.301985f
C53 AVSS D<4> 0.301985f
C54 AVDD XA4/MP0/a_216_n18# -0.311772f
C55 XA6/A XA5/B 0.263519f
C56 AVDD AVSS 6.228554f
C57 XA6/B AVSS 0.54117f
C58 XF11/XA7/C D<3> 0.159126f
C59 DONE D<0> 0.29654f
C60 ENABLE XA5/B 0.10479f
C61 CK_SAMPLE EN 0.28401f
C62 DO<0> AVSS 0.192871f
C63 XA6/B CKS 0.066782f
C64 DO<5> AVSS 0.187665f
C65 AVDD XA5/B 0.083886f
C66 XA5/B XA6/B 0.187691f
C67 DO<7> AVSS 0.186597f
C68 XA6/XA2/A XA6/B 0.172524f
C69 AVDD D<1> 0.137402f
C70 DONE D<2> 0.295113f
C71 CKS AVSS 1.512398f
C72 AVDD XA5a/MP0/a_216_n18# -0.313603f
C73 D<0> XI14/XA7/C 0.159126f
C74 D<5> DONE 0.295113f
C75 XA5/B AVSS 0.356101f
C76 XI14/XA7/C XH13/XA7/C 0.233892f
C77 DONE D<6> 0.295113f
C78 XE10/XA7/C XD09/XA7/C 0.233892f
C79 EN CK_SAMPLE_BSSW 0.080252f
C80 DO<2> AVSS 0.187666f
C81 DO<4> AVSS 0.187665f
C82 XA6/B XA6/XA1/MN1/S 0.057307f
C83 AVDD XA4/MP1/a_216_334# -0.311908f
C84 AVSS D<1> 0.301985f
C85 AVSS DO<6> 0.187666f
C86 AVDD EN 0.458465f
C87 XA6/B EN 0.176334f
C88 D<5> D<6> 0.12805f
C89 XA6/A XA4/MP1/G 0.091672f
C90 XD09/XA7/C D<5> 0.159126f
C91 XG12/XA7/C XH13/XA7/C 0.060806f
C92 D<7> DONE 0.292286f
C93 CK_SAMPLE XA5/XA2/A 0.123914f
C94 EN AVSS 0.334598f
C95 XA5/B CKS 0.210661f
C96 XA6/A XA5/XA2/A 0.06853f
C97 AVDD D<0> 0.142353f
C98 XE10/XA7/C D<4> 0.159127f
C99 XF11/XA7/C 0 2.352415f
C100 XF11/QN 0 0.966414f
C101 DO<3> 0 0.963071f
C102 XF11/XA8/MN0/a_324_334# 0 0.422f
C103 XF11/XA8/MP0/a_216_334# 0 0.091271f
C104 XF11/XA8/MN0/a_324_n18# 0 0.360407f
C105 XF11/XA7/MN0/a_324_n18# 0 0.360407f
C106 XF11/XA6/MN0/a_324_n18# 0 0.360407f
C107 XF11/XA5/A 0 0.896691f
C108 XF11/XA6/A 0 1.098676f
C109 XF11/XA5/MN0/a_324_n18# 0 0.360407f
C110 XF11/XA4/MN0/a_324_n18# 0 0.360407f
C111 D<3> 0 0.918631f
C112 XF11/XA3/MN0/a_324_n18# 0 0.360407f
C113 XF11/XA6/C 0 1.328497f
C114 XF11/XA2/MN0/a_324_n18# 0 0.360407f
C115 XF11/XA1/MN0/a_324_n18# 0 0.360407f
C116 XF11/XA0/MN1/a_324_n18# 0 0.422415f
C117 XF11/XA0/MP1/a_216_n18# 0 0.091271f
C118 CK_SAMPLE_BSSW 0 0.351307f
C119 XA6/XA2/MN0/a_324_n18# 0 0.360407f
C120 XA2/MN0/a_324_n18# 0 0.359492f
C121 XA5a/MN0/a_324_334# 0 0.359492f
C122 XA6/XA2/A 0 0.871363f
C123 XA6/B 0 1.026141f
C124 XH13/XA7/C 0 2.352415f
C125 XH13/QN 0 0.966414f
C126 DO<1> 0 0.963071f
C127 XH13/XA8/MN0/a_324_334# 0 0.422f
C128 XH13/XA8/MP0/a_216_334# 0 0.091271f
C129 XH13/XA8/MN0/a_324_n18# 0 0.360407f
C130 XH13/XA7/MN0/a_324_n18# 0 0.360407f
C131 XH13/XA6/MN0/a_324_n18# 0 0.360407f
C132 XH13/XA5/A 0 0.896691f
C133 XH13/XA6/A 0 1.098676f
C134 XH13/XA5/MN0/a_324_n18# 0 0.360407f
C135 XH13/XA4/MN0/a_324_n18# 0 0.360407f
C136 D<1> 0 0.918631f
C137 XH13/XA3/MN0/a_324_n18# 0 0.360407f
C138 XH13/XA6/C 0 1.328497f
C139 XH13/XA2/MN0/a_324_n18# 0 0.360407f
C140 XH13/XA1/MN0/a_324_n18# 0 0.360407f
C141 XH13/XA0/MN1/a_324_n18# 0 0.422415f
C142 XH13/XA0/MP1/a_216_n18# 0 0.091271f
C143 XA4/MP1/G 0 0.884568f
C144 CKS 0 0.801993f
C145 CK_SAMPLE 0 0.805485f
C146 XA5/XA2/MN0/a_324_n18# 0 0.360407f
C147 XA5a/MN0/a_324_n18# 0 0.359492f
C148 XA5/XA2/A 0 0.888056f
C149 XA4/MN1/a_324_334# 0 0.359492f
C150 XA5/B 0 1.456308f
C151 XA6/A 0 1.690748f
C152 XA3/MN0/a_324_n18# 0 0.359492f
C153 XA4/MN0/a_324_n18# 0 0.359492f
C154 EN 0 0.153136f
C155 XA2/MP0/G 0 0.708335f
C156 TIE_L 0 0.1839f
C157 XA2/MN0/a_324_334# 0 0.422f
C158 XA2/MP0/a_216_334# 0 0.091271f
C159 XA1/MN1/a_324_n18# 0 0.422415f
C160 XA1/MP1/a_216_n18# 0 0.091271f
C161 XC08/XA7/C 0 2.352415f
C162 XC08/QN 0 0.966414f
C163 DO<6> 0 0.963071f
C164 XC08/XA8/MN0/a_324_334# 0 0.422f
C165 XC08/XA8/MP0/a_216_334# 0 0.091271f
C166 XC08/XA8/MN0/a_324_n18# 0 0.360407f
C167 XC08/XA7/MN0/a_324_n18# 0 0.360407f
C168 XC08/XA6/MN0/a_324_n18# 0 0.360407f
C169 XC08/XA5/A 0 0.896691f
C170 XC08/XA6/A 0 1.098676f
C171 XC08/XA5/MN0/a_324_n18# 0 0.360407f
C172 XC08/XA4/MN0/a_324_n18# 0 0.360407f
C173 D<6> 0 0.918631f
C174 XC08/XA3/MN0/a_324_n18# 0 0.360407f
C175 XC08/XA6/C 0 1.328497f
C176 XC08/XA2/MN0/a_324_n18# 0 0.360407f
C177 XC08/XA1/MN0/a_324_n18# 0 0.360407f
C178 AVSS 0 -8.464533f
C179 XC08/XA0/MN1/a_324_n18# 0 0.422415f
C180 AVDD 0 0.152305p
C181 XC08/XA0/MP1/a_216_n18# 0 0.091271f
C182 XE10/XA7/C 0 2.352415f
C183 XE10/QN 0 0.966414f
C184 DO<4> 0 0.963071f
C185 XE10/XA8/MN0/a_324_334# 0 0.422f
C186 XE10/XA8/MP0/a_216_334# 0 0.091271f
C187 XE10/XA8/MN0/a_324_n18# 0 0.360407f
C188 XE10/XA7/MN0/a_324_n18# 0 0.360407f
C189 XE10/XA6/MN0/a_324_n18# 0 0.360407f
C190 XE10/XA5/A 0 0.896691f
C191 XE10/XA6/A 0 1.098676f
C192 XE10/XA5/MN0/a_324_n18# 0 0.360407f
C193 XE10/XA4/MN0/a_324_n18# 0 0.360407f
C194 D<4> 0 0.918631f
C195 XE10/XA3/MN0/a_324_n18# 0 0.360407f
C196 XE10/XA6/C 0 1.328497f
C197 XE10/XA2/MN0/a_324_n18# 0 0.360407f
C198 XE10/XA1/MN0/a_324_n18# 0 0.360407f
C199 XE10/XA0/MN1/a_324_n18# 0 0.422415f
C200 XE10/XA0/MP1/a_216_n18# 0 0.091271f
C201 XG12/XA7/C 0 2.352415f
C202 XG12/QN 0 0.966414f
C203 DO<2> 0 0.963071f
C204 XG12/XA8/MN0/a_324_334# 0 0.422f
C205 XG12/XA8/MP0/a_216_334# 0 0.091271f
C206 XG12/XA8/MN0/a_324_n18# 0 0.360407f
C207 XG12/XA7/MN0/a_324_n18# 0 0.360407f
C208 XG12/XA6/MN0/a_324_n18# 0 0.360407f
C209 XG12/XA5/A 0 0.896691f
C210 XG12/XA6/A 0 1.098676f
C211 XG12/XA5/MN0/a_324_n18# 0 0.360407f
C212 XG12/XA4/MN0/a_324_n18# 0 0.360407f
C213 D<2> 0 0.918631f
C214 XG12/XA3/MN0/a_324_n18# 0 0.360407f
C215 XG12/XA6/C 0 1.328497f
C216 XG12/XA2/MN0/a_324_n18# 0 0.360407f
C217 XG12/XA1/MN0/a_324_n18# 0 0.360407f
C218 XG12/XA0/MN1/a_324_n18# 0 0.422415f
C219 XG12/XA0/MP1/a_216_n18# 0 0.091271f
C220 XI14/XA7/C 0 2.352415f
C221 XI14/QN 0 0.966414f
C222 DO<0> 0 0.960285f
C223 XI14/XA8/MN0/a_324_334# 0 0.422f
C224 XI14/XA8/MP0/a_216_334# 0 0.091271f
C225 XI14/XA8/MN0/a_324_n18# 0 0.360407f
C226 XI14/XA7/MN0/a_324_n18# 0 0.360407f
C227 XI14/XA6/MN0/a_324_n18# 0 0.360407f
C228 XI14/XA5/A 0 0.896691f
C229 XI14/XA6/A 0 1.098676f
C230 XI14/XA5/MN0/a_324_n18# 0 0.360407f
C231 XI14/XA4/MN0/a_324_n18# 0 0.360407f
C232 D<0> 0 1.011141f
C233 XI14/XA3/MN0/a_324_n18# 0 0.360407f
C234 XI14/XA6/C 0 1.328497f
C235 XI14/XA2/MN0/a_324_n18# 0 0.360407f
C236 XI14/XA1/MN0/a_324_n18# 0 0.360407f
C237 XI14/XA0/MN1/a_324_n18# 0 0.422415f
C238 XI14/XA0/MP1/a_216_n18# 0 0.091271f
C239 ENABLE 0 0.918187f
C240 XA1/MN1/a_324_334# 0 0.359492f
C241 XB07/XA7/C 0 2.352415f
C242 XB07/QN 0 0.966414f
C243 DO<7> 0 0.973878f
C244 XB07/XA8/MN0/a_324_334# 0 0.422f
C245 XB07/XA8/MP0/a_216_334# 0 0.091271f
C246 XB07/XA8/MN0/a_324_n18# 0 0.360407f
C247 XB07/XA7/MN0/a_324_n18# 0 0.360407f
C248 XB07/XA6/MN0/a_324_n18# 0 0.360407f
C249 XB07/XA5/A 0 0.896691f
C250 XB07/XA6/A 0 1.098676f
C251 XB07/XA5/MN0/a_324_n18# 0 0.360407f
C252 XB07/XA4/MN0/a_324_n18# 0 0.360407f
C253 D<7> 0 1.10231f
C254 XB07/XA3/MN0/a_324_n18# 0 0.360407f
C255 XB07/XA6/C 0 1.328497f
C256 XB07/XA2/MN0/a_324_n18# 0 0.360407f
C257 DONE 0 9.575078f
C258 XB07/XA1/MN0/a_324_n18# 0 0.360407f
C259 XB07/XA0/MN1/a_324_n18# 0 0.422415f
C260 XB07/XA0/MP1/a_216_n18# 0 0.091271f
C261 XD09/XA7/C 0 2.352415f
C262 XD09/QN 0 0.966414f
C263 DO<5> 0 0.965307f
C264 XD09/XA8/MN0/a_324_334# 0 0.422f
C265 XD09/XA8/MP0/a_216_334# 0 0.091271f
C266 XD09/XA8/MN0/a_324_n18# 0 0.360407f
C267 XD09/XA7/MN0/a_324_n18# 0 0.360407f
C268 XD09/XA6/MN0/a_324_n18# 0 0.360407f
C269 XD09/XA5/A 0 0.896691f
C270 XD09/XA6/A 0 1.098676f
C271 XD09/XA5/MN0/a_324_n18# 0 0.360407f
C272 XD09/XA4/MN0/a_324_n18# 0 0.360407f
C273 D<5> 0 0.918631f
C274 XD09/XA3/MN0/a_324_n18# 0 0.360407f
C275 XD09/XA6/C 0 1.328497f
C276 XD09/XA2/MN0/a_324_n18# 0 0.360407f
C277 XD09/XA1/MN0/a_324_n18# 0 0.360407f
C278 XD09/XA0/MN1/a_324_n18# 0 0.422415f
C279 XD09/XA0/MP1/a_216_n18# 0 0.091271f
.ends

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5]
*+ ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7]
*+ uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
*+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
*+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
*+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
*+ VPWR VGND
XTT06SAR_NDIO_0 VGND clk TT06SAR_NDIO
XTT06SAR_NDIO_1 VGND SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW TT06SAR_NDIO
XTT06SAR_NDIO_2 VGND ui_in[0] TT06SAR_NDIO
Xtt_um_TT06_SAR_done_0 SUNSAR_SAR8B_CV_0/DONE uio_out[0] uio_oe[0] VPWR VGND tt_um_TT06_SAR_done
Xsky130_fd_pr__cap_mim_m3_1_XS736D_0 VPWR VGND VGND sky130_fd_pr__cap_mim_m3_1_XS736D
XSUNSAR_SAR8B_CV_0 ua[1] ua[0] SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/D<4>
+ SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/XA3/CEO SUNSAR_SAR8B_CV_0/XA6/CN0
+ SUNSAR_SAR8B_CV_0/XA6/CP0 SUNSAR_SAR8B_CV_0/XA3/CN0 SUNSAR_SAR8B_CV_0/XA20/XA9/A
+ SUNSAR_SAR8B_CV_0/XA3/CP0 SUNSAR_SAR8B_CV_0/XA4/DONE SUNSAR_SAR8B_CV_0/XA0/XA9/B
+ SUNSAR_SAR8B_CV_0/XA7/CEO SUNSAR_SAR8B_CV_0/XA0/CP0 SUNSAR_SAR8B_CV_0/XA4/CEO SUNSAR_SAR8B_CV_0/XA7/CN0
+ SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/XA1/CEO SUNSAR_SAR8B_CV_0/XA7/CP0 SUNSAR_SAR8B_CV_0/XA4/CN0
+ SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA0/CEIN SUNSAR_SAR8B_CV_0/XA4/CP0 SUNSAR_SAR8B_CV_0/XA1/CN0
+ SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA2/DONE SUNSAR_SAR8B_CV_0/XA1/CP0 SUNSAR_SAR8B_CV_0/XA5/CEO
+ SUNSAR_SAR8B_CV_0/XA20/XA4/MP0/S SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/XA2/CEO
+ SUNSAR_SAR8B_CV_0/SARP SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0/XA5/CN0
+ SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA0/CEO SUNSAR_SAR8B_CV_0/XA5/CP0 SUNSAR_SAR8B_CV_0/XA6/DONE
+ SUNSAR_SAR8B_CV_0/XA0/XA4/A SUNSAR_SAR8B_CV_0/XA2/CN0 SUNSAR_SAR8B_CV_0/D<5> VPWR
+ SUNSAR_SAR8B_CV_0/XA2/CP0 SUNSAR_SAR8B_CV_0/SARN VPWR SUNSAR_SAR8B_CV_0/XA6/CEO
+ VGND SUNSAR_SAR8B_CV
XSUNSAR_CAPT8B_CV_0 clk ui_in[0] SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW
+ SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/D<5>
+ SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/D<1>
+ SUNSAR_SAR8B_CV_0/D<0> uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2]
+ uo_out[1] uo_out[0] TIE_L SUNSAR_SAR8B_CV_0/DONE VGND VPWR SUNSAR_CAPT8B_CV
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R1 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R2 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R3 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R4 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R5 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R6 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R7 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R8 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R9 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R10 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R11 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R12 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R13 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R14 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R15 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
C0 uo_out[4] uio_oe[0] 0.550054f
C1 TIE_L1 uo_out[5] 0.275794f
C2 VPWR TIE_L 0.370965f
C3 VGND SUNSAR_SAR8B_CV_0/D<2> 3.643656f
C4 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW ui_in[0] 0.097118f
C5 TIE_L uo_out[4] 0.31941f
C6 SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/XA3/XA9/B 0.058103f
C7 VGND SUNSAR_SAR8B_CV_0/XA1/CP0 -0.221564f
C8 SUNSAR_SAR8B_CV_0/XA3/CEO SUNSAR_SAR8B_CV_0/D<4> 0.05126f
C9 VGND SUNSAR_SAR8B_CV_0/DONE 1.348305f
C10 VGND uo_out[6] 0.199834f
C11 VGND SUNSAR_SAR8B_CV_0/XA1/CN0 -0.15266f
C12 SUNSAR_SAR8B_CV_0/XA0/XA4/A SUNSAR_SAR8B_CV_0/D<7> 0.103251f
C13 uo_out[7] uio_out[0] 0.07272f
C14 SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/D<0> 0.315767f
C15 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW uio_oe[0] 0.135493f
C16 VGND VPWR 24.268234f
C17 uo_out[6] uo_out[5] 0.318994f
C18 uio_oe[0] uio_out[0] 1.555271f
C19 SUNSAR_SAR8B_CV_0/XA20/XA9/A SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.09352f
C20 TIE_L uio_out[0] 0.44106f
C21 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA5/XA9/B 0.058103f
C22 uo_out[2] uo_out[1] 0.060561f
C23 SUNSAR_SAR8B_CV_0/XA5/CP0 SUNSAR_SAR8B_CV_0/D<2> 0.151875f
C24 ua[1] SUNSAR_SAR8B_CV_0/XA0/CEIN 0.312742f
C25 uo_out[4] uo_out[5] 1.133807f
C26 VPWR SUNSAR_SAR8B_CV_0/D<4> 1.689756f
C27 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA5/CEO 0.05126f
C28 VGND SUNSAR_SAR8B_CV_0/D<5> 3.751857f
C29 uo_out[1] uo_out[0] 0.328349f
C30 SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/XA7/XA9/B 0.058103f
C31 SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/D<0> 0.193713f
C32 SUNSAR_SAR8B_CV_0/XA5/CN0 SUNSAR_SAR8B_CV_0/D<2> 0.411523f
C33 SUNSAR_SAR8B_CV_0/XA0/CEIN ua[0] 0.982813f
C34 SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.494615f
C35 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW VGND 3.243993f
C36 VGND uio_out[0] 0.384239f
C37 VPWR SUNSAR_SAR8B_CV_0/D<0> 1.952988f
C38 VGND SUNSAR_SAR8B_CV_0/D<1> 3.727024f
C39 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<2> 0.074477f
C40 uio_out[0] uo_out[5] 0.109219f
C41 VGND SUNSAR_SAR8B_CV_0/D<6> 3.637564f
C42 VPWR clk 0.185197f
C43 SUNSAR_SAR8B_CV_0/XA2/CP0 SUNSAR_SAR8B_CV_0/D<5> 0.477434f
C44 VPWR SUNSAR_SAR8B_CV_0/D<3> 1.692954f
C45 SUNSAR_SAR8B_CV_0/XA2/CN0 SUNSAR_SAR8B_CV_0/D<5> 0.251493f
C46 VGND SUNSAR_SAR8B_CV_0/XA6/CN0 -0.260744f
C47 SUNSAR_SAR8B_CV_0/DONE SUNSAR_SAR8B_CV_0/XA7/CEO 0.123345f
C48 VPWR SUNSAR_SAR8B_CV_0/D<7> 0.570534f
C49 uo_out[7] uio_oe[0] 0.43252f
C50 SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/XA6/CP0 0.151117f
C51 TIE_L uo_out[7] 0.471918f
C52 uo_out[1] uio_out[0] 0.064738f
C53 SUNSAR_SAR8B_CV_0/XA2/CEO SUNSAR_SAR8B_CV_0/D<4> 0.075193f
C54 VPWR SUNSAR_SAR8B_CV_0/CK_SAMPLE 2.139971f
C55 SUNSAR_CAPT8B_CV_0/XA2/MP0/G uio_oe[0] 0.064035f
C56 SUNSAR_SAR8B_CV_0/XA0/CEIN VPWR 1.427229f
C57 TIE_L uio_oe[0] 1.219126f
C58 ua[1] ua[0] 3.839995f
C59 VGND ui_in[0] 0.595812f
C60 clk uio_out[0] 0.120689f
C61 VGND SUNSAR_SAR8B_CV_0/XA4/CP0 -0.063096f
C62 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<5> 0.073932f
C63 uo_out[2] uo_out[3] 0.08287f
C64 VGND SUNSAR_SAR8B_CV_0/XA4/CN0 -0.260744f
C65 SUNSAR_SAR8B_CV_0/XA0/CEO SUNSAR_SAR8B_CV_0/D<6> 0.075193f
C66 VGND uo_out[7] 0.057608f
C67 SUNSAR_SAR8B_CV_0/XA6/CEO SUNSAR_SAR8B_CV_0/D<0> 0.07415f
C68 VGND uio_oe[0] 0.366251f
C69 SUNSAR_SAR8B_CV_0/XA20/XA4/MP0/S SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.061422f
C70 uo_out[7] uo_out[5] 1.578182f
C71 VGND TIE_L 0.100247f
C72 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/DONE 0.054848f
C73 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<1> 0.073932f
C74 VPWR uo_out[3] 0.234367f
C75 uo_out[4] uo_out[3] 0.846609f
C76 uio_oe[0] uo_out[5] 1.553295f
C77 ua[1] VPWR 0.257135f
C78 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<6> 0.074477f
C79 VGND SUNSAR_SAR8B_CV_0/XA3/CN0 -0.26062f
C80 TIE_L uo_out[5] 1.309194f
C81 SUNSAR_SAR8B_CV_0/XA1/CEO SUNSAR_SAR8B_CV_0/D<6> 0.05126f
C82 SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/DONE 0.131506f
C83 SUNSAR_SAR8B_CV_0/XA0/XA9/B SUNSAR_SAR8B_CV_0/D<7> 0.082644f
C84 clk ui_in[0] 0.217403f
C85 SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA1/XA9/B 0.058103f
C86 VPWR ua[0] 0.537238f
C87 VPWR TIE_L1 0.114647f
C88 VPWR SUNSAR_SAR8B_CV_0/EN 7.947423f
C89 uo_out[1] uio_oe[0] 0.432143f
C90 SUNSAR_SAR8B_CV_0/XA3/CN0 SUNSAR_SAR8B_CV_0/D<4> 0.411522f
C91 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/CP0 0.151117f
C92 SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/XA6/DONE 0.054848f
C93 SUNSAR_SAR8B_CV_0/D<0> SUNSAR_SAR8B_CV_0/XA7/CN0 0.08663f
C94 TIE_L uo_out[1] 0.50141f
C95 SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/XA0/CP0 0.068981f
C96 VGND SUNSAR_SAR8B_CV_0/XA3/CP0 -0.062957f
C97 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/CN0 0.410141f
C98 uo_out[3] uio_out[0] 0.057862f
C99 VPWR SUNSAR_SAR8B_CV_0/D<2> 1.705346f
C100 ua[1] SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0.221633f
C101 ui_in[0] SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.079428f
C102 clk uio_oe[0] 0.260056f
C103 VGND SUNSAR_SAR8B_CV_0/D<4> 3.598254f
C104 TIE_L clk 0.13612f
C105 SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/XA3/CP0 0.151875f
C106 VPWR SUNSAR_SAR8B_CV_0/DONE 0.952355f
C107 VGND SUNSAR_SAR8B_CV_0/XA6/CP0 -0.063096f
C108 VPWR uo_out[6] 0.323007f
C109 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW ua[0] 0.437286f
C110 SUNSAR_SAR8B_CV_0/SARN SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.077154f
C111 VGND SUNSAR_SAR8B_CV_0/XA2/CP0 -0.222661f
C112 uo_out[4] uo_out[6] 0.843602f
C113 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0/EN 0.147251f
C114 VGND SUNSAR_SAR8B_CV_0/XA2/CN0 -0.152784f
C115 VGND SUNSAR_SAR8B_CV_0/D<0> 3.041315f
C116 VGND SUNSAR_SAR8B_CV_0/XA5/CP0 -0.062957f
C117 TIE_L2 VPWR 0.09991f
C118 VGND clk 0.197311f
C119 uo_out[2] uio_out[0] 0.052955f
C120 VGND SUNSAR_SAR8B_CV_0/D<3> 3.719566f
C121 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/XA4/CEO 0.075193f
C122 SUNSAR_SAR8B_CV_0/D<2> SUNSAR_SAR8B_CV_0/D<1> 0.050961f
C123 VGND SUNSAR_SAR8B_CV_0/XA5/CN0 -0.26062f
C124 VPWR SUNSAR_SAR8B_CV_0/D<5> 1.686887f
C125 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0/DONE 0.094851f
C126 uo_out[0] uio_out[0] 0.201579f
C127 SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/XA6/CEO 0.075291f
C128 VGND SUNSAR_SAR8B_CV_0/D<7> 1.927649f
C129 SUNSAR_SAR8B_CV_0/D<4> SUNSAR_SAR8B_CV_0/D<3> 0.054939f
C130 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW VPWR 0.168521f
C131 VGND SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.679423f
C132 SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA1/CP0 0.476574f
C133 VPWR uio_out[0] 0.145655f
C134 SUNSAR_SAR8B_CV_0/D<6> SUNSAR_SAR8B_CV_0/XA1/CN0 0.252238f
C135 SUNSAR_SAR8B_CV_0/EN ui_in[0] 0.968121f
C136 uo_out[3] uio_oe[0] 0.21235f
C137 VPWR SUNSAR_SAR8B_CV_0/D<1> 1.714778f
C138 TIE_L uo_out[3] 0.185334f
C139 VGND SUNSAR_SAR8B_CV_0/XA7/CP0 -0.065363f
C140 VPWR SUNSAR_SAR8B_CV_0/D<6> 1.725454f
C141 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<4> 0.074477f
C142 TIE_L1 uo_out[7] 0.206895f
C143 SUNSAR_SAR8B_CV_0/SARP SUNSAR_SAR8B_CV_0/SARN 0.059854f
C144 TIE_L1 uio_oe[0] 0.902557f
C145 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW uio_out[0] 0.088825f
C146 TIE_L TIE_L1 0.257793f
C147 ui_in[0] SUNSAR_SAR8B_CV_0/DONE 0.159434f
C148 SUNSAR_SAR8B_CV_0/XA7/CEO SUNSAR_SAR8B_CV_0/D<0> 0.075015f
C149 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<0> 0.075213f
C150 ua[1] VGND 0.26469f
C151 VPWR ui_in[0] 1.386636f
C152 SUNSAR_SAR8B_CV_0/D<1> SUNSAR_SAR8B_CV_0/XA6/XA9/B 0.058072f
C153 uo_out[2] uio_oe[0] 0.267753f
C154 SUNSAR_SAR8B_CV_0/XA2/XA9/B SUNSAR_SAR8B_CV_0/D<5> 0.058072f
C155 SUNSAR_SAR8B_CV_0/CK_SAMPLE SUNSAR_SAR8B_CV_0/D<3> 0.073932f
C156 uo_out[6] uo_out[7] 2.362091f
C157 SUNSAR_SAR8B_CV_0/XA7/CP0 SUNSAR_SAR8B_CV_0/D<0> 0.155245f
C158 uo_out[2] TIE_L 0.156661f
C159 SUNSAR_SAR8B_CV_0/EN SUNSAR_SAR8B_CV_0/XA7/XA2/A 0.050875f
C160 uo_out[0] uio_oe[0] 0.670799f
C161 SUNSAR_SAR8B_CV_0/D<3> SUNSAR_SAR8B_CV_0/XA4/XA9/B 0.058072f
C162 uo_out[6] uio_oe[0] 0.057603f
C163 TIE_L uo_out[0] 0.278654f
C164 VGND ua[0] 0.823969f
C165 SUNSAR_SAR8B_CV_0/D<7> SUNSAR_SAR8B_CV_0/CK_SAMPLE 0.174845f
C166 SUNSAR_SAR8B_CV_0/XA6/CN0 SUNSAR_SAR8B_CV_0/D<1> 0.410141f
C167 VPWR uo_out[7] 0.253367f
C168 SUNSAR_SAR8B_CV_0/XA0/CEIN SUNSAR_SAR8B_CV_0/D<7> 0.093457f
C169 VGND SUNSAR_SAR8B_CV_0/EN 0.497831f
C170 TIE_L uo_out[6] 0.204625f
C171 uo_out[4] uo_out[7] 0.121648f
C172 SUNSAR_SAR8B_CV_0/XA2/DONE SUNSAR_SAR8B_CV_0/D<5> 0.054848f
C173 TIE_L2 uo_out[7] 0.100011f
C174 VPWR uio_oe[0] 1.039709f
C175 ua[2] 0 0.119794f
C176 ua[3] 0 0.119794f
C177 ua[4] 0 0.121038f
C178 ua[5] 0 0.122428f
C179 ua[6] 0 0.122428f
C180 ua[7] 0 0.111009f
C181 ena 0 0.073297f
C182 uio_oe[7] 0 0.062293f
C183 TIE_L1 0 1.51307f
C184 TIE_L2 0 1.83212f
C185 m1_14848_7490# 0 0.145721f $ **FLOATING
C186 SUNSAR_CAPT8B_CV_0/XF11/XA7/C 0 2.352415f
C187 SUNSAR_CAPT8B_CV_0/XF11/QN 0 0.966414f
C188 uo_out[3] 0 1.33751f
C189 SUNSAR_CAPT8B_CV_0/XF11/XA8/MN0/a_324_334# 0 0.422f
C190 SUNSAR_CAPT8B_CV_0/XF11/XA8/MP0/a_216_334# 0 0.091271f
C191 SUNSAR_CAPT8B_CV_0/XF11/XA8/MN0/a_324_n18# 0 0.360407f
C192 SUNSAR_CAPT8B_CV_0/XF11/XA7/MN0/a_324_n18# 0 0.360407f
C193 SUNSAR_CAPT8B_CV_0/XF11/XA6/MN0/a_324_n18# 0 0.360407f
C194 SUNSAR_CAPT8B_CV_0/XF11/XA5/A 0 0.896691f
C195 SUNSAR_CAPT8B_CV_0/XF11/XA6/A 0 1.098676f
C196 SUNSAR_CAPT8B_CV_0/XF11/XA5/MN0/a_324_n18# 0 0.360407f
C197 SUNSAR_CAPT8B_CV_0/XF11/XA4/MN0/a_324_n18# 0 0.360407f
C198 SUNSAR_CAPT8B_CV_0/XF11/XA3/MN0/a_324_n18# 0 0.360407f
C199 SUNSAR_CAPT8B_CV_0/XF11/XA6/C 0 1.328497f
C200 SUNSAR_CAPT8B_CV_0/XF11/XA2/MN0/a_324_n18# 0 0.360407f
C201 SUNSAR_CAPT8B_CV_0/XF11/XA1/MN0/a_324_n18# 0 0.360407f
C202 SUNSAR_CAPT8B_CV_0/XF11/XA0/MN1/a_324_n18# 0 0.422415f
C203 SUNSAR_CAPT8B_CV_0/XF11/XA0/MP1/a_216_n18# 0 0.091271f
C204 SUNSAR_CAPT8B_CV_0/XA6/XA2/MN0/a_324_n18# 0 0.360407f
C205 SUNSAR_CAPT8B_CV_0/XA2/MN0/a_324_n18# 0 0.359492f
C206 SUNSAR_CAPT8B_CV_0/XA5a/MN0/a_324_334# 0 0.359492f
C207 SUNSAR_CAPT8B_CV_0/XA6/XA2/A 0 0.871363f
C208 SUNSAR_CAPT8B_CV_0/XA6/B 0 1.026141f
C209 SUNSAR_CAPT8B_CV_0/XH13/XA7/C 0 2.352415f
C210 SUNSAR_CAPT8B_CV_0/XH13/QN 0 0.966414f
C211 uo_out[1] 0 1.194172f
C212 SUNSAR_CAPT8B_CV_0/XH13/XA8/MN0/a_324_334# 0 0.422f
C213 SUNSAR_CAPT8B_CV_0/XH13/XA8/MP0/a_216_334# 0 0.091271f
C214 SUNSAR_CAPT8B_CV_0/XH13/XA8/MN0/a_324_n18# 0 0.360407f
C215 SUNSAR_CAPT8B_CV_0/XH13/XA7/MN0/a_324_n18# 0 0.360407f
C216 SUNSAR_CAPT8B_CV_0/XH13/XA6/MN0/a_324_n18# 0 0.360407f
C217 SUNSAR_CAPT8B_CV_0/XH13/XA5/A 0 0.896691f
C218 SUNSAR_CAPT8B_CV_0/XH13/XA6/A 0 1.098676f
C219 SUNSAR_CAPT8B_CV_0/XH13/XA5/MN0/a_324_n18# 0 0.360407f
C220 SUNSAR_CAPT8B_CV_0/XH13/XA4/MN0/a_324_n18# 0 0.360407f
C221 SUNSAR_CAPT8B_CV_0/XH13/XA3/MN0/a_324_n18# 0 0.360407f
C222 SUNSAR_CAPT8B_CV_0/XH13/XA6/C 0 1.328497f
C223 SUNSAR_CAPT8B_CV_0/XH13/XA2/MN0/a_324_n18# 0 0.360407f
C224 SUNSAR_CAPT8B_CV_0/XH13/XA1/MN0/a_324_n18# 0 0.360407f
C225 SUNSAR_CAPT8B_CV_0/XH13/XA0/MN1/a_324_n18# 0 0.422415f
C226 SUNSAR_CAPT8B_CV_0/XH13/XA0/MP1/a_216_n18# 0 0.091271f
C227 SUNSAR_CAPT8B_CV_0/XA4/MP1/G 0 0.884568f
C228 clk 0 3.641592f
C229 SUNSAR_CAPT8B_CV_0/XA5/XA2/MN0/a_324_n18# 0 0.360407f
C230 SUNSAR_CAPT8B_CV_0/XA5a/MN0/a_324_n18# 0 0.359492f
C231 SUNSAR_CAPT8B_CV_0/XA5/XA2/A 0 0.888056f
C232 SUNSAR_CAPT8B_CV_0/XA4/MN1/a_324_334# 0 0.359492f
C233 SUNSAR_CAPT8B_CV_0/XA5/B 0 1.456308f
C234 SUNSAR_CAPT8B_CV_0/XA6/A 0 1.690748f
C235 SUNSAR_CAPT8B_CV_0/XA3/MN0/a_324_n18# 0 0.359492f
C236 SUNSAR_CAPT8B_CV_0/XA4/MN0/a_324_n18# 0 0.359492f
C237 SUNSAR_CAPT8B_CV_0/XA2/MP0/G 0 0.708335f
C238 TIE_L 0 0.99989f
C239 SUNSAR_CAPT8B_CV_0/XA2/MN0/a_324_334# 0 0.422f
C240 SUNSAR_CAPT8B_CV_0/XA2/MP0/a_216_334# 0 0.091271f
C241 SUNSAR_CAPT8B_CV_0/XA1/MN1/a_324_n18# 0 0.422415f
C242 SUNSAR_CAPT8B_CV_0/XA1/MP1/a_216_n18# 0 0.091271f
C243 SUNSAR_CAPT8B_CV_0/XC08/XA7/C 0 2.352415f
C244 SUNSAR_CAPT8B_CV_0/XC08/QN 0 0.966414f
C245 uo_out[6] 0 1.372751f
C246 SUNSAR_CAPT8B_CV_0/XC08/XA8/MN0/a_324_334# 0 0.422f
C247 SUNSAR_CAPT8B_CV_0/XC08/XA8/MP0/a_216_334# 0 0.091271f
C248 SUNSAR_CAPT8B_CV_0/XC08/XA8/MN0/a_324_n18# 0 0.360407f
C249 SUNSAR_CAPT8B_CV_0/XC08/XA7/MN0/a_324_n18# 0 0.360407f
C250 SUNSAR_CAPT8B_CV_0/XC08/XA6/MN0/a_324_n18# 0 0.360407f
C251 SUNSAR_CAPT8B_CV_0/XC08/XA5/A 0 0.896691f
C252 SUNSAR_CAPT8B_CV_0/XC08/XA6/A 0 1.098676f
C253 SUNSAR_CAPT8B_CV_0/XC08/XA5/MN0/a_324_n18# 0 0.360407f
C254 SUNSAR_CAPT8B_CV_0/XC08/XA4/MN0/a_324_n18# 0 0.360407f
C255 SUNSAR_CAPT8B_CV_0/XC08/XA3/MN0/a_324_n18# 0 0.360407f
C256 SUNSAR_CAPT8B_CV_0/XC08/XA6/C 0 1.328497f
C257 SUNSAR_CAPT8B_CV_0/XC08/XA2/MN0/a_324_n18# 0 0.360407f
C258 SUNSAR_CAPT8B_CV_0/XC08/XA1/MN0/a_324_n18# 0 0.360407f
C259 SUNSAR_CAPT8B_CV_0/XC08/XA0/MN1/a_324_n18# 0 0.422415f
C260 SUNSAR_CAPT8B_CV_0/XC08/XA0/MP1/a_216_n18# 0 0.091271f
C261 SUNSAR_CAPT8B_CV_0/XE10/XA7/C 0 2.352415f
C262 SUNSAR_CAPT8B_CV_0/XE10/QN 0 0.966414f
C263 uo_out[4] 0 1.095506f
C264 SUNSAR_CAPT8B_CV_0/XE10/XA8/MN0/a_324_334# 0 0.422f
C265 SUNSAR_CAPT8B_CV_0/XE10/XA8/MP0/a_216_334# 0 0.091271f
C266 SUNSAR_CAPT8B_CV_0/XE10/XA8/MN0/a_324_n18# 0 0.360407f
C267 SUNSAR_CAPT8B_CV_0/XE10/XA7/MN0/a_324_n18# 0 0.360407f
C268 SUNSAR_CAPT8B_CV_0/XE10/XA6/MN0/a_324_n18# 0 0.360407f
C269 SUNSAR_CAPT8B_CV_0/XE10/XA5/A 0 0.896691f
C270 SUNSAR_CAPT8B_CV_0/XE10/XA6/A 0 1.098676f
C271 SUNSAR_CAPT8B_CV_0/XE10/XA5/MN0/a_324_n18# 0 0.360407f
C272 SUNSAR_CAPT8B_CV_0/XE10/XA4/MN0/a_324_n18# 0 0.360407f
C273 SUNSAR_CAPT8B_CV_0/XE10/XA3/MN0/a_324_n18# 0 0.360407f
C274 SUNSAR_CAPT8B_CV_0/XE10/XA6/C 0 1.328497f
C275 SUNSAR_CAPT8B_CV_0/XE10/XA2/MN0/a_324_n18# 0 0.360407f
C276 SUNSAR_CAPT8B_CV_0/XE10/XA1/MN0/a_324_n18# 0 0.360407f
C277 SUNSAR_CAPT8B_CV_0/XE10/XA0/MN1/a_324_n18# 0 0.422415f
C278 SUNSAR_CAPT8B_CV_0/XE10/XA0/MP1/a_216_n18# 0 0.091271f
C279 SUNSAR_CAPT8B_CV_0/XG12/XA7/C 0 2.352415f
C280 SUNSAR_CAPT8B_CV_0/XG12/QN 0 0.966414f
C281 uo_out[2] 0 1.120428f
C282 SUNSAR_CAPT8B_CV_0/XG12/XA8/MN0/a_324_334# 0 0.422f
C283 SUNSAR_CAPT8B_CV_0/XG12/XA8/MP0/a_216_334# 0 0.091271f
C284 SUNSAR_CAPT8B_CV_0/XG12/XA8/MN0/a_324_n18# 0 0.360407f
C285 SUNSAR_CAPT8B_CV_0/XG12/XA7/MN0/a_324_n18# 0 0.360407f
C286 SUNSAR_CAPT8B_CV_0/XG12/XA6/MN0/a_324_n18# 0 0.360407f
C287 SUNSAR_CAPT8B_CV_0/XG12/XA5/A 0 0.896691f
C288 SUNSAR_CAPT8B_CV_0/XG12/XA6/A 0 1.098676f
C289 SUNSAR_CAPT8B_CV_0/XG12/XA5/MN0/a_324_n18# 0 0.360407f
C290 SUNSAR_CAPT8B_CV_0/XG12/XA4/MN0/a_324_n18# 0 0.360407f
C291 SUNSAR_CAPT8B_CV_0/XG12/XA3/MN0/a_324_n18# 0 0.360407f
C292 SUNSAR_CAPT8B_CV_0/XG12/XA6/C 0 1.328497f
C293 SUNSAR_CAPT8B_CV_0/XG12/XA2/MN0/a_324_n18# 0 0.360407f
C294 SUNSAR_CAPT8B_CV_0/XG12/XA1/MN0/a_324_n18# 0 0.360407f
C295 SUNSAR_CAPT8B_CV_0/XG12/XA0/MN1/a_324_n18# 0 0.422415f
C296 SUNSAR_CAPT8B_CV_0/XG12/XA0/MP1/a_216_n18# 0 0.091271f
C297 SUNSAR_CAPT8B_CV_0/XI14/XA7/C 0 2.352415f
C298 SUNSAR_CAPT8B_CV_0/XI14/QN 0 0.966414f
C299 uo_out[0] 0 1.493281f
C300 SUNSAR_CAPT8B_CV_0/XI14/XA8/MN0/a_324_334# 0 0.422f
C301 SUNSAR_CAPT8B_CV_0/XI14/XA8/MP0/a_216_334# 0 0.091271f
C302 SUNSAR_CAPT8B_CV_0/XI14/XA8/MN0/a_324_n18# 0 0.360407f
C303 SUNSAR_CAPT8B_CV_0/XI14/XA7/MN0/a_324_n18# 0 0.360407f
C304 SUNSAR_CAPT8B_CV_0/XI14/XA6/MN0/a_324_n18# 0 0.360407f
C305 SUNSAR_CAPT8B_CV_0/XI14/XA5/A 0 0.896691f
C306 SUNSAR_CAPT8B_CV_0/XI14/XA6/A 0 1.098676f
C307 SUNSAR_CAPT8B_CV_0/XI14/XA5/MN0/a_324_n18# 0 0.360407f
C308 SUNSAR_CAPT8B_CV_0/XI14/XA4/MN0/a_324_n18# 0 0.360407f
C309 SUNSAR_CAPT8B_CV_0/XI14/XA3/MN0/a_324_n18# 0 0.360407f
C310 SUNSAR_CAPT8B_CV_0/XI14/XA6/C 0 1.328497f
C311 SUNSAR_CAPT8B_CV_0/XI14/XA2/MN0/a_324_n18# 0 0.360407f
C312 SUNSAR_CAPT8B_CV_0/XI14/XA1/MN0/a_324_n18# 0 0.360407f
C313 SUNSAR_CAPT8B_CV_0/XI14/XA0/MN1/a_324_n18# 0 0.422415f
C314 SUNSAR_CAPT8B_CV_0/XI14/XA0/MP1/a_216_n18# 0 0.091271f
C315 ui_in[0] 0 3.522175f
C316 SUNSAR_CAPT8B_CV_0/XA1/MN1/a_324_334# 0 0.359492f
C317 SUNSAR_CAPT8B_CV_0/XB07/XA7/C 0 2.352415f
C318 SUNSAR_CAPT8B_CV_0/XB07/QN 0 0.966414f
C319 uo_out[7] 0 1.986758f
C320 SUNSAR_CAPT8B_CV_0/XB07/XA8/MN0/a_324_334# 0 0.422f
C321 SUNSAR_CAPT8B_CV_0/XB07/XA8/MP0/a_216_334# 0 0.091271f
C322 SUNSAR_CAPT8B_CV_0/XB07/XA8/MN0/a_324_n18# 0 0.360407f
C323 SUNSAR_CAPT8B_CV_0/XB07/XA7/MN0/a_324_n18# 0 0.360407f
C324 SUNSAR_CAPT8B_CV_0/XB07/XA6/MN0/a_324_n18# 0 0.360407f
C325 SUNSAR_CAPT8B_CV_0/XB07/XA5/A 0 0.896691f
C326 SUNSAR_CAPT8B_CV_0/XB07/XA6/A 0 1.098676f
C327 SUNSAR_CAPT8B_CV_0/XB07/XA5/MN0/a_324_n18# 0 0.360407f
C328 SUNSAR_CAPT8B_CV_0/XB07/XA4/MN0/a_324_n18# 0 0.360407f
C329 SUNSAR_CAPT8B_CV_0/XB07/XA3/MN0/a_324_n18# 0 0.360407f
C330 SUNSAR_CAPT8B_CV_0/XB07/XA6/C 0 1.328497f
C331 SUNSAR_CAPT8B_CV_0/XB07/XA2/MN0/a_324_n18# 0 0.360407f
C332 SUNSAR_SAR8B_CV_0/DONE 0 12.858106f
C333 SUNSAR_CAPT8B_CV_0/XB07/XA1/MN0/a_324_n18# 0 0.360407f
C334 SUNSAR_CAPT8B_CV_0/XB07/XA0/MN1/a_324_n18# 0 0.422415f
C335 SUNSAR_CAPT8B_CV_0/XB07/XA0/MP1/a_216_n18# 0 0.091271f
C336 SUNSAR_CAPT8B_CV_0/XD09/XA7/C 0 2.352415f
C337 SUNSAR_CAPT8B_CV_0/XD09/QN 0 0.966414f
C338 uo_out[5] 0 1.119996f
C339 SUNSAR_CAPT8B_CV_0/XD09/XA8/MN0/a_324_334# 0 0.422f
C340 SUNSAR_CAPT8B_CV_0/XD09/XA8/MP0/a_216_334# 0 0.091271f
C341 SUNSAR_CAPT8B_CV_0/XD09/XA8/MN0/a_324_n18# 0 0.360407f
C342 SUNSAR_CAPT8B_CV_0/XD09/XA7/MN0/a_324_n18# 0 0.360407f
C343 SUNSAR_CAPT8B_CV_0/XD09/XA6/MN0/a_324_n18# 0 0.360407f
C344 SUNSAR_CAPT8B_CV_0/XD09/XA5/A 0 0.896691f
C345 SUNSAR_CAPT8B_CV_0/XD09/XA6/A 0 1.098676f
C346 SUNSAR_CAPT8B_CV_0/XD09/XA5/MN0/a_324_n18# 0 0.360407f
C347 SUNSAR_CAPT8B_CV_0/XD09/XA4/MN0/a_324_n18# 0 0.360407f
C348 SUNSAR_CAPT8B_CV_0/XD09/XA3/MN0/a_324_n18# 0 0.360407f
C349 SUNSAR_CAPT8B_CV_0/XD09/XA6/C 0 1.328497f
C350 SUNSAR_CAPT8B_CV_0/XD09/XA2/MN0/a_324_n18# 0 0.360407f
C351 SUNSAR_CAPT8B_CV_0/XD09/XA1/MN0/a_324_n18# 0 0.360407f
C352 SUNSAR_CAPT8B_CV_0/XD09/XA0/MN1/a_324_n18# 0 0.422415f
C353 SUNSAR_CAPT8B_CV_0/XD09/XA0/MP1/a_216_n18# 0 0.091271f
C354 SUNSAR_SAR8B_CV_0/XA7/XA9/MN1/a_324_334# 0 0.360407f
C355 SUNSAR_SAR8B_CV_0/XA7/XA9/MN0/a_324_n18# 0 0.360407f
C356 SUNSAR_SAR8B_CV_0/XA7/XA9/A 0 1.250071f
C357 SUNSAR_SAR8B_CV_0/XA7/XA7/MN0/a_324_n18# 0 0.360407f
C358 SUNSAR_SAR8B_CV_0/XA7/XA8/MN0/a_324_n18# 0 0.360407f
C359 SUNSAR_SAR8B_CV_0/XA7/XA9/B 0 1.15806f
C360 SUNSAR_SAR8B_CV_0/XA7/XA6/MN0/a_324_n18# 0 0.360407f
C361 SUNSAR_SAR8B_CV_0/XA7/XA4/A 0 2.621765f
C362 SUNSAR_SAR8B_CV_0/XA7/XA4/MN0/a_324_n18# 0 0.360407f
C363 SUNSAR_SAR8B_CV_0/XA7/CP0 0 2.4163f
C364 SUNSAR_SAR8B_CV_0/XA7/CN0 0 0.312365f
C365 SUNSAR_SAR8B_CV_0/XA7/XA5/MN0/a_324_n18# 0 0.360407f
C366 SUNSAR_SAR8B_CV_0/XA7/CN1 0 2.428168f
C367 SUNSAR_SAR8B_CV_0/D<0> 0 1.87393f
C368 SUNSAR_SAR8B_CV_0/XA7/XA3/MN0/a_324_n18# 0 0.360407f
C369 SUNSAR_SAR8B_CV_0/XA7/XA2/A 0 2.030764f
C370 SUNSAR_SAR8B_CV_0/XA7/XA2/MN0/a_324_n18# 0 0.360407f
C371 SUNSAR_SAR8B_CV_0/XA7/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C372 SUNSAR_SAR8B_CV_0/XA7/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C373 SUNSAR_SAR8B_CV_0/XA7/XA1/XA2/Y 0 1.060197f
C374 SUNSAR_SAR8B_CV_0/XA7/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C375 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C376 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C377 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C378 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MP3/G 0 0.827484f
C379 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN2/S 0 0.200627f
C380 SUNSAR_SAR8B_CV_0/XA7/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C381 SUNSAR_SAR8B_CV_0/XA7/ENO 0 1.582724f
C382 SUNSAR_SAR8B_CV_0/XA7/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C383 SUNSAR_SAR8B_CV_0/XA7/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C384 SUNSAR_SAR8B_CV_0/XA7/XA13/MN1/a_324_334# 0 0.422f
C385 SUNSAR_SAR8B_CV_0/XA7/XA13/MP1/a_216_334# 0 0.091271f
C386 SUNSAR_SAR8B_CV_0/XA7/CEO 0 1.316615f
C387 SUNSAR_SAR8B_CV_0/XA7/XA12/MN0/a_324_n18# 0 0.360407f
C388 SUNSAR_SAR8B_CV_0/XA7/XA13/MN1/a_324_n18# 0 0.360407f
C389 SUNSAR_SAR8B_CV_0/XA7/XA12/A 0 0.755669f
C390 SUNSAR_SAR8B_CV_0/XA7/XA11/MN0/a_324_n18# 0 0.360407f
C391 SUNSAR_SAR8B_CV_0/XA6/CEO 0 1.009021f
C392 SUNSAR_SAR8B_CV_0/XA7/XA11/A 0 0.662715f
C393 SUNSAR_SAR8B_CV_0/XA7/XA9/Y 0 0.718246f
C394 SUNSAR_SAR8B_CV_0/XA6/XA9/MN1/a_324_334# 0 0.360407f
C395 SUNSAR_SAR8B_CV_0/XA6/XA9/MN0/a_324_n18# 0 0.360407f
C396 SUNSAR_SAR8B_CV_0/XA6/XA9/A 0 1.250071f
C397 SUNSAR_SAR8B_CV_0/XA6/DONE 0 0.13094f
C398 SUNSAR_SAR8B_CV_0/XA6/XA7/MN0/a_324_n18# 0 0.360407f
C399 SUNSAR_SAR8B_CV_0/XA6/XA8/MN0/a_324_n18# 0 0.360407f
C400 SUNSAR_SAR8B_CV_0/XA6/XA9/B 0 1.15806f
C401 SUNSAR_SAR8B_CV_0/XA6/XA6/MN0/a_324_n18# 0 0.360407f
C402 SUNSAR_SAR8B_CV_0/XA6/XA4/A 0 2.621765f
C403 SUNSAR_SAR8B_CV_0/XA6/XA4/MN0/a_324_n18# 0 0.360407f
C404 SUNSAR_SAR8B_CV_0/XA6/CP0 0 2.4163f
C405 SUNSAR_SAR8B_CV_0/XA6/CN0 0 4.160099f
C406 SUNSAR_SAR8B_CV_0/XA6/XA5/MN0/a_324_n18# 0 0.360407f
C407 SUNSAR_SAR8B_CV_0/XA6/CN1 0 2.428168f
C408 SUNSAR_SAR8B_CV_0/D<1> 0 5.818007f
C409 SUNSAR_SAR8B_CV_0/XA6/XA3/MN0/a_324_n18# 0 0.360407f
C410 SUNSAR_SAR8B_CV_0/XA6/XA2/A 0 2.030764f
C411 SUNSAR_SAR8B_CV_0/XA6/XA2/MN0/a_324_n18# 0 0.360407f
C412 SUNSAR_SAR8B_CV_0/XA6/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C413 SUNSAR_SAR8B_CV_0/XA6/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C414 SUNSAR_SAR8B_CV_0/XA6/XA1/XA2/Y 0 1.060197f
C415 SUNSAR_SAR8B_CV_0/XA6/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C416 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C417 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C418 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C419 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MP3/G 0 0.827484f
C420 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN2/S 0 0.200627f
C421 SUNSAR_SAR8B_CV_0/XA6/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C422 SUNSAR_SAR8B_CV_0/XA7/EN 0 3.856368f
C423 SUNSAR_SAR8B_CV_0/XA6/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C424 SUNSAR_SAR8B_CV_0/XA6/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C425 SUNSAR_SAR8B_CV_0/XA6/XA13/MN1/a_324_334# 0 0.422f
C426 SUNSAR_SAR8B_CV_0/XA6/XA13/MP1/a_216_334# 0 0.091271f
C427 SUNSAR_SAR8B_CV_0/XA6/XA12/MN0/a_324_n18# 0 0.360407f
C428 SUNSAR_SAR8B_CV_0/XA6/XA13/MN1/a_324_n18# 0 0.360407f
C429 SUNSAR_SAR8B_CV_0/XA6/XA12/A 0 0.755669f
C430 SUNSAR_SAR8B_CV_0/XA6/XA11/MN0/a_324_n18# 0 0.360407f
C431 SUNSAR_SAR8B_CV_0/XA5/CEO 0 1.104751f
C432 SUNSAR_SAR8B_CV_0/XA6/XA11/A 0 0.662715f
C433 SUNSAR_SAR8B_CV_0/XA6/XA9/Y 0 0.718246f
C434 SUNSAR_SAR8B_CV_0/XA5/XA9/MN1/a_324_334# 0 0.360407f
C435 SUNSAR_SAR8B_CV_0/XA5/XA9/MN0/a_324_n18# 0 0.360407f
C436 SUNSAR_SAR8B_CV_0/XA5/XA9/A 0 1.250071f
C437 SUNSAR_SAR8B_CV_0/XA5/DONE 0 0.123486f
C438 SUNSAR_SAR8B_CV_0/XA5/XA7/MN0/a_324_n18# 0 0.360407f
C439 SUNSAR_SAR8B_CV_0/XA5/XA8/MN0/a_324_n18# 0 0.360407f
C440 SUNSAR_SAR8B_CV_0/XA5/XA9/B 0 1.15806f
C441 SUNSAR_SAR8B_CV_0/XA5/XA6/MN0/a_324_n18# 0 0.360407f
C442 SUNSAR_SAR8B_CV_0/XA5/XA4/A 0 2.621765f
C443 SUNSAR_SAR8B_CV_0/XA5/XA4/MN0/a_324_n18# 0 0.360407f
C444 SUNSAR_SAR8B_CV_0/XA5/CP0 0 2.4163f
C445 SUNSAR_SAR8B_CV_0/XA5/CN0 0 3.052303f
C446 SUNSAR_SAR8B_CV_0/XA5/XA5/MN0/a_324_n18# 0 0.360407f
C447 SUNSAR_SAR8B_CV_0/XA5/CN1 0 2.428168f
C448 SUNSAR_SAR8B_CV_0/D<2> 0 5.190204f
C449 SUNSAR_SAR8B_CV_0/XA5/XA3/MN0/a_324_n18# 0 0.360407f
C450 SUNSAR_SAR8B_CV_0/XA5/XA2/A 0 2.030764f
C451 SUNSAR_SAR8B_CV_0/XA5/XA2/MN0/a_324_n18# 0 0.360407f
C452 SUNSAR_SAR8B_CV_0/XA5/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C453 SUNSAR_SAR8B_CV_0/XA5/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C454 SUNSAR_SAR8B_CV_0/XA5/XA1/XA2/Y 0 1.060197f
C455 SUNSAR_SAR8B_CV_0/XA5/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C456 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C457 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C458 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C459 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MP3/G 0 0.827484f
C460 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN2/S 0 0.200627f
C461 SUNSAR_SAR8B_CV_0/XA5/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C462 SUNSAR_SAR8B_CV_0/XA6/EN 0 3.679756f
C463 SUNSAR_SAR8B_CV_0/XA5/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C464 SUNSAR_SAR8B_CV_0/XA5/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C465 SUNSAR_SAR8B_CV_0/XA5/XA13/MN1/a_324_334# 0 0.422f
C466 SUNSAR_SAR8B_CV_0/XA5/XA13/MP1/a_216_334# 0 0.091271f
C467 SUNSAR_SAR8B_CV_0/XA5/XA12/MN0/a_324_n18# 0 0.360407f
C468 SUNSAR_SAR8B_CV_0/XA5/XA13/MN1/a_324_n18# 0 0.360407f
C469 SUNSAR_SAR8B_CV_0/XA5/XA12/A 0 0.755669f
C470 SUNSAR_SAR8B_CV_0/XA5/XA11/MN0/a_324_n18# 0 0.360407f
C471 SUNSAR_SAR8B_CV_0/XA4/CEO 0 1.086041f
C472 SUNSAR_SAR8B_CV_0/XA5/XA11/A 0 0.662715f
C473 SUNSAR_SAR8B_CV_0/XA5/XA9/Y 0 0.718246f
C474 SUNSAR_SAR8B_CV_0/XA4/XA9/MN1/a_324_334# 0 0.360407f
C475 SUNSAR_SAR8B_CV_0/XA4/XA9/MN0/a_324_n18# 0 0.360407f
C476 SUNSAR_SAR8B_CV_0/XA4/XA9/A 0 1.250071f
C477 SUNSAR_SAR8B_CV_0/XA4/DONE 0 0.13094f
C478 SUNSAR_SAR8B_CV_0/XA4/XA7/MN0/a_324_n18# 0 0.360407f
C479 SUNSAR_SAR8B_CV_0/XA4/XA8/MN0/a_324_n18# 0 0.360407f
C480 SUNSAR_SAR8B_CV_0/XA4/XA9/B 0 1.15806f
C481 SUNSAR_SAR8B_CV_0/XA4/XA6/MN0/a_324_n18# 0 0.360407f
C482 SUNSAR_SAR8B_CV_0/XA4/XA4/A 0 2.621765f
C483 SUNSAR_SAR8B_CV_0/XA4/XA4/MN0/a_324_n18# 0 0.360407f
C484 SUNSAR_SAR8B_CV_0/XA4/CP0 0 2.4163f
C485 SUNSAR_SAR8B_CV_0/XA4/CN0 0 2.237548f
C486 SUNSAR_SAR8B_CV_0/XA4/XA5/MN0/a_324_n18# 0 0.360407f
C487 SUNSAR_SAR8B_CV_0/XA4/CN1 0 2.428168f
C488 SUNSAR_SAR8B_CV_0/D<3> 0 4.013408f
C489 SUNSAR_SAR8B_CV_0/XA4/XA3/MN0/a_324_n18# 0 0.360407f
C490 SUNSAR_SAR8B_CV_0/XA4/XA2/A 0 2.030764f
C491 SUNSAR_SAR8B_CV_0/XA4/XA2/MN0/a_324_n18# 0 0.360407f
C492 SUNSAR_SAR8B_CV_0/XA4/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C493 SUNSAR_SAR8B_CV_0/XA4/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C494 SUNSAR_SAR8B_CV_0/XA4/XA1/XA2/Y 0 1.060197f
C495 SUNSAR_SAR8B_CV_0/XA4/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C496 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C497 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C498 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C499 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MP3/G 0 0.827484f
C500 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN2/S 0 0.200627f
C501 SUNSAR_SAR8B_CV_0/XA4/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C502 SUNSAR_SAR8B_CV_0/XA5/EN 0 3.635208f
C503 SUNSAR_SAR8B_CV_0/XA4/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C504 SUNSAR_SAR8B_CV_0/XA4/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C505 SUNSAR_SAR8B_CV_0/XA4/XA13/MN1/a_324_334# 0 0.422f
C506 SUNSAR_SAR8B_CV_0/XA4/XA13/MP1/a_216_334# 0 0.091271f
C507 SUNSAR_SAR8B_CV_0/XA4/XA12/MN0/a_324_n18# 0 0.360407f
C508 SUNSAR_SAR8B_CV_0/XA4/XA13/MN1/a_324_n18# 0 0.360407f
C509 SUNSAR_SAR8B_CV_0/XA4/XA12/A 0 0.755669f
C510 SUNSAR_SAR8B_CV_0/XA4/XA11/MN0/a_324_n18# 0 0.360407f
C511 SUNSAR_SAR8B_CV_0/XA3/CEO 0 1.107611f
C512 SUNSAR_SAR8B_CV_0/XA4/XA11/A 0 0.662715f
C513 SUNSAR_SAR8B_CV_0/XA4/XA9/Y 0 0.718246f
C514 SUNSAR_SAR8B_CV_0/XA3/XA9/MN1/a_324_334# 0 0.360407f
C515 SUNSAR_SAR8B_CV_0/XA3/XA9/MN0/a_324_n18# 0 0.360407f
C516 SUNSAR_SAR8B_CV_0/XA3/XA9/A 0 1.250071f
C517 SUNSAR_SAR8B_CV_0/XA3/DONE 0 0.123486f
C518 SUNSAR_SAR8B_CV_0/XA3/XA7/MN0/a_324_n18# 0 0.360407f
C519 SUNSAR_SAR8B_CV_0/XA3/XA8/MN0/a_324_n18# 0 0.360407f
C520 SUNSAR_SAR8B_CV_0/XA3/XA9/B 0 1.15806f
C521 SUNSAR_SAR8B_CV_0/XA3/XA6/MN0/a_324_n18# 0 0.360407f
C522 SUNSAR_SAR8B_CV_0/XA3/XA4/A 0 2.621765f
C523 SUNSAR_SAR8B_CV_0/XA3/XA4/MN0/a_324_n18# 0 0.360407f
C524 SUNSAR_SAR8B_CV_0/XA3/CP0 0 2.4163f
C525 SUNSAR_SAR8B_CV_0/XA3/CN0 0 3.224855f
C526 SUNSAR_SAR8B_CV_0/XA3/XA5/MN0/a_324_n18# 0 0.360407f
C527 SUNSAR_SAR8B_CV_0/XA3/CN1 0 2.428168f
C528 SUNSAR_SAR8B_CV_0/D<4> 0 4.549352f
C529 SUNSAR_SAR8B_CV_0/XA3/XA3/MN0/a_324_n18# 0 0.360407f
C530 SUNSAR_SAR8B_CV_0/XA3/XA2/A 0 2.030764f
C531 SUNSAR_SAR8B_CV_0/XA3/XA2/MN0/a_324_n18# 0 0.360407f
C532 SUNSAR_SAR8B_CV_0/XA3/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C533 SUNSAR_SAR8B_CV_0/XA3/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C534 SUNSAR_SAR8B_CV_0/XA3/XA1/XA2/Y 0 1.060197f
C535 SUNSAR_SAR8B_CV_0/XA3/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C536 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C537 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C538 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C539 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MP3/G 0 0.827484f
C540 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN2/S 0 0.200627f
C541 SUNSAR_SAR8B_CV_0/XA3/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C542 SUNSAR_SAR8B_CV_0/XA4/EN 0 3.720665f
C543 SUNSAR_SAR8B_CV_0/XA3/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C544 SUNSAR_SAR8B_CV_0/XA3/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C545 SUNSAR_SAR8B_CV_0/XA3/XA13/MN1/a_324_334# 0 0.422f
C546 SUNSAR_SAR8B_CV_0/XA3/XA13/MP1/a_216_334# 0 0.091271f
C547 SUNSAR_SAR8B_CV_0/XA3/XA12/MN0/a_324_n18# 0 0.360407f
C548 SUNSAR_SAR8B_CV_0/XA3/XA13/MN1/a_324_n18# 0 0.360407f
C549 SUNSAR_SAR8B_CV_0/XA3/XA12/A 0 0.755669f
C550 SUNSAR_SAR8B_CV_0/XA3/XA11/MN0/a_324_n18# 0 0.360407f
C551 SUNSAR_SAR8B_CV_0/XA2/CEO 0 1.085281f
C552 SUNSAR_SAR8B_CV_0/XA3/XA11/A 0 0.662715f
C553 SUNSAR_SAR8B_CV_0/XA3/XA9/Y 0 0.718246f
C554 SUNSAR_SAR8B_CV_0/XA2/XA9/MN1/a_324_334# 0 0.360407f
C555 SUNSAR_SAR8B_CV_0/XA2/XA9/MN0/a_324_n18# 0 0.360407f
C556 SUNSAR_SAR8B_CV_0/XA2/XA9/A 0 1.250071f
C557 SUNSAR_SAR8B_CV_0/XA2/DONE 0 0.13094f
C558 SUNSAR_SAR8B_CV_0/XA2/XA7/MN0/a_324_n18# 0 0.360407f
C559 SUNSAR_SAR8B_CV_0/XA2/XA8/MN0/a_324_n18# 0 0.360407f
C560 SUNSAR_SAR8B_CV_0/XA2/XA9/B 0 1.15806f
C561 SUNSAR_SAR8B_CV_0/XA2/XA6/MN0/a_324_n18# 0 0.360407f
C562 SUNSAR_SAR8B_CV_0/XA2/XA4/A 0 2.621765f
C563 SUNSAR_SAR8B_CV_0/XA2/XA4/MN0/a_324_n18# 0 0.360407f
C564 SUNSAR_SAR8B_CV_0/XA2/CP0 0 4.49437f
C565 SUNSAR_SAR8B_CV_0/XA2/CN0 0 2.820252f
C566 SUNSAR_SAR8B_CV_0/XA2/XA5/MN0/a_324_n18# 0 0.360407f
C567 SUNSAR_SAR8B_CV_0/XA2/CN1 0 6.112935f
C568 SUNSAR_SAR8B_CV_0/XA2/XA3/MN0/a_324_n18# 0 0.360407f
C569 SUNSAR_SAR8B_CV_0/XA2/XA2/A 0 2.030764f
C570 SUNSAR_SAR8B_CV_0/XA2/XA2/MN0/a_324_n18# 0 0.360407f
C571 SUNSAR_SAR8B_CV_0/XA2/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C572 SUNSAR_SAR8B_CV_0/XA2/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C573 SUNSAR_SAR8B_CV_0/XA2/XA1/XA2/Y 0 1.060197f
C574 SUNSAR_SAR8B_CV_0/XA2/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C575 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C576 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C577 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C578 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MP3/G 0 0.827484f
C579 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN2/S 0 0.200627f
C580 SUNSAR_SAR8B_CV_0/XA2/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C581 SUNSAR_SAR8B_CV_0/XA3/EN 0 3.784028f
C582 SUNSAR_SAR8B_CV_0/XA2/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C583 SUNSAR_SAR8B_CV_0/XA2/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C584 SUNSAR_SAR8B_CV_0/XA2/XA13/MN1/a_324_334# 0 0.422f
C585 SUNSAR_SAR8B_CV_0/XA2/XA13/MP1/a_216_334# 0 0.091271f
C586 SUNSAR_SAR8B_CV_0/XA2/XA12/MN0/a_324_n18# 0 0.360407f
C587 SUNSAR_SAR8B_CV_0/XA2/XA13/MN1/a_324_n18# 0 0.360407f
C588 SUNSAR_SAR8B_CV_0/XA2/XA12/A 0 0.755669f
C589 SUNSAR_SAR8B_CV_0/XA2/XA11/MN0/a_324_n18# 0 0.360407f
C590 SUNSAR_SAR8B_CV_0/XA1/CEO 0 1.104751f
C591 SUNSAR_SAR8B_CV_0/XA2/XA11/A 0 0.662715f
C592 SUNSAR_SAR8B_CV_0/XA2/XA9/Y 0 0.718246f
C593 SUNSAR_SAR8B_CV_0/XA1/XA9/MN1/a_324_334# 0 0.360407f
C594 SUNSAR_SAR8B_CV_0/XA1/XA9/MN0/a_324_n18# 0 0.360407f
C595 SUNSAR_SAR8B_CV_0/XA1/XA9/A 0 1.250071f
C596 SUNSAR_SAR8B_CV_0/XA1/DONE 0 0.123486f
C597 SUNSAR_SAR8B_CV_0/XA1/XA7/MN0/a_324_n18# 0 0.360407f
C598 SUNSAR_SAR8B_CV_0/XA1/XA8/MN0/a_324_n18# 0 0.360407f
C599 SUNSAR_SAR8B_CV_0/XA1/XA9/B 0 1.15806f
C600 SUNSAR_SAR8B_CV_0/XA1/XA6/MN0/a_324_n18# 0 0.360407f
C601 SUNSAR_SAR8B_CV_0/XA1/XA4/A 0 2.621765f
C602 SUNSAR_SAR8B_CV_0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C603 SUNSAR_SAR8B_CV_0/XA1/CP0 0 4.486094f
C604 SUNSAR_SAR8B_CV_0/XA1/CN0 0 2.798774f
C605 SUNSAR_SAR8B_CV_0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C606 SUNSAR_SAR8B_CV_0/XA1/CN1 0 4.70217f
C607 SUNSAR_SAR8B_CV_0/D<6> 0 4.492109f
C608 SUNSAR_SAR8B_CV_0/XA1/XA3/MN0/a_324_n18# 0 0.360407f
C609 SUNSAR_SAR8B_CV_0/XA1/XA2/A 0 2.030764f
C610 SUNSAR_SAR8B_CV_0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C611 SUNSAR_SAR8B_CV_0/XA1/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C612 SUNSAR_SAR8B_CV_0/XA1/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C613 SUNSAR_SAR8B_CV_0/XA1/XA1/XA2/Y 0 1.060197f
C614 SUNSAR_SAR8B_CV_0/XA1/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C615 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C616 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C617 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C618 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MP3/G 0 0.827484f
C619 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN2/S 0 0.200627f
C620 SUNSAR_SAR8B_CV_0/XA1/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C621 SUNSAR_SAR8B_CV_0/XA2/EN 0 3.720665f
C622 SUNSAR_SAR8B_CV_0/XA1/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C623 SUNSAR_SAR8B_CV_0/XA1/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C624 SUNSAR_SAR8B_CV_0/XA1/XA13/MN1/a_324_334# 0 0.422f
C625 SUNSAR_SAR8B_CV_0/XA1/XA13/MP1/a_216_334# 0 0.091271f
C626 SUNSAR_SAR8B_CV_0/XA1/XA12/MN0/a_324_n18# 0 0.360407f
C627 SUNSAR_SAR8B_CV_0/XA1/XA13/MN1/a_324_n18# 0 0.360407f
C628 SUNSAR_SAR8B_CV_0/XA1/XA12/A 0 0.755669f
C629 SUNSAR_SAR8B_CV_0/XA1/XA11/MN0/a_324_n18# 0 0.360407f
C630 SUNSAR_SAR8B_CV_0/XA0/CEO 0 1.083361f
C631 SUNSAR_SAR8B_CV_0/XA1/XA11/A 0 0.662715f
C632 SUNSAR_SAR8B_CV_0/XA1/XA9/Y 0 0.718246f
C633 SUNSAR_SAR8B_CV_0/XB2/XA7/MN1/a_324_n18# 0 0.359583f
C634 SUNSAR_SAR8B_CV_0/XB2/XA5b/MN1/a_324_n18# 0 0.422415f
C635 SUNSAR_SAR8B_CV_0/XB2/XA5b/MP1/a_216_n18# 0 0.091271f
C636 SUNSAR_SAR8B_CV_0/XB2/XA1/Y 0 0.690197f
C637 SUNSAR_SAR8B_CV_0/XB2/CKN 0 1.768971f
C638 SUNSAR_SAR8B_CV_0/XB2/XA4/MN0/a_324_n18# 0 0.359583f
C639 SUNSAR_SAR8B_CV_0/XB2/XA5/MN1/a_324_334# 0 0.422f
C640 SUNSAR_SAR8B_CV_0/XB2/XA5/MP1/a_216_334# 0 0.091271f
C641 SUNSAR_SAR8B_CV_0/XB2/XA3/MP0/S 0 0.743486f
C642 SUNSAR_SAR8B_CV_0/XB2/XA3/MN0/a_324_n18# 0 0.359583f
C643 SUNSAR_SAR8B_CV_0/XB2/XA2/MP0/G 0 0.708335f
C644 SUNSAR_SAR8B_CV_0/XB2/XA7/MN1/a_324_334# 0 0.359583f
C645 SUNSAR_SAR8B_CV_0/XB2/XA5/MN1/a_324_n18# 0 0.360407f
C646 SUNSAR_SAR8B_CV_0/XB2/XA1/MP0/G 0 0.788614f
C647 SUNSAR_SAR8B_CV_0/XB2/XA4/MN1/a_324_334# 0 0.359583f
C648 SUNSAR_SAR8B_CV_0/XB2/XA0/MN0/a_324_n18# 0 0.359583f
C649 SUNSAR_SAR8B_CV_0/XB2/M8/a_324_n18# 0 0.356977f
C650 SUNSAR_SAR8B_CV_0/XB2/M8/a_324_334# 0 0.422f
C651 SUNSAR_SAR8B_CV_0/XB2/M6/a_324_n18# 0 0.356977f
C652 SUNSAR_SAR8B_CV_0/XB2/M7/a_324_n18# 0 0.356977f
C653 SUNSAR_SAR8B_CV_0/XB2/XA3/B 0 54.41209f
C654 SUNSAR_SAR8B_CV_0/XB2/XA4/GNG 0 53.065117f
C655 SUNSAR_SAR8B_CV_0/XB2/M5/a_324_n18# 0 0.356977f
C656 SUNSAR_SAR8B_CV_0/XB2/M3/a_324_n18# 0 0.356977f
C657 SUNSAR_SAR8B_CV_0/XB2/M4/a_324_n18# 0 0.356977f
C658 SUNSAR_SAR8B_CV_0/XB2/M4/G 0 2.475647f
C659 ua[0] 0 2.335287f
C660 SUNSAR_SAR8B_CV_0/XB2/M1/a_324_n18# 0 0.422415f
C661 SUNSAR_SAR8B_CV_0/XB2/M2/a_324_n18# 0 0.356977f
C662 SUNSAR_SAR8B_CV_0/XA0/XA9/MN1/a_324_334# 0 0.360407f
C663 SUNSAR_SAR8B_CV_0/XA0/XA9/MN0/a_324_n18# 0 0.360407f
C664 SUNSAR_SAR8B_CV_0/XA0/XA9/A 0 1.250071f
C665 SUNSAR_SAR8B_CV_0/XA0/DONE 0 0.134046f
C666 SUNSAR_SAR8B_CV_0/XA0/XA7/MN0/a_324_n18# 0 0.360407f
C667 SUNSAR_SAR8B_CV_0/XA0/XA8/MN0/a_324_n18# 0 0.360407f
C668 SUNSAR_SAR8B_CV_0/XA0/XA9/B 0 1.15806f
C669 SUNSAR_SAR8B_CV_0/CK_SAMPLE 0 17.082773f
C670 SUNSAR_SAR8B_CV_0/XA0/XA6/MN0/a_324_n18# 0 0.360407f
C671 SUNSAR_SAR8B_CV_0/XA0/XA4/A 0 2.621765f
C672 SUNSAR_SAR8B_CV_0/XA0/XA4/MN0/a_324_n18# 0 0.360407f
C673 SUNSAR_SAR8B_CV_0/XA0/CP0 0 8.48089f
C674 SUNSAR_SAR8B_CV_0/XA0/XA5/MN0/a_324_n18# 0 0.360407f
C675 SUNSAR_SAR8B_CV_0/D<7> 0 9.577809f
C676 SUNSAR_SAR8B_CV_0/XA0/XA3/MN0/a_324_n18# 0 0.360407f
C677 SUNSAR_SAR8B_CV_0/XA0/XA2/A 0 2.030764f
C678 SUNSAR_SAR8B_CV_0/XA0/XA2/MN0/a_324_n18# 0 0.360407f
C679 SUNSAR_SAR8B_CV_0/XA0/XA1/XA5/MN0/a_324_n18# 0 0.360407f
C680 SUNSAR_SAR8B_CV_0/EN 0 5.97155f
C681 SUNSAR_SAR8B_CV_0/XA0/XA1/XA4/MN0/a_324_n18# 0 0.360407f
C682 SUNSAR_SAR8B_CV_0/XA0/XA1/XA2/Y 0 1.060197f
C683 SUNSAR_SAR8B_CV_0/XA0/XA1/XA2/MN0/a_324_n18# 0 0.360407f
C684 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN3/a_324_n18# 0 0.355196f
C685 SUNSAR_SAR8B_CV_0/XA20/CPO 0 11.091676f
C686 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN2/a_324_n18# 0 0.355196f
C687 SUNSAR_SAR8B_CV_0/XA20/CNO 0 12.667546f
C688 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN1/a_324_n18# 0 0.355196f
C689 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MP3/G 0 0.827484f
C690 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN2/S 0 0.200627f
C691 SUNSAR_SAR8B_CV_0/XA0/XA1/XA1/MN0/a_324_n18# 0 0.360407f
C692 SUNSAR_SAR8B_CV_0/XA1/EN 0 3.794638f
C693 SUNSAR_SAR8B_CV_0/XA0/XA1/XA0/MN1/a_324_n18# 0 0.422415f
C694 VPWR 0 0.724279p
C695 SUNSAR_SAR8B_CV_0/XA0/XA1/XA0/MP1/a_216_n18# 0 0.091271f
C696 SUNSAR_SAR8B_CV_0/XA0/XA13/MN1/a_324_334# 0 0.422f
C697 SUNSAR_SAR8B_CV_0/XA0/XA13/MP1/a_216_334# 0 0.091271f
C698 SUNSAR_SAR8B_CV_0/XA0/XA12/MN0/a_324_n18# 0 0.360407f
C699 SUNSAR_SAR8B_CV_0/XA0/XA13/MN1/a_324_n18# 0 0.360407f
C700 SUNSAR_SAR8B_CV_0/XA0/XA12/A 0 0.755669f
C701 SUNSAR_SAR8B_CV_0/XA0/XA11/MN0/a_324_n18# 0 0.360407f
C702 SUNSAR_SAR8B_CV_0/XA0/XA11/A 0 0.662715f
C703 SUNSAR_SAR8B_CV_0/XA0/XA9/Y 0 0.718246f
C704 SUNSAR_SAR8B_CV_0/XB1/XA7/MN1/a_324_n18# 0 0.359583f
C705 VGND 0 0.221901p
C706 SUNSAR_SAR8B_CV_0/XB1/XA5b/MN1/a_324_n18# 0 0.422415f
C707 SUNSAR_SAR8B_CV_0/XB1/XA5b/MP1/a_216_n18# 0 0.091271f
C708 SUNSAR_SAR8B_CV_0/XB1/XA1/Y 0 0.690197f
C709 SUNSAR_SAR8B_CV_0/XB1/CKN 0 1.768971f
C710 SUNSAR_SAR8B_CV_0/XB1/XA4/MN0/a_324_n18# 0 0.359583f
C711 SUNSAR_SAR8B_CV_0/XB1/XA5/MN1/a_324_334# 0 0.422f
C712 SUNSAR_SAR8B_CV_0/XB1/XA5/MP1/a_216_334# 0 0.091271f
C713 SUNSAR_SAR8B_CV_0/XB1/XA3/MP0/S 0 0.743486f
C714 SUNSAR_SAR8B_CV_0/XB1/XA3/MN0/a_324_n18# 0 0.359583f
C715 SUNSAR_SAR8B_CV_0/XB1/XA2/MP0/G 0 0.708335f
C716 SUNSAR_SAR8B_CV_0/XB1/XA7/MN1/a_324_334# 0 0.359583f
C717 SUNSAR_SAR8B_CV_0/XB1/XA5/MN1/a_324_n18# 0 0.360407f
C718 SUNSAR_SAR8B_CV_0/XB1/XA1/MP0/G 0 0.788614f
C719 SUNSAR_SAR8B_CV_0/XB1/XA4/MN1/a_324_334# 0 0.359583f
C720 SUNSAR_SAR8B_CV_0/CK_SAMPLE_BSSW 0 6.759625f
C721 SUNSAR_SAR8B_CV_0/XB1/XA0/MN0/a_324_n18# 0 0.359583f
C722 SUNSAR_SAR8B_CV_0/XB1/M8/a_324_n18# 0 0.356977f
C723 SUNSAR_SAR8B_CV_0/XB1/M8/a_324_334# 0 0.422f
C724 SUNSAR_SAR8B_CV_0/XB1/M6/a_324_n18# 0 0.356977f
C725 SUNSAR_SAR8B_CV_0/XB1/M7/a_324_n18# 0 0.356977f
C726 SUNSAR_SAR8B_CV_0/XB1/XA3/B 0 54.41209f
C727 SUNSAR_SAR8B_CV_0/XB1/XA4/GNG 0 53.065117f
C728 SUNSAR_SAR8B_CV_0/XA0/CEIN 0 19.901903f
C729 SUNSAR_SAR8B_CV_0/XB1/M5/a_324_n18# 0 0.356977f
C730 SUNSAR_SAR8B_CV_0/XB1/M3/a_324_n18# 0 0.356977f
C731 SUNSAR_SAR8B_CV_0/XB1/M4/a_324_n18# 0 0.356977f
C732 SUNSAR_SAR8B_CV_0/XB1/M4/G 0 2.475647f
C733 ua[1] 0 3.007717f
C734 SUNSAR_SAR8B_CV_0/XB1/M1/a_324_n18# 0 0.422415f
C735 SUNSAR_SAR8B_CV_0/XB1/M2/a_324_n18# 0 0.356977f
C736 SUNSAR_SAR8B_CV_0/XA20/XA9/MN0/a_324_n18# 0 0.360407f
C737 SUNSAR_SAR8B_CV_0/XA20/XA3/CO 0 2.703497f
C738 SUNSAR_SAR8B_CV_0/XA20/XA2/MN6/a_324_334# 0 0.360407f
C739 SUNSAR_SAR8B_CV_0/XA20/XA3a/A 0 2.536943f
C740 SUNSAR_SAR8B_CV_0/XA20/XA3/MN0/a_324_n18# 0 0.360407f
C741 SUNSAR_SAR8B_CV_0/XA20/XA3a/MN0/a_324_n18# 0 0.360407f
C742 SUNSAR_SAR8B_CV_0/XA20/XA4/MN0/a_324_n18# 0 0.360407f
C743 SUNSAR_SAR8B_CV_0/XA20/XA4/MP0/S 0 0.397005f
C744 SUNSAR_SAR8B_CV_0/SARN 0 30.043571f
C745 SUNSAR_SAR8B_CV_0/XA20/XA3/N2 0 0.234927f
C746 SUNSAR_SAR8B_CV_0/XA20/XA9/Y 0 3.176436f
C747 SUNSAR_SAR8B_CV_0/XA20/XA2/N2 0 0.234927f
C748 SUNSAR_SAR8B_CV_0/XA20/XA2/MN0/a_324_n18# 0 0.360407f
C749 SUNSAR_SAR8B_CV_0/XA20/XA3/N1 0 0.905385f
C750 SUNSAR_SAR8B_CV_0/SARP 0 30.653925f
C751 SUNSAR_SAR8B_CV_0/XA20/XA1/MN0/a_324_n18# 0 0.360407f
C752 SUNSAR_SAR8B_CV_0/XA20/XA1/MP0/S 0 0.397005f
C753 SUNSAR_SAR8B_CV_0/XA20/XA9/A 0 3.508213f
C754 SUNSAR_SAR8B_CV_0/XA20/XA0/MN1/a_324_n18# 0 0.422415f
C755 SUNSAR_SAR8B_CV_0/XA20/XA0/MP1/a_216_n18# 0 0.091271f
C756 SUNSAR_SAR8B_CV_0/XA20/XA13/MN1/a_324_n18# 0 0.360407f
C757 SUNSAR_SAR8B_CV_0/XA20/XA13/MN1/a_324_334# 0 0.422f
C758 SUNSAR_SAR8B_CV_0/XA20/XA13/MP1/a_216_334# 0 0.091271f
C759 SUNSAR_SAR8B_CV_0/XA20/XA12/MN0/a_324_n18# 0 0.360407f
C760 SUNSAR_SAR8B_CV_0/XA20/XA11/MN0/a_324_n18# 0 0.360407f
C761 SUNSAR_SAR8B_CV_0/XA20/XA9/MN0/a_324_334# 0 0.360407f
C762 SUNSAR_SAR8B_CV_0/XA20/XA12/Y 0 0.623344f
C763 SUNSAR_SAR8B_CV_0/XA20/XA11/Y 0 0.759612f
C764 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES2/B 0 3.1129f
C765 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES4/B 0 3.516117f
C766 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES8/B 0 3.933522f
C767 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES16/B 0 4.664508f
C768 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES1B/B 0 2.892833f
C769 SUNSAR_SAR8B_CV_0/XDAC2/XC32a<0>/XRES1A/B 0 1.735354f
C770 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES2/B 0 3.1129f
C771 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES4/B 0 3.516117f
C772 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES8/B 0 3.933522f
C773 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES16/B 0 4.664508f
C774 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES1B/B 0 2.892833f
C775 SUNSAR_SAR8B_CV_0/XDAC2/XC1/XRES1A/B 0 1.735354f
C776 SUNSAR_SAR8B_CV_0/XA0/CN0 0 6.776559f
C777 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES2/B 0 3.1129f
C778 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES4/B 0 3.516117f
C779 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES8/B 0 3.933522f
C780 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES16/B 0 4.664508f
C781 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES1B/B 0 2.892833f
C782 SUNSAR_SAR8B_CV_0/XDAC2/XC0/XRES1A/B 0 1.735354f
C783 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES2/B 0 3.1129f
C784 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES4/B 0 3.516117f
C785 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES8/B 0 3.933522f
C786 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES16/B 0 4.664508f
C787 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES1B/B 0 2.892833f
C788 SUNSAR_SAR8B_CV_0/XDAC2/X16ab/XRES1A/B 0 1.735354f
C789 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES2/B 0 3.1129f
C790 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES4/B 0 3.516117f
C791 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES8/B 0 3.933522f
C792 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES16/B 0 4.664508f
C793 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES1B/B 0 2.892833f
C794 SUNSAR_SAR8B_CV_0/XDAC1/XC32a<0>/XRES1A/B 0 1.735354f
C795 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES2/B 0 3.1129f
C796 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES4/B 0 3.516117f
C797 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES8/B 0 3.933522f
C798 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES16/B 0 4.664508f
C799 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES1B/B 0 2.892833f
C800 SUNSAR_SAR8B_CV_0/XDAC1/XC1/XRES1A/B 0 1.735354f
C801 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES2/B 0 3.1129f
C802 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES4/B 0 3.516117f
C803 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES8/B 0 3.933522f
C804 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES16/B 0 4.664508f
C805 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES1B/B 0 2.892833f
C806 SUNSAR_SAR8B_CV_0/XDAC1/XC0/XRES1A/B 0 1.735354f
C807 SUNSAR_SAR8B_CV_0/D<5> 0 5.830972f
C808 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES2/B 0 3.1129f
C809 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES4/B 0 3.516117f
C810 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES8/B 0 3.933522f
C811 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES16/B 0 4.664508f
C812 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES1B/B 0 2.892833f
C813 SUNSAR_SAR8B_CV_0/XDAC1/X16ab/XRES1A/B 0 1.735354f
C814 SUNSAR_SAR8B_CV_0/XA0/CP1 0 4.930175f
C815 tt_um_TT06_SAR_done_0/x5/MN1/a_324_334# 0 0.422f
C816 tt_um_TT06_SAR_done_0/x5/MP1/a_216_334# 0 0.091271f
C817 tt_um_TT06_SAR_done_0/x4/MP0/G 0 0.782647f
C818 tt_um_TT06_SAR_done_0/x5/MN1/a_324_n18# 0 0.360407f
C819 uio_oe[0] 0 1.551274f
C820 uio_out[0] 0 1.059239f
C821 tt_um_TT06_SAR_done_0/x3/MN1/a_324_n18# 0 0.355196f
C822 tt_um_TT06_SAR_done_0/x4/MN0/a_324_n18# 0 0.360407f
C823 tt_um_TT06_SAR_done_0/x3/MP1/G 0 0.95314f
C824 tt_um_TT06_SAR_done_0/x3/MN0/a_324_n18# 0 0.422415f
C825 tt_um_TT06_SAR_done_0/x3/MP0/a_216_n18# 0 0.091271f
.ends

