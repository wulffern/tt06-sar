* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1]
*+ uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1]
*+ uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7]
*+ ui_in[0] uo_out[6] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA4.A SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=240.8616 ps=1.269k w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=244.62 ps=1.28028k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X51 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X52 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X56 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X58 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X63 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X65 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X66 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X72 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X74 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X76 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X77 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X78 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X79 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 VPWR SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X88 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X90 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X95 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X96 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X97 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X98 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R8 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X99 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X100 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X101 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_CAPT8B_CV_0.XE10.XA4.A SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X106 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X107 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X108 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X114 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X115 SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X116 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 VGND SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X118 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R10 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X119 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X120 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X121 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X122 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X124 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X125 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X130 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X131 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X132 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X134 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X135 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X136 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X137 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X146 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X147 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X148 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X149 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X150 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X155 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R13 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X158 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X160 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X163 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X166 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R14 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X167 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X169 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X174 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X175 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R15 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X176 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X177 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X178 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X181 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X182 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X185 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X186 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X188 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X193 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X194 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X195 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X198 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R16 uio_oe[0] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
R17 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X199 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X201 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R18 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X205 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X206 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X207 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 VGND SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R19 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X212 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X213 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X214 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X216 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X221 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X223 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA3.XA11.Y SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X225 SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X228 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X229 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X230 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X232 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X233 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X235 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X236 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X237 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X239 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X246 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X247 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X250 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X252 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X253 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X255 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X256 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X258 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X259 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X261 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X263 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X264 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X266 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X268 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X270 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X274 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X275 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X276 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X277 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X278 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X279 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X280 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X281 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X282 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R23 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R24 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X283 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X284 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X286 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X292 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X294 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X299 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X300 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X301 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X304 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X306 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X307 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X308 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X309 VPWR SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X310 VGND SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X311 SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X312 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X313 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X314 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X315 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X316 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R25 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R26 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X317 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X318 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X319 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X320 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X321 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X322 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X323 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X324 SUNSAR_SAR8B_CV_0.XB2.XA3.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X327 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X328 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R27 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X329 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X330 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X331 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X332 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X333 SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X334 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X336 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X337 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X338 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X340 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X341 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X342 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X344 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X345 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X346 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R29 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X347 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X348 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X349 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X350 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X351 SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X352 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X354 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X355 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X359 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R30 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X360 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X361 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X364 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X365 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R31 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X366 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X367 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X368 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R32 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X369 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X370 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X371 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X372 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X373 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X374 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X375 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X376 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X377 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X378 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X379 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X381 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R34 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X382 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X384 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X385 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X386 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X387 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X389 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R35 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X390 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X391 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X393 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X394 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X395 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X396 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X397 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X400 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X402 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X404 SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X406 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X407 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R36 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R37 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X409 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X410 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X411 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X413 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X414 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X416 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X417 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X418 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X419 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X420 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X421 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X422 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X423 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X424 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R38 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X425 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X426 SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X427 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X428 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X429 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X431 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X433 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X434 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X435 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X436 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X437 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X438 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X440 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X441 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X442 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X443 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X444 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA7.CEO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R41 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X446 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X447 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X449 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X450 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X452 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X453 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X454 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X455 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X456 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X457 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X458 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X459 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R42 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X460 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R43 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X461 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X462 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X463 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X465 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X468 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X470 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X471 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X472 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R44 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X473 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X474 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X475 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X476 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X477 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X478 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X479 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X480 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X481 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X482 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 VGND SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X486 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X487 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X488 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X489 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X491 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X492 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X493 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X494 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X495 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X496 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X497 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X498 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X499 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X500 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R46 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X501 SUNSAR_CAPT8B_CV_0.XD09.XA4.A SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X502 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X503 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X505 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X506 SUNSAR_SAR8B_CV_0.XA5.XA11.Y SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X508 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X509 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X510 SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X511 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R48 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X512 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X513 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X514 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X515 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X516 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X517 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X519 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X520 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X521 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X522 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X523 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X525 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X526 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X527 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X528 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R49 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X529 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X530 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X531 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X532 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X533 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X536 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X537 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X540 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X541 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA20.XA10.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X544 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X545 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X548 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R51 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X549 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X550 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X552 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X553 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X554 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X556 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X557 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X558 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X559 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X560 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X561 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X562 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X564 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X565 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X567 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X568 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X569 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X570 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X571 SUNSAR_CAPT8B_CV_0.XA2.MN0.G SUNSAR_CAPT8B_CV_0.XA2.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X572 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X573 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X574 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X575 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X576 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X577 ua[1] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X578 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X579 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X580 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X581 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X582 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X583 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X584 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X585 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X587 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X588 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X589 SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X590 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R53 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X591 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X592 SUNSAR_SAR8B_CV_0.XA2.XA11.Y SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X593 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X594 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X595 VGND SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X596 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R54 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X598 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X599 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X600 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X601 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X602 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X603 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X604 VGND SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X605 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X606 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X609 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X610 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X611 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X613 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X614 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X616 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X618 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X619 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X621 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X624 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X626 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X630 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X631 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X637 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R55 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X640 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X642 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X644 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X645 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X647 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X648 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X649 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X650 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X652 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X653 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X654 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X655 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X656 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X657 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X658 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X659 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X660 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X661 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R57 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R58 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X662 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X663 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X664 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X665 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X666 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X667 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X669 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X670 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X674 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X675 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X676 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 SUNSAR_CAPT8B_CV_0.XC08.XA4.A SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X680 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X681 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X682 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X683 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X684 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X685 SUNSAR_SAR8B_CV_0.XA4.XA11.Y SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X686 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X687 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X688 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X690 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R60 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X691 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X692 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X693 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X694 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X695 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X696 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X697 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X699 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X700 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X701 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X704 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X705 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X706 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X707 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X709 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X710 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R61 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X711 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X712 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X713 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X714 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X715 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X716 SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X717 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X718 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X719 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R62 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X720 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X721 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X722 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X724 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X725 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X726 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X727 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X728 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X729 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X730 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X731 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X732 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 SUNSAR_CAPT8B_CV_0.XI14.XA4.A SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X734 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X735 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X736 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X737 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X738 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X739 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X740 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X741 ua[0] SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X742 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X744 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X745 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R65 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X746 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X747 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X748 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X749 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X750 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X751 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X752 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X753 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X754 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X755 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X756 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X759 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X760 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X762 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X763 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R67 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X764 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X765 VGND SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X766 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X767 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X768 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X769 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X770 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X771 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X772 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X773 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X774 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R68 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X777 VGND SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X778 SUNSAR_SAR8B_CV_0.XA1.XA11.Y SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X779 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X780 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X782 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X783 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X786 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X787 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X788 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X789 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X790 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X791 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X792 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X793 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X795 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X798 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA6.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X800 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X801 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X802 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X807 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X808 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X809 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X810 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X813 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X814 VGND SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X815 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X816 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X817 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X818 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X819 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X821 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X822 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X823 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X824 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X825 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X827 ua[1] SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X828 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X829 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X830 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X831 VGND SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X832 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X833 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X834 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X835 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R70 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X836 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X837 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X838 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X839 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R71 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X841 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X842 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X843 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X844 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X845 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X847 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X848 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X849 SUNSAR_SAR8B_CV_0.XA7.XA11.Y SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X850 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X852 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X853 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X854 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X855 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X858 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X859 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X862 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 SUNSAR_CAPT8B_CV_0.XB07.XA4.A SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X864 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 VGND SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X867 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X868 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_CAPT8B_CV_0.XH13.XA4.A SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X872 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X873 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X874 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X875 VGND SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X876 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X878 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X879 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 VGND SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X882 VPWR SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X883 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X884 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X885 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X886 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R72 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X887 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X890 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X892 VGND SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X893 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X894 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X895 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R73 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X896 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X897 VGND SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X899 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R74 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X900 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA6.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X901 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X902 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X903 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R75 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X905 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X906 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X907 VGND SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X909 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X910 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R76 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X911 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X912 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X913 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X914 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X915 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X916 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X917 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X918 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X920 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R77 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XA4.GNG sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X923 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X924 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X925 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.D SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X926 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X928 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X929 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X930 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X931 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X932 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X933 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X934 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X935 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R78 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X936 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X937 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X939 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R79 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X940 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X941 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X942 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X944 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X945 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X946 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X947 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X948 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA3.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X949 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X950 SUNSAR_SAR8B_CV_0.XB1.XA3.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X951 SUNSAR_CAPT8B_CV_0.XF11.XA4.A SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X953 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X954 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R80 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X955 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X956 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X957 VGND SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X959 VGND SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X961 TIE_L SUNSAR_CAPT8B_CV_0.XA2.MN0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X962 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X963 SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X964 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X965 SUNSAR_SAR8B_CV_0.XA6.XA11.Y SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R81 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XA3.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X967 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X969 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X970 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X971 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X972 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X974 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X975 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X976 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X978 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X979 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X980 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X982 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X984 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X985 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R82 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X986 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X987 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X988 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X992 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X993 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X994 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X995 ua[0] SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X996 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X997 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X999 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R83 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1000 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1001 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1002 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN0.D SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1004 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1005 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1006 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1007 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R84 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1008 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1012 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1013 VGND SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1014 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.D SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1016 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1017 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1018 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA0.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1019 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1020 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1021 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1022 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA6.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R85 uio_out[0] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X1025 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1031 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1033 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1034 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1035 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1036 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1037 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1038 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1039 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1040 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1041 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1042 VGND SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1043 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1044 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.D SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1045 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1046 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.649845f
C1 a_9990_4566# VPWR 0.413433f
C2 TIE_L TIE_L1 0.284231f
C3 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.55251f
C4 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.07164f
C5 a_13842_27148# VPWR 0.471462f
C6 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.433299f
C7 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.CEO 0.432008f
C8 a_5130_32076# VPWR 0.436368f
C9 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y a_17750_41000# 0.114097f
C10 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C11 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VPWR 1.77562f
C12 a_5130_28204# VPWR 0.361706f
C13 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.267144f
C14 SUNSAR_SAR8B_CV_0.XA5.CEO VPWR 1.0603f
C15 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C16 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y uo_out[3] 0.309657f
C17 SUNSAR_CAPT8B_CV_0.XF11.QN uo_out[3] 0.267395f
C18 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR 0.112858f
C19 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VPWR 2.95307f
C20 SUNSAR_CAPT8B_CV_0.XB07.QN VPWR 0.901622f
C21 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VPWR 0.452478f
C22 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y a_6302_42408# 0.113479f
C23 a_5130_35068# VPWR 0.394528f
C24 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.158152f
C25 a_15230_41352# VPWR 0.394053f
C26 a_5130_35948# VPWR 0.417826f
C27 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 3.57448f
C28 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_3762_35420# 0.133834f
C29 a_3762_32076# VPWR 0.436368f
C30 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP0.D VPWR 0.106927f
C31 a_3762_28204# VPWR 0.36179f
C32 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.702226f
C33 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C34 SUNSAR_SAR8B_CV_0.XA4.ENO a_12690_28556# 0.132757f
C35 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA4.Y 0.504864f
C36 a_10190_42760# SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.111734f
C37 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C38 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VPWR 0.723728f
C39 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y uo_out[3] 0.249907f
C40 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR 4.24834f
C41 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VPWR 1.77562f
C42 SUNSAR_CAPT8B_CV_0.XA2.MN0.G VPWR 0.667429f
C43 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.145483f
C44 a_10190_40648# VPWR 0.492624f
C45 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.57155f
C46 a_3762_35068# VPWR 0.394528f
C47 a_20270_41880# SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.100592f
C48 a_13862_41352# VPWR 0.394053f
C49 a_3762_35948# VPWR 0.417826f
C50 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35420# 0.160931f
C51 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C52 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.327909f
C53 uo_out[6] uo_out[7] 2.38922f
C54 SUNSAR_SAR8B_CV_0.XA4.CEO VPWR 2.30385f
C55 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.QN 0.318734f
C56 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.M3.G 0.263588f
C57 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP0.D VPWR 0.106927f
C58 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.D VPWR 0.104609f
C59 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.112859f
C60 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.449584f
C61 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_3728# 0.172147f
C62 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.589705f
C63 a_8822_40648# VPWR 0.491225f
C64 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.55251f
C65 SUNSAR_SAR8B_CV_0.XA7.XA8.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C66 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VPWR 0.271482f
C67 a_10170_27148# VPWR 0.470364f
C68 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.98135f
C69 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.375196f
C70 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA11.Y 0.220689f
C71 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VPWR 0.618979f
C72 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6519f
C73 a_5150_42760# VPWR 0.391454f
C74 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VPWR 0.429492f
C75 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.74594f
C76 SUNSAR_SAR8B_CV_0.XA3.ENO a_11322_28556# 0.135353f
C77 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C78 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.09966f
C79 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VPWR 0.720133f
C80 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G 0.22339f
C81 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.11263f
C82 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VPWR 0.519052f
C83 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.145483f
C84 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.ENO 0.409858f
C85 a_8802_27148# VPWR 0.471462f
C86 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.294852f
C87 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.437693f
C88 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 0.595738f
C89 SUNSAR_SAR8B_CV_0.XA20.XA10.B VPWR 1.13456f
C90 SUNSAR_SAR8B_CV_0.XA4.XA6.Y SUNSAR_SAR8B_CV_0.XA4.XA8.A 0.527529f
C91 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR 0.324111f
C92 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y a_16382_41000# 0.115667f
C93 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.DONE 0.372578f
C94 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR 0.137646f
C95 a_3782_42760# VPWR 0.391454f
C96 a_20270_44168# VPWR 0.340085f
C97 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.204048f
C98 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.17528f
C99 SUNSAR_SAR8B_CV_0.XA3.CEO VPWR 1.06031f
C100 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C101 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y a_13862_41000# 0.15757f
C102 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR 4.25569f
C103 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VPWR 1.77562f
C104 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.112859f
C105 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y a_2630_42408# 0.111909f
C106 a_16542_4918# VPWR 0.470354f
C107 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.449584f
C108 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.41635f
C109 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VPWR 2.1352f
C110 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.26537f
C111 a_10190_41352# VPWR 0.394053f
C112 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.377598f
C113 SUNSAR_CAPT8B_CV_0.XH13.QN uo_out[1] 0.254135f
C114 SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR 0.774301f
C115 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.746324f
C116 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VPWR 2.30036f
C117 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y a_15230_41000# 0.156079f
C118 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C119 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VPWR 1.06002f
C120 a_18902_44168# VPWR 0.3405f
C121 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.748719f
C122 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C123 a_8822_42760# SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.113305f
C124 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VPWR 0.723762f
C125 VPWR uo_out[7] 1.27659f
C126 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.297363f
C127 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y a_12710_41000# 0.114097f
C128 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.310451f
C129 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.11263f
C130 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.649845f
C131 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.145483f
C132 a_5150_40648# VPWR 0.492592f
C133 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y uo_out[1] 0.305961f
C134 SUNSAR_SAR8B_CV_0.XA6.DONE VPWR 0.246222f
C135 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.ENO 0.144331f
C136 a_20250_30316# VPWR 0.403745f
C137 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.268769f
C138 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233744f
C139 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C140 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.383512f
C141 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.744161f
C142 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.437693f
C143 a_8822_41352# VPWR 0.394053f
C144 SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR 0.780003f
C145 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VPWR 2.31184f
C146 SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR 9.39958f
C147 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR 0.138148f
C148 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y uo_out[7] 0.308722f
C149 SUNSAR_SAR8B_CV_0.XA2.CEO VPWR 2.30393f
C150 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.19724f
C151 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.426291f
C152 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.15234f
C153 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.112859f
C154 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VPWR 0.519052f
C155 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.744161f
C156 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_4688# 0.172147f
C157 a_3782_40648# VPWR 0.491225f
C158 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y uo_out[1] 0.248461f
C159 SUNSAR_SAR8B_CV_0.XA5.DONE VPWR 0.245452f
C160 a_18882_30316# VPWR 0.403802f
C161 a_5130_27148# VPWR 0.470364f
C162 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.649845f
C163 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA11.Y 0.293159f
C164 SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR 0.779986f
C165 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VPWR 2.31184f
C166 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.55251f
C167 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.165965f
C168 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.136678f
C169 SUNSAR_SAR8B_CV_0.EN VPWR 41.9239f
C170 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VPWR 1.06875f
C171 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C172 SUNSAR_SAR8B_CV_0.XA2.ENO a_7650_28556# 0.132757f
C173 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y uo_out[7] 0.248979f
C174 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VPWR 0.720114f
C175 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80606f
C176 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.D VPWR 0.104609f
C177 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y uo_out[5] 0.245678f
C178 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.340491f
C179 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.11263f
C180 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VPWR 0.452478f
C181 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.145483f
C182 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.ENO 0.438277f
C183 VPWR uo_out[6] 1.34623f
C184 SUNSAR_SAR8B_CV_0.XA4.DONE VPWR 0.246222f
C185 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.2165f
C186 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.12241f
C187 a_3762_27148# VPWR 0.471462f
C188 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.SARP 0.435464f
C189 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D 0.252966f
C190 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.CEO 0.432008f
C191 SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR 0.780003f
C192 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.625035f
C193 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VPWR 2.31184f
C194 a_23942_43112# VPWR 0.393308f
C195 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR 0.137646f
C196 a_15230_44168# VPWR 0.340085f
C197 SUNSAR_SAR8B_CV_0.XA1.CEO VPWR 1.0603f
C198 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.665724f
C199 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.242472f
C200 SUNSAR_SAR8B_CV_0.DONE VPWR 7.82915f
C201 ui_in[0] clk 0.169609f
C202 SUNSAR_SAR8B_CV_0.XA3.DONE VPWR 0.245452f
C203 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.297144f
C204 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.07223f
C205 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA0.XA11.Y 0.158152f
C206 SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR 0.779986f
C207 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VPWR 2.31184f
C208 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VPWR 1.05322f
C209 a_13862_44168# VPWR 0.3405f
C210 SUNSAR_SAR8B_CV_0.XA1.ENO a_6282_28556# 0.135353f
C211 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.441867f
C212 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VPWR 0.728492f
C213 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y a_11342_41000# 0.115667f
C214 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR 0.112858f
C215 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARP 0.506551f
C216 a_9990_4918# VPWR 0.468783f
C217 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.145483f
C218 a_23942_41000# VPWR 0.390551f
C219 SUNSAR_SAR8B_CV_0.XA2.DONE VPWR 0.246222f
C220 a_15210_30316# VPWR 0.404384f
C221 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.55251f
C222 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.276413f
C223 SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR 0.780003f
C224 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VPWR 2.31184f
C225 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR 0.138148f
C226 SUNSAR_SAR8B_CV_0.XA0.CEO VPWR 2.30575f
C227 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.34383f
C228 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y a_10190_41000# 0.156079f
C229 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR 0.112858f
C230 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.D VPWR 0.104609f
C231 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C232 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.40569f
C233 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_5648# 0.172147f
C234 SUNSAR_SAR8B_CV_0.XA1.DONE VPWR 0.245452f
C235 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.ENO 0.144331f
C236 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35068# 0.129098f
C237 a_13842_30316# VPWR 0.404384f
C238 a_20250_27500# VPWR 0.382397f
C239 SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR 0.779986f
C240 SUNSAR_SAR8B_CV_0.XA3.XA6.Y SUNSAR_SAR8B_CV_0.XA3.XA8.A 0.527529f
C241 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S 0.300065f
C242 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VPWR 2.31184f
C243 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.55251f
C244 SUNSAR_CAPT8B_CV_0.XI14.XA4.A VPWR 1.63909f
C245 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VPWR 1.06875f
C246 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.107567f
C247 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.441867f
C248 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.39041f
C249 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR 4.2492f
C250 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VPWR 1.77562f
C251 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_2928# 0.105547f
C252 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.145483f
C253 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.ENO 0.503825f
C254 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.86675f
C255 SUNSAR_SAR8B_CV_0.XA0.DONE VPWR 0.247527f
C256 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.12241f
C257 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C258 a_18882_27500# VPWR 0.382189f
C259 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.D 0.152518f
C260 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C261 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.D<5> 0.393076f
C262 SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR 0.784656f
C263 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 0.625175f
C264 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VPWR 2.31184f
C265 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.109613f
C266 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR 0.137646f
C267 a_20250_37180# VPWR 0.469114f
C268 a_22790_42408# SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.10248f
C269 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.11641f
C270 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VPWR 2.9531f
C271 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C272 a_16542_5270# VPWR 0.489055f
C273 a_20270_41000# VPWR 0.388156f
C274 a_23922_35420# VPWR 0.416528f
C275 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.671839f
C276 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA3.Y 0.432466f
C277 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.375025f
C278 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.284482f
C279 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.649845f
C280 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y a_5150_41880# 0.100592f
C281 a_23922_36300# VPWR 0.472384f
C282 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VPWR 4.6743f
C283 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.63636f
C284 uo_out[5] uo_out[4] 1.16362f
C285 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VPWR 1.05322f
C286 SUNSAR_SAR8B_CV_0.XA0.ENO a_2610_28556# 0.132757f
C287 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.131536f
C288 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.109137f
C289 a_18882_37180# VPWR 0.473682f
C290 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA2.Y 0.63636f
C291 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.143675f
C292 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.152052f
C293 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR 0.765792f
C294 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.145483f
C295 a_18902_41000# VPWR 0.388256f
C296 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.ENO 0.144331f
C297 a_10170_30316# VPWR 0.404384f
C298 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 54.2165f
C299 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.D 0.150467f
C300 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.744161f
C301 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C302 a_15230_41880# SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.100592f
C303 SUNSAR_SAR8B_CV_0.EN a_20250_29612# 0.142592f
C304 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.16676f
C305 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR 0.138148f
C306 SUNSAR_CAPT8B_CV_0.XH13.XA4.A VPWR 1.63909f
C307 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189112f
C308 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.52234f
C309 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR 4.27988f
C310 a_21422_42408# SUNSAR_CAPT8B_CV_0.XI14.XA3.Y 0.113479f
C311 a_13862_43288# VPWR 0.394205f
C312 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.144778f
C313 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.180903f
C314 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.339883f
C315 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_6608# 0.172147f
C316 VPWR uo_out[3] 1.25759f
C317 a_8802_30316# VPWR 0.404384f
C318 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.372599f
C319 a_15210_27500# VPWR 0.382397f
C320 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.587991f
C321 SUNSAR_SAR8B_CV_0.EN a_18882_29612# 0.143959f
C322 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.137975f
C323 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.393665f
C324 a_20250_32956# VPWR 0.433941f
C325 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.2165f
C326 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C327 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.45828f
C328 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VPWR 1.06875f
C329 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.143023f
C330 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA4.Y 0.107823f
C331 SUNSAR_SAR8B_CV_0.SARP VPWR 0.139564f
C332 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.139471f
C333 a_9990_5270# VPWR 0.490626f
C334 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_3888# 0.105547f
C335 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.ENO 0.438277f
C336 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.176792f
C337 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA10.Y 0.293873f
C338 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1615f
C339 a_20250_35420# VPWR 0.39661f
C340 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35068# 0.127528f
C341 a_13842_27500# VPWR 0.382189f
C342 a_20250_36300# VPWR 0.395776f
C343 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.625035f
C344 SUNSAR_SAR8B_CV_0.XA2.XA6.Y SUNSAR_SAR8B_CV_0.XA2.XA8.A 0.527529f
C345 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.241356f
C346 a_18882_32956# VPWR 0.436368f
C347 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.109613f
C348 SUNSAR_SAR8B_CV_0.XB2.XA3.B ua[0] 0.241597f
C349 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR 0.137646f
C350 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_3334# 0.120042f
C351 a_15210_37180# VPWR 0.474036f
C352 TIE_L1 uo_out[7] 0.461734f
C353 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VPWR 0.808658f
C354 a_15230_41000# VPWR 0.388156f
C355 a_18882_35420# VPWR 0.39968f
C356 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.791379f
C357 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.252047f
C358 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D 0.104122f
C359 a_18882_36300# VPWR 0.399161f
C360 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S ua[0] 0.100365f
C361 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VPWR 1.05322f
C362 SUNSAR_CAPT8B_CV_0.XG12.XA4.A VPWR 1.63909f
C363 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.110962f
C364 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_3334# 0.113134f
C365 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_OP 1.15994f
C366 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.142977f
C367 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.419738f
C368 a_13842_37180# VPWR 0.473697f
C369 a_10190_43288# VPWR 0.394205f
C370 a_20250_29612# VPWR 0.398044f
C371 a_23942_41880# VPWR 0.398828f
C372 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.154232f
C373 a_13862_41000# VPWR 0.388256f
C374 a_5130_30316# VPWR 0.404384f
C375 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 6.86675f
C376 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.11884f
C377 SUNSAR_SAR8B_CV_0.XB1.TIE_L ua[0] 1.05246f
C378 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C379 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.D 0.155821f
C380 SUNSAR_SAR8B_CV_0.EN a_15210_29612# 0.143959f
C381 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.D<6> 0.39306f
C382 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.105016f
C383 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C384 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR 0.138148f
C385 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.133602f
C386 a_17750_42408# SUNSAR_CAPT8B_CV_0.XH13.XA3.Y 0.111909f
C387 a_8822_43288# VPWR 0.394205f
C388 a_18882_29612# VPWR 0.397362f
C389 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.3401f
C390 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C391 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.ENO 0.144331f
C392 a_3762_30316# VPWR 0.404384f
C393 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C394 SUNSAR_SAR8B_CV_0.XB1.TIE_L ua[1] 0.704356f
C395 a_10170_27500# VPWR 0.382397f
C396 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON a_20250_30316# 0.127528f
C397 SUNSAR_SAR8B_CV_0.EN a_13842_29612# 0.143959f
C398 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_SAR8B_CV_0.D<6> 0.241356f
C399 a_15210_32956# VPWR 0.436368f
C400 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.86675f
C401 SUNSAR_SAR8B_CV_0.XB1.XA3.B ua[1] 0.241597f
C402 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VPWR 1.06875f
C403 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C404 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_2982# 0.158066f
C405 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.142956f
C406 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.419738f
C407 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR 0.112858f
C408 a_16542_5622# VPWR 0.472384f
C409 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_4848# 0.105547f
C410 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.ENO 0.503825f
C411 a_15210_35420# VPWR 0.39968f
C412 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6519f
C413 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03123f
C414 a_8802_27500# VPWR 0.382189f
C415 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.276413f
C416 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.D 0.150467f
C417 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.744161f
C418 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C419 a_15210_36300# VPWR 0.398846f
C420 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 0.625175f
C421 ua[1] ua[0] 3.85017f
C422 a_13842_32956# VPWR 0.436368f
C423 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S ua[1] 0.100365f
C424 a_23922_28556# VPWR 0.499441f
C425 SUNSAR_CAPT8B_CV_0.XF11.XA4.A VPWR 1.63909f
C426 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.133602f
C427 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.118152f
C428 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.10225f
C429 a_10170_37180# VPWR 0.474068f
C430 a_16382_42408# SUNSAR_CAPT8B_CV_0.XG12.XA3.Y 0.113479f
C431 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR 0.112858f
C432 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.ENO 0.793076f
C433 a_20270_41880# VPWR 0.395781f
C434 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C435 a_10190_41000# VPWR 0.388175f
C436 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA10.Y 0.381914f
C437 a_13842_35420# VPWR 0.39968f
C438 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35068# 0.129098f
C439 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VPWR 6.88568f
C440 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C441 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.62595f
C442 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON a_18882_30316# 0.129098f
C443 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.200058f
C444 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.12241f
C445 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.11099f
C446 a_13842_36300# VPWR 0.399161f
C447 VPWR uo_out[1] 1.02322f
C448 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.170578f
C449 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.142977f
C450 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.301485f
C451 a_8802_37180# VPWR 0.473729f
C452 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR 4.24508f
C453 a_5150_43288# VPWR 0.394205f
C454 a_18902_41880# VPWR 0.395781f
C455 a_15210_29612# VPWR 0.397362f
C456 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_2768# 0.172147f
C457 a_16542_5974# VPWR 0.449888f
C458 SUNSAR_CAPT8B_CV_0.XC08.XA4.A a_5150_42760# 0.111734f
C459 a_8822_41000# VPWR 0.388256f
C460 TIE_L1 VPWR 0.115195f
C461 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.ENO 0.144331f
C462 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 27.1615f
C463 a_23922_30844# VPWR 0.425847f
C464 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03123f
C465 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C466 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C467 SUNSAR_SAR8B_CV_0.EN a_10170_29612# 0.143959f
C468 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_SAR8B_CV_0.EN 0.176398f
C469 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA2.Y 0.432466f
C470 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.180455f
C471 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.241356f
C472 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.189429f
C473 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.133602f
C474 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.166192f
C475 a_3782_43288# VPWR 0.394205f
C476 a_13842_29612# VPWR 0.397362f
C477 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.290432f
C478 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.18612f
C479 a_5130_27500# VPWR 0.382397f
C480 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.284482f
C481 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D 0.104122f
C482 SUNSAR_SAR8B_CV_0.EN a_8802_29612# 0.143959f
C483 SUNSAR_SAR8B_CV_0.XA1.XA6.Y SUNSAR_SAR8B_CV_0.XA1.XA8.A 0.527529f
C484 TIE_L uo_out[5] 1.32477f
C485 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.393049f
C486 a_10170_32956# VPWR 0.436368f
C487 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 27.1615f
C488 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARN 0.64474f
C489 SUNSAR_CAPT8B_CV_0.XE10.XA4.A VPWR 1.63909f
C490 a_20250_28556# VPWR 0.406628f
C491 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.191868f
C492 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.11826f
C493 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.379175p
C494 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_2982# 0.158066f
C495 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.166272f
C496 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.142956f
C497 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.155424f
C498 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.146492f
C499 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_5808# 0.105547f
C500 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VPWR 0.808658f
C501 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.ENO 0.434116f
C502 a_10170_35420# VPWR 0.39968f
C503 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.55251f
C504 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VPWR 2.45124f
C505 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 1.03107f
C506 a_3762_27500# VPWR 0.382189f
C507 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.D 0.155821f
C508 a_10170_36300# VPWR 0.398846f
C509 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.08082f
C510 a_8802_32956# VPWR 0.436368f
C511 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.137745f
C512 a_18882_28556# VPWR 0.406628f
C513 SUNSAR_SAR8B_CV_0.XA20.XA2.CO a_23922_30844# 0.100515f
C514 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.133602f
C515 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.B 0.26479f
C516 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.166192f
C517 a_5130_37180# VPWR 0.474051f
C518 TIE_L2 uo_out[7] 0.106093f
C519 a_12710_42408# SUNSAR_CAPT8B_CV_0.XF11.XA3.Y 0.111909f
C520 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR 4.25322f
C521 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.ENO 1.2771f
C522 a_15230_41880# VPWR 0.395781f
C523 a_5150_41000# VPWR 0.388161f
C524 a_8802_35420# VPWR 0.39968f
C525 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARN 0.538639f
C526 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VPWR 2.44986f
C527 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON a_15210_30316# 0.127528f
C528 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.474658f
C529 a_8802_36300# VPWR 0.399161f
C530 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.412143f
C531 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.162703f
C532 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C533 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3334# 0.163985f
C534 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_3334# 0.114704f
C535 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.669708f
C536 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.166272f
C537 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.142977f
C538 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.449584f
C539 a_3762_37180# VPWR 0.473713f
C540 SUNSAR_CAPT8B_CV_0.XA3.Y VPWR 0.86364f
C541 a_13862_41880# VPWR 0.395781f
C542 a_10170_29612# VPWR 0.397362f
C543 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.152052f
C544 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_3728# 0.172147f
C545 a_9990_5622# VPWR 0.470814f
C546 a_3782_41000# VPWR 0.388256f
C547 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA10.Y 0.303978f
C548 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35068# 0.127528f
C549 SUNSAR_SAR8B_CV_0.XA20.XA10.A SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.321724f
C550 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6519f
C551 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VPWR 2.45309f
C552 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.791351f
C553 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C554 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.106828f
C555 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.D 0.150467f
C556 SUNSAR_SAR8B_CV_0.SARN ua[0] 1.02347f
C557 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.432466f
C558 SUNSAR_SAR8B_CV_0.EN a_5130_29612# 0.143959f
C559 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.CKN 0.102131f
C560 SUNSAR_CAPT8B_CV_0.XD09.XA4.A VPWR 1.63909f
C561 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON 0.133602f
C562 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_3334# 0.118471f
C563 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.166192f
C564 a_11342_42408# SUNSAR_CAPT8B_CV_0.XE10.XA3.Y 0.113479f
C565 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.545186f
C566 a_23942_43640# VPWR 0.412992f
C567 a_8802_29612# VPWR 0.397362f
C568 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.339883f
C569 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C570 SUNSAR_SAR8B_CV_0.EN ui_in[0] 0.969482f
C571 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.13078f
C572 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.ENO 0.144331f
C573 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VPWR 2.45309f
C574 a_20250_27852# VPWR 0.358413f
C575 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON a_13842_30316# 0.129098f
C576 TIE_L uo_out[2] 0.162449f
C577 SUNSAR_SAR8B_CV_0.SARN ua[1] 0.806872f
C578 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA1.Y 0.12241f
C579 SUNSAR_SAR8B_CV_0.EN a_3762_29612# 0.143959f
C580 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.199516f
C581 a_5130_32956# VPWR 0.436368f
C582 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6519f
C583 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.175642f
C584 a_15210_28556# VPWR 0.406628f
C585 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.105035f
C586 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.206912f
C587 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.142956f
C588 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.449584f
C589 a_16542_2630# VPWR 0.448659f
C590 TIE_L uo_out[4] 0.333172f
C591 SUNSAR_SAR8B_CV_0.XA7.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C592 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR 0.112858f
C593 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.724217f
C594 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y a_3782_41000# 0.15757f
C595 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG m3_18054_6768# 0.105547f
C596 a_9990_5974# VPWR 0.451043f
C597 a_23942_41352# VPWR 0.376408f
C598 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.ENO 0.491653f
C599 a_5130_35420# VPWR 0.39968f
C600 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.55251f
C601 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VPWR 2.45309f
C602 a_18882_27852# VPWR 0.358599f
C603 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.449584f
C604 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_4390# 0.15559f
C605 a_5130_36300# VPWR 0.398846f
C606 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.20727f
C607 SUNSAR_SAR8B_CV_0.XA0.XA6.Y SUNSAR_SAR8B_CV_0.XA0.XA8.A 0.527529f
C608 a_3762_32956# VPWR 0.436368f
C609 SUNSAR_SAR8B_CV_0.DONE ui_in[0] 0.175856f
C610 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C611 a_13842_28556# VPWR 0.406628f
C612 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON 0.133602f
C613 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_4038# 0.135393f
C614 a_20250_37532# VPWR 0.454392f
C615 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y 0.342913f
C616 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR 0.112858f
C617 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.ENO 1.2771f
C618 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y a_2630_41000# 0.114097f
C619 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C620 a_23922_26796# VPWR 0.442318f
C621 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA10.Y 0.352238f
C622 a_3762_35420# VPWR 0.39968f
C623 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VPWR 2.45309f
C624 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.TIE_L 4.28648f
C625 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D 0.104122f
C626 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_4390# 0.15559f
C627 a_3762_36300# VPWR 0.399161f
C628 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.215251f
C629 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.205884f
C630 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.393063f
C631 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y clk 0.210661f
C632 SUNSAR_CAPT8B_CV_0.XC08.XA4.A VPWR 1.63909f
C633 SUNSAR_SAR8B_CV_0.XB2.M3.G a_13950_3686# 0.16579f
C634 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.432466f
C635 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3334# 0.163985f
C636 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.142977f
C637 a_18882_37532# VPWR 0.458267f
C638 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y SUNSAR_SAR8B_CV_0.D<3> 0.241356f
C639 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP0.D VPWR 0.106927f
C640 a_5130_29612# VPWR 0.397362f
C641 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.722427f
C642 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.154232f
C643 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_4688# 0.172147f
C644 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.A 0.111867f
C645 TIE_L2 VPWR 0.106973f
C646 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.ENO 0.144331f
C647 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VPWR 2.45309f
C648 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.55251f
C649 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.10132f
C650 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.791379f
C651 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.276413f
C652 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.D 0.155821f
C653 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.449584f
C654 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[0] 0.247314f
C655 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.178111f
C656 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.241356f
C657 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18344f
C658 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VPWR 4.93712f
C659 VPWR ui_in[0] 1.38894f
C660 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON 0.133602f
C661 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.183415f
C662 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA1.Y 0.12241f
C663 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_22790_43640# 0.127669f
C664 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.D<3> 0.393049f
C665 a_7670_42408# SUNSAR_CAPT8B_CV_0.XD09.XA3.Y 0.111909f
C666 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR 3.09787f
C667 a_3762_29612# VPWR 0.397362f
C668 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.3401f
C669 a_20270_41352# VPWR 0.394053f
C670 SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.D VPWR 0.106794f
C671 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35068# 0.129098f
C672 SUNSAR_SAR8B_CV_0.XA6.XA8.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.143554f
C673 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VPWR 2.45309f
C674 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.34399f
C675 a_15210_27852# VPWR 0.358413f
C676 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON a_10170_30316# 0.127528f
C677 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.CKN 0.102131f
C678 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.12241f
C679 a_23922_36652# VPWR 0.449853f
C680 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.50324f
C681 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.EN 0.315968f
C682 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.55549f
C683 a_23922_33132# VPWR 0.415713f
C684 a_10170_28556# VPWR 0.406628f
C685 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C686 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.26479f
C687 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C688 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.4271f
C689 SUNSAR_SAR8B_CV_0.XA6.XA10.Y SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C690 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.103734f
C691 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.722417f
C692 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.QN 0.318734f
C693 a_20250_26796# VPWR 0.441753f
C694 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.ENO 0.11341f
C695 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.182408f
C696 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 54.2165f
C697 SUNSAR_SAR8B_CV_0.XA20.XA10.A VPWR 0.658328f
C698 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.193518f
C699 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.209352f
C700 a_13842_27852# VPWR 0.358599f
C701 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.204048f
C702 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.D 0.150467f
C703 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA2.Y 0.432466f
C704 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_34540# 0.103065f
C705 a_8802_28556# VPWR 0.406628f
C706 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON 0.133602f
C707 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.XA3.B 0.379175p
C708 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.669708f
C709 a_9990_2630# VPWR 0.447504f
C710 a_15210_37532# VPWR 0.459479f
C711 a_20250_34716# VPWR 0.396749f
C712 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.ENO 1.2771f
C713 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR 0.337652f
C714 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.CO 1.43919f
C715 a_23942_44344# VPWR 0.342053f
C716 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.DONE 0.492001f
C717 a_18882_26796# VPWR 0.442908f
C718 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA6.Y 0.291229f
C719 a_20250_31196# VPWR 0.437f
C720 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.238862f
C721 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.284482f
C722 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON a_8802_30316# 0.129098f
C723 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[5] 0.248535f
C724 TIE_L uo_out[0] 0.280844f
C725 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB2.M3.G 0.151329f
C726 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 1.62434f
C727 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VPWR 0.718455f
C728 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.228326f
C729 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.205884f
C730 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C731 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR 2.66621f
C732 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.175642f
C733 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.Y 0.178114f
C734 SUNSAR_SAR8B_CV_0.XB1.M3.G a_12582_3686# 0.16579f
C735 a_16542_2982# VPWR 0.490338f
C736 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C737 a_13842_37532# VPWR 0.458324f
C738 SUNSAR_SAR8B_CV_0.XA5.XA10.Y SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C739 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y a_10190_41880# 0.100592f
C740 a_18882_34716# VPWR 0.399819f
C741 a_23922_29964# VPWR 0.429137f
C742 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.233892f
C743 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.722427f
C744 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_5648# 0.172147f
C745 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA10.Y 0.303978f
C746 SUNSAR_SAR8B_CV_0.XA7.XA8.A VPWR 1.20972f
C747 SUNSAR_CAPT8B_CV_0.XG12.QN uo_out[2] 0.254418f
C748 a_18882_31196# VPWR 0.44007f
C749 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.55251f
C750 SUNSAR_SAR8B_CV_0.XA7.XA11.MP0.D VPWR 0.101562f
C751 SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR 2.64055f
C752 SUNSAR_SAR8B_CV_0.XB2.M3.G ua[0] 0.765539f
C753 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.143148f
C754 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.12241f
C755 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C756 SUNSAR_SAR8B_CV_0.D<0> VPWR 5.48841f
C757 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.13078f
C758 SUNSAR_SAR8B_CV_0.XA7.XA11.Y a_21402_36828# 0.104051f
C759 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VPWR 0.924613f
C760 a_10170_27852# VPWR 0.358413f
C761 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.126354f
C762 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.SARP 0.122781f
C763 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.238636f
C764 SUNSAR_SAR8B_CV_0.XA6.XA11.MP0.D VPWR 0.119314f
C765 SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR 2.64054f
C766 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C767 a_5130_28556# VPWR 0.406628f
C768 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.SARP 0.147435f
C769 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA2.Y 0.432466f
C770 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.40569f
C771 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y uo_out[0] 0.245915f
C772 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.722417f
C773 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.QN 0.318734f
C774 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.DONE 0.297507f
C775 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.D VPWR 0.106927f
C776 SUNSAR_CAPT8B_CV_0.XA4.Y clk 0.206733f
C777 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 6.86675f
C778 SUNSAR_SAR8B_CV_0.XA6.XA8.A VPWR 1.22023f
C779 SUNSAR_SAR8B_CV_0.XA5.XA8.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.145738f
C780 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35068# 0.127528f
C781 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D SUNSAR_SAR8B_CV_0.SARN 0.253395f
C782 a_8802_27852# VPWR 0.358599f
C783 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C784 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.XB1.M3.G 0.1501f
C785 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VPWR 0.725614f
C786 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C787 SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR 2.64055f
C788 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.11536f
C789 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[4] 0.249063f
C790 a_3762_28556# VPWR 0.406628f
C791 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.179089f
C792 SUNSAR_CAPT8B_CV_0.XA4.MN0.S SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.138433f
C793 a_10170_37532# VPWR 0.459599f
C794 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.D<4> 0.393055f
C795 a_15210_34716# VPWR 0.399819f
C796 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y uo_out[0] 0.307374f
C797 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.D VPWR 0.108436f
C798 a_5150_42408# VPWR 0.391292f
C799 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C800 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C801 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP0.D VPWR 0.106927f
C802 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA10.Y 0.352238f
C803 a_15210_31196# VPWR 0.44007f
C804 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C805 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON a_5130_30316# 0.127528f
C806 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VPWR 0.722887f
C807 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.228332f
C808 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA6.Y 0.205884f
C809 SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR 2.64054f
C810 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP 0.123668f
C811 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31666f
C812 a_8802_37532# VPWR 0.458443f
C813 SUNSAR_SAR8B_CV_0.XA4.XA10.Y SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C814 SUNSAR_SAR8B_CV_0.XA7.XA10.Y a_21402_36300# 0.13402f
C815 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_SAR8B_CV_0.D<4> 0.241356f
C816 a_13842_34716# VPWR 0.399819f
C817 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y uo_out[2] 0.246879f
C818 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VPWR 0.279205f
C819 a_3782_42408# VPWR 0.391292f
C820 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.63636f
C821 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.152052f
C822 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.738812f
C823 SUNSAR_SAR8B_CV_0.XB1.XA3.B m3_2358_6608# 0.172147f
C824 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_2928# 0.105547f
C825 SUNSAR_SAR8B_CV_0.D<1> VPWR 5.18522f
C826 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VPWR 0.930839f
C827 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_21402_35420# 0.160931f
C828 SUNSAR_CAPT8B_CV_0.XI14.QN uo_out[0] 0.25785f
C829 a_13842_31196# VPWR 0.44007f
C830 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.2165f
C831 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.791351f
C832 TIE_L clk 0.150303f
C833 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C834 SUNSAR_SAR8B_CV_0.XA5.XA11.MP0.D VPWR 0.101979f
C835 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.CKN 0.153964f
C836 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR 2.7271f
C837 SUNSAR_SAR8B_CV_0.XB1.M3.G ua[1] 0.762388f
C838 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_4038# 0.135393f
C839 a_9990_2982# VPWR 0.491909f
C840 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y uo_out[2] 0.305131f
C841 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.339883f
C842 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.280191f
C843 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.DONE 0.297715f
C844 SUNSAR_SAR8B_CV_0.XA4.XA8.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.143554f
C845 SUNSAR_SAR8B_CV_0.XA7.XA8.A a_20250_35420# 0.133834f
C846 a_5130_27852# VPWR 0.358413f
C847 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y uo_out[5] 0.30523f
C848 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON a_3762_30316# 0.129098f
C849 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.204048f
C850 SUNSAR_SAR8B_CV_0.XA4.XA11.MP0.D VPWR 0.119314f
C851 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C852 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR 2.72582f
C853 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y uo_out[4] 0.246349f
C854 a_20250_28908# VPWR 0.395394f
C855 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.178114f
C856 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.432466f
C857 a_16542_3334# VPWR 0.380282f
C858 SUNSAR_SAR8B_CV_0.XA3.XA10.Y SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C859 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y a_2630_42408# 0.100131f
C860 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.D VPWR 0.104609f
C861 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR 0.686731f
C862 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.738798f
C863 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.152045f
C864 SUNSAR_SAR8B_CV_0.XA6.XA11.Y a_17730_36828# 0.10248f
C865 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1615f
C866 SUNSAR_SAR8B_CV_0.XA5.XA8.A VPWR 1.2202f
C867 uo_out[7] uo_out[5] 1.57818f
C868 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.331207f
C869 a_3762_27852# VPWR 0.358599f
C870 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.276252f
C871 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_4742# 0.156331f
C872 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VPWR 0.725614f
C873 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR 2.72889f
C874 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y uo_out[4] 0.305131f
C875 a_18882_28908# VPWR 0.395394f
C876 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.464697f
C877 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.159359f
C878 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 0.635098f
C879 a_21422_43816# SUNSAR_CAPT8B_CV_0.XI14.QN 0.129239f
C880 a_5130_37532# VPWR 0.459538f
C881 a_10170_34716# VPWR 0.399819f
C882 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VPWR 0.898003f
C883 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C884 SUNSAR_SAR8B_CV_0.D<2> VPWR 5.20829f
C885 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VPWR 0.93081f
C886 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35068# 0.129098f
C887 a_10170_31196# VPWR 0.44007f
C888 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C889 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_4742# 0.156331f
C890 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.301485f
C891 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VPWR 0.722887f
C892 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.M3.G 0.36754f
C893 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.228326f
C894 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA6.Y 0.205884f
C895 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.GNG 0.250503f
C896 a_3762_37532# VPWR 0.458382f
C897 a_8802_34716# VPWR 0.399819f
C898 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.CK 1.59176f
C899 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.154232f
C900 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VPWR 0.898003f
C901 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.740872f
C902 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.DONE 0.297504f
C903 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_3888# 0.105547f
C904 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP0.D VPWR 0.106927f
C905 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA2.XA10.Y 0.303978f
C906 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C907 SUNSAR_SAR8B_CV_0.XA4.XA8.A VPWR 1.22023f
C908 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_18882_35420# 0.133834f
C909 a_8802_31196# VPWR 0.44007f
C910 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.86675f
C911 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.108751f
C912 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 3.86364f
C913 SUNSAR_SAR8B_CV_0.XA3.XA11.MP0.D VPWR 0.101979f
C914 a_20250_33836# VPWR 0.407174f
C915 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C916 uo_out[6] uo_out[5] 0.327382f
C917 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.179089f
C918 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.324243f
C919 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.CKN 0.41624f
C920 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.3401f
C921 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VPWR 0.898003f
C922 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C923 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.419738f
C924 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP0.D VPWR 0.106927f
C925 a_10190_41880# VPWR 0.395781f
C926 SUNSAR_SAR8B_CV_0.XA5.XA11.Y a_16362_36828# 0.104051f
C927 SUNSAR_SAR8B_CV_0.XA1.CEO SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.13078f
C928 a_17750_42408# SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.100131f
C929 SUNSAR_SAR8B_CV_0.XA6.XA8.A a_17730_35420# 0.160931f
C930 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_CAPT8B_CV_0.XA4.MN0.S 0.206292f
C931 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.204048f
C932 SUNSAR_SAR8B_CV_0.XA2.XA11.MP0.D VPWR 0.119314f
C933 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.CKN 0.153964f
C934 a_18882_33836# VPWR 0.409601f
C935 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.174995f
C936 a_15210_28908# VPWR 0.395394f
C937 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C938 SUNSAR_SAR8B_CV_0.XB2.M3.G SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D 0.101001f
C939 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.63636f
C940 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C941 a_23942_40296# VPWR 0.453754f
C942 SUNSAR_SAR8B_CV_0.XA2.XA10.Y SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C943 SUNSAR_SAR8B_CV_0.XA6.XA10.Y a_17730_36300# 0.13253f
C944 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y SUNSAR_SAR8B_CV_0.D<5> 0.241356f
C945 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VPWR 0.271482f
C946 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VPWR 0.898003f
C947 SUNSAR_SAR8B_CV_0.D<3> VPWR 5.17056f
C948 a_8822_41880# VPWR 0.395781f
C949 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6519f
C950 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VPWR 0.930839f
C951 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y uo_out[6] 0.251051f
C952 SUNSAR_SAR8B_CV_0.XA3.XA8.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.145738f
C953 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VPWR 2.95303f
C954 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C955 a_23942_42760# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.101843f
C956 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB1.M3.G 0.175967f
C957 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VPWR 0.725614f
C958 uo_out[7] uo_out[4] 0.121957f
C959 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.475004f
C960 a_13842_28908# VPWR 0.395394f
C961 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C962 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.CMP_ON 2.96993f
C963 a_17750_43816# SUNSAR_CAPT8B_CV_0.XH13.QN 0.127669f
C964 a_9990_3334# VPWR 0.380282f
C965 a_5130_34716# VPWR 0.399819f
C966 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VPWR 0.898003f
C967 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.DONE 0.297602f
C968 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.QN 0.318734f
C969 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.419738f
C970 SUNSAR_SAR8B_CV_0.XA0.CEO SUNSAR_SAR8B_CV_0.XA1.XA10.Y 0.352238f
C971 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C972 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y uo_out[6] 0.306905f
C973 a_5130_31196# VPWR 0.44007f
C974 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.118161f
C975 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.30776f
C976 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.SARP 0.257526f
C977 a_22790_42760# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.13379f
C978 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.301485f
C979 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VPWR 0.722887f
C980 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.228332f
C981 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA6.Y 0.205884f
C982 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C983 VPWR uo_out[5] 1.0281f
C984 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.178114f
C985 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C986 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA7.CN1 0.466806f
C987 SUNSAR_SAR8B_CV_0.XA1.XA10.Y SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C988 SUNSAR_SAR8B_CV_0.XA5.XA10.Y a_16362_36300# 0.13402f
C989 a_3762_34716# VPWR 0.399819f
C990 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA6.ENO 0.291697f
C991 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.D VPWR 0.104609f
C992 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VPWR 0.898003f
C993 SUNSAR_CAPT8B_CV_0.XA4.MN0.S clk 0.438597f
C994 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_4848# 0.105547f
C995 SUNSAR_SAR8B_CV_0.XA3.XA8.A VPWR 1.2202f
C996 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP0.D VPWR 0.106927f
C997 SUNSAR_SAR8B_CV_0.XA0.XA8.A a_2610_35068# 0.127528f
C998 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1615f
C999 a_3762_31196# VPWR 0.44007f
C1000 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.13041f
C1001 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S 0.128204f
C1002 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.ENO 0.116058f
C1003 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C1004 SUNSAR_SAR8B_CV_0.XA1.XA11.MP0.D VPWR 0.101979f
C1005 a_15210_33836# VPWR 0.409601f
C1006 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C1007 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XB1.CKN 0.143148f
C1008 a_16382_43816# SUNSAR_CAPT8B_CV_0.XG12.QN 0.129239f
C1009 a_20270_40296# VPWR 0.455248f
C1010 uo_out[6] uo_out[4] 0.84361f
C1011 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VPWR 0.271482f
C1012 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C1013 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VPWR 0.898003f
C1014 SUNSAR_SAR8B_CV_0.D<4> VPWR 5.15123f
C1015 a_5150_41880# VPWR 0.395781f
C1016 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VPWR 0.93081f
C1017 SUNSAR_SAR8B_CV_0.XA2.XA8.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.143554f
C1018 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VPWR 2.95305f
C1019 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.118161f
C1020 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.ENO 0.111173f
C1021 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.849501f
C1022 SUNSAR_SAR8B_CV_0.XA0.XA11.MP0.D VPWR 0.119314f
C1023 a_13842_33836# VPWR 0.409601f
C1024 a_10170_28908# VPWR 0.395394f
C1025 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1026 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA6.CN1 0.466806f
C1027 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA1.Y 0.233892f
C1028 SUNSAR_SAR8B_CV_0.XB2.XA3.B VPWR 1.56028f
C1029 a_18902_40296# VPWR 0.457343f
C1030 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.42393f
C1031 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VPWR 3.91346f
C1032 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.26609f
C1033 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VPWR 0.898003f
C1034 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.DONE 0.297941f
C1035 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y 0.386305f
C1036 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP0.D VPWR 0.106927f
C1037 a_3782_41880# VPWR 0.395781f
C1038 SUNSAR_SAR8B_CV_0.XA4.XA11.Y a_12690_36828# 0.10248f
C1039 SUNSAR_SAR8B_CV_0.XA0.XA11.Y SUNSAR_SAR8B_CV_0.XB1.TIE_L 0.215804f
C1040 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.55251f
C1041 SUNSAR_SAR8B_CV_0.XA2.XA8.A VPWR 1.22023f
C1042 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VPWR 1.77562f
C1043 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_16362_35420# 0.160931f
C1044 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VPWR 6.94539f
C1045 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP 0.129613f
C1046 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S 0.363295f
C1047 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.ENO 0.111217f
C1048 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.ENO 0.893904f
C1049 a_12710_42408# SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.100131f
C1050 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VPWR 0.728421f
C1051 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1052 a_8802_28908# VPWR 0.395394f
C1053 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.179089f
C1054 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.30589f
C1055 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.CKN 0.200119f
C1056 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.437693f
C1057 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR 0.183853f
C1058 a_23922_34892# VPWR 0.395601f
C1059 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.432466f
C1060 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C1061 a_23942_42760# VPWR 0.388156f
C1062 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP0.D VPWR 0.106927f
C1063 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA1.Y 0.233892f
C1064 SUNSAR_CAPT8B_CV_0.XB07.XA4.A a_3782_42760# 0.113305f
C1065 a_10190_44168# VPWR 0.340085f
C1066 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP0.D VPWR 0.106927f
C1067 SUNSAR_SAR8B_CV_0.XA5.XA8.A a_15210_35420# 0.133834f
C1068 a_23922_31724# VPWR 0.412398f
C1069 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.118226f
C1070 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.ENO 0.111173f
C1071 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.ENO 0.952619f
C1072 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_5094# 0.160184f
C1073 VPWR uo_out[2] 1.02322f
C1074 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.301485f
C1075 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.227341f
C1076 SUNSAR_SAR8B_CV_0.XB1.TIE_L VPWR 7.37316f
C1077 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA6.Y 0.205884f
C1078 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA5.CN1 0.466806f
C1079 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.231927f
C1080 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D 0.101001f
C1081 SUNSAR_SAR8B_CV_0.XB1.XA3.B VPWR 1.5612f
C1082 SUNSAR_SAR8B_CV_0.XA0.XA10.Y SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C1083 VPWR uo_out[4] 1.03096f
C1084 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA3.Y 0.12241f
C1085 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.D VPWR 0.104609f
C1086 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.473354f
C1087 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.152052f
C1088 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_5808# 0.105547f
C1089 SUNSAR_SAR8B_CV_0.D<5> VPWR 5.14531f
C1090 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP0.D VPWR 0.118162f
C1091 a_8822_44168# VPWR 0.3405f
C1092 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VPWR 0.930839f
C1093 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6519f
C1094 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.530644f
C1095 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP 0.13041f
C1096 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 4.0111f
C1097 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.ENO 1.02916f
C1098 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.ENO 0.111217f
C1099 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C1100 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_5094# 0.160184f
C1101 a_10170_33836# VPWR 0.409601f
C1102 SUNSAR_SAR8B_CV_0.XA20.XA2.CO SUNSAR_SAR8B_CV_0.XA0.CMP_ON 0.504801f
C1103 VPWR ua[0] 0.51729f
C1104 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.CKN 0.41624f
C1105 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR 0.183853f
C1106 a_12710_43816# SUNSAR_CAPT8B_CV_0.XF11.QN 0.127669f
C1107 a_15230_40296# VPWR 0.455577f
C1108 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.55251f
C1109 SUNSAR_SAR8B_CV_0.XA7.ENO VPWR 4.77251f
C1110 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.149144f
C1111 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145339f
C1112 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.DONE 0.298165f
C1113 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y a_22790_41000# 0.11811f
C1114 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.386137f
C1115 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.QN 0.318734f
C1116 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.449584f
C1117 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VPWR 1.20019f
C1118 SUNSAR_SAR8B_CV_0.XA3.XA11.Y a_11322_36828# 0.104051f
C1119 SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR 2.62711f
C1120 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.118161f
C1121 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C1122 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.ENO 0.952619f
C1123 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.ENO 0.111173f
C1124 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.316693f
C1125 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.204048f
C1126 a_20250_36828# VPWR 0.392512f
C1127 a_8802_33836# VPWR 0.409601f
C1128 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.174845f
C1129 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.SARN 0.591428f
C1130 a_5130_28908# VPWR 0.395394f
C1131 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.178114f
C1132 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA4.CN1 0.466806f
C1133 VPWR ua[1] 0.225132f
C1134 SUNSAR_SAR8B_CV_0.XB1.M3.G SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 0.250503f
C1135 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_CAPT8B_CV_0.XH13.XA2.Y 0.63636f
C1136 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.437693f
C1137 a_16542_4038# VPWR 0.379979f
C1138 a_13862_40296# VPWR 0.457343f
C1139 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.232115f
C1140 SUNSAR_SAR8B_CV_0.XA4.XA10.Y a_12690_36300# 0.13253f
C1141 SUNSAR_SAR8B_CV_0.XA6.ENO VPWR 5.54203f
C1142 a_20270_42760# VPWR 0.391454f
C1143 a_15210_26796# VPWR 0.441753f
C1144 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.182595f
C1145 SUNSAR_SAR8B_CV_0.XA1.XA8.A VPWR 1.2202f
C1146 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 3.55251f
C1147 SUNSAR_SAR8B_CV_0.XA1.XA8.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C1148 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_13842_35420# 0.133834f
C1149 SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR 2.62329f
C1150 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP 0.129613f
C1151 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.2199f
C1152 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.ENO 1.02916f
C1153 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.ENO 0.111217f
C1154 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S 0.126806f
C1155 a_20270_42760# SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.111734f
C1156 a_18882_36828# VPWR 0.395703f
C1157 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.EN 0.343905f
C1158 a_3762_28908# VPWR 0.395394f
C1159 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.SARP 0.524159f
C1160 a_11342_43816# SUNSAR_CAPT8B_CV_0.XE10.QN 0.129239f
C1161 SUNSAR_SAR8B_CV_0.XA5.ENO VPWR 4.84607f
C1162 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C1163 a_18902_42760# VPWR 0.391454f
C1164 a_13842_26796# VPWR 0.442908f
C1165 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.SARN 0.108405f
C1166 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.449584f
C1167 SUNSAR_SAR8B_CV_0.D<6> VPWR 5.17441f
C1168 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP0.D VPWR 0.106927f
C1169 SUNSAR_CAPT8B_CV_0.XA4.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.104933f
C1170 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VPWR 0.93081f
C1171 SUNSAR_SAR8B_CV_0.XA4.XA8.A a_12690_35420# 0.160931f
C1172 SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR 2.62342f
C1173 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.118226f
C1174 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.398331f
C1175 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.ENO 0.952619f
C1176 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.ENO 0.111173f
C1177 uo_out[2] uo_out[3] 0.110956f
C1178 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_23922_29964# 0.151031f
C1179 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.301485f
C1180 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.227352f
C1181 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA6.Y 0.205884f
C1182 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C1183 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.CN1 0.466806f
C1184 a_23942_42408# VPWR 0.3915f
C1185 uo_out[3] uo_out[4] 0.862834f
C1186 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.726497f
C1187 SUNSAR_SAR8B_CV_0.XA3.XA10.Y a_11322_36300# 0.13402f
C1188 SUNSAR_SAR8B_CV_0.XA4.ENO VPWR 5.52623f
C1189 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VPWR 0.271482f
C1190 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.DONE 0.294651f
C1191 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y 0.375196f
C1192 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG m3_9126_6768# 0.105547f
C1193 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP0.D VPWR 0.106927f
C1194 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP0.D VPWR 0.106927f
C1195 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.XA11.Y 0.324105f
C1196 SUNSAR_SAR8B_CV_0.XA0.XA8.A VPWR 1.22398f
C1197 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.55251f
C1198 SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR 2.62342f
C1199 SUNSAR_SAR8B_CV_0.XB1.TIE_L SUNSAR_SAR8B_CV_0.SARP 0.596437f
C1200 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP 0.13041f
C1201 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.25689f
C1202 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.ENO 1.04628f
C1203 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.XA2.Y 0.63636f
C1204 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S 0.363295f
C1205 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR a_22770_29964# 0.134249f
C1206 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XF11.QN 0.318734f
C1207 TIE_L uo_out[7] 0.462706f
C1208 a_5130_33836# VPWR 0.409601f
C1209 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D 0.107674f
C1210 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA3.Y 0.134182f
C1211 a_10190_40296# VPWR 0.455675f
C1212 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.SARP 0.102632f
C1213 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 54.2165f
C1214 SUNSAR_SAR8B_CV_0.XA3.ENO VPWR 4.84607f
C1215 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C1216 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP0.D VPWR 0.106927f
C1217 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.107427f
C1218 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.QN 0.318734f
C1219 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA7.CEO 0.138f
C1220 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y a_8822_41000# 0.15757f
C1221 SUNSAR_SAR8B_CV_0.XA0.XA8.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C1222 SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR 2.62342f
C1223 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.118161f
C1224 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.79343f
C1225 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C1226 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.204048f
C1227 VPWR uo_out[0] 1.19196f
C1228 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.694484f
C1229 a_15210_36828# VPWR 0.395582f
C1230 a_3762_33836# VPWR 0.409601f
C1231 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.174995f
C1232 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.D VPWR 0.104609f
C1233 SUNSAR_CAPT8B_CV_0.XB07.XA4.A VPWR 1.63909f
C1234 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.535136f
C1235 SUNSAR_SAR8B_CV_0.XB2.XA1.Y SUNSAR_SAR8B_CV_0.XB2.M3.G 0.224309f
C1236 a_8822_40296# VPWR 0.457343f
C1237 SUNSAR_SAR8B_CV_0.XA2.ENO VPWR 5.52623f
C1238 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.D VPWR 0.104609f
C1239 a_15230_42760# VPWR 0.391454f
C1240 a_10170_26796# VPWR 0.441753f
C1241 SUNSAR_SAR8B_CV_0.D<7> VPWR 3.61291f
C1242 SUNSAR_SAR8B_CV_0.XA2.XA11.Y a_7650_36828# 0.10248f
C1243 SUNSAR_SAR8B_CV_0.XA6.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.158152f
C1244 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y a_7670_41000# 0.114097f
C1245 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 54.2173f
C1246 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VPWR 0.94014f
C1247 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR 2.62393f
C1248 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP 0.129613f
C1249 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_13950_5446# 0.102604f
C1250 a_18902_42760# SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.113305f
C1251 SUNSAR_SAR8B_CV_0.SARP ua[1] 1.01251f
C1252 a_13842_36828# VPWR 0.395703f
C1253 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.744161f
C1254 TIE_L1 uo_out[5] 0.366299f
C1255 a_20270_42408# VPWR 0.391292f
C1256 a_9990_4038# VPWR 0.379979f
C1257 TIE_L uo_out[6] 0.203535f
C1258 SUNSAR_SAR8B_CV_0.XA1.ENO VPWR 4.84607f
C1259 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VPWR 0.271482f
C1260 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.303428f
C1261 a_13862_42760# VPWR 0.391454f
C1262 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y SUNSAR_SAR8B_CV_0.D<7> 0.241356f
C1263 a_8802_26796# VPWR 0.442908f
C1264 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.233892f
C1265 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y 0.383512f
C1266 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP0.D VPWR 0.106927f
C1267 a_23922_35948# VPWR 0.390687f
C1268 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR 2.62403f
C1269 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.118226f
C1270 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.316693f
C1271 SUNSAR_SAR8B_CV_0.XB1.TIE_L a_12582_5446# 0.101033f
C1272 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y SUNSAR_CAPT8B_CV_0.XE10.XA4.A 0.301485f
C1273 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.638386f
C1274 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CP0 0.331282f
C1275 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA6.Y 0.205884f
C1276 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C1277 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_CAPT8B_CV_0.XB07.XA4.A 0.649845f
C1278 SUNSAR_SAR8B_CV_0.SARN VPWR 0.132799f
C1279 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.D VPWR 0.104609f
C1280 SUNSAR_CAPT8B_CV_0.XA4.Y VPWR 1.18734f
C1281 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.559553f
C1282 a_18902_42408# VPWR 0.391292f
C1283 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VPWR 2.50821f
C1284 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C1285 SUNSAR_SAR8B_CV_0.XA0.ENO VPWR 5.52718f
C1286 a_5150_44168# VPWR 0.340085f
C1287 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.244517f
C1288 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y SUNSAR_SAR8B_CV_0.D<7> 0.393125f
C1289 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.EN 0.208884f
C1290 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP0.D VPWR 0.106927f
C1291 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA6.XA11.Y 0.220689f
C1292 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_11322_35420# 0.160931f
C1293 SUNSAR_SAR8B_CV_0.XA7.XA6.Y SUNSAR_SAR8B_CV_0.XA7.XA8.A 0.527529f
C1294 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.55251f
C1295 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.394834f
C1296 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP 0.13041f
C1297 SUNSAR_SAR8B_CV_0.XA0.CMP_ON SUNSAR_SAR8B_CV_0.XA0.CMP_OP 7.93512f
C1298 SUNSAR_SAR8B_CV_0.XA20.XA1.CK a_22770_28556# 0.140127f
C1299 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S 0.126806f
C1300 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_CAPT8B_CV_0.XE10.QN 0.318734f
C1301 a_5150_43816# VPWR 0.391817f
C1302 SUNSAR_SAR8B_CV_0.XB2.CKN VPWR 2.34497f
C1303 a_5150_40296# VPWR 0.455605f
C1304 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 6.86675f
C1305 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C1306 a_20270_43816# VPWR 0.391817f
C1307 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C1308 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.386137f
C1309 SUNSAR_SAR8B_CV_0.XA1.XA11.Y a_6282_36828# 0.104051f
C1310 SUNSAR_SAR8B_CV_0.XA3.XA8.A a_10170_35420# 0.133834f
C1311 a_20250_32076# VPWR 0.433941f
C1312 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP 0.118161f
C1313 a_20250_28204# VPWR 0.361706f
C1314 a_10170_36828# VPWR 0.396003f
C1315 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C1316 a_3782_43816# VPWR 0.391817f
C1317 a_20270_43288# VPWR 0.394205f
C1318 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.649845f
C1319 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y SUNSAR_CAPT8B_CV_0.XG12.XA1.Y 0.63636f
C1320 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C1321 a_3782_40296# VPWR 0.457343f
C1322 TIE_L VPWR 0.401306f
C1323 SUNSAR_SAR8B_CV_0.XA2.XA10.Y a_7650_36300# 0.13253f
C1324 a_20250_35068# VPWR 0.391458f
C1325 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.D VPWR 0.104609f
C1326 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.18614f
C1327 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA2.CO 0.205975f
C1328 a_10190_42760# VPWR 0.391454f
C1329 a_18902_43816# VPWR 0.391817f
C1330 a_5130_26796# VPWR 0.441753f
C1331 SUNSAR_SAR8B_CV_0.XA5.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.377598f
C1332 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y a_6302_41000# 0.115667f
C1333 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 6.86675f
C1334 a_20250_35948# VPWR 0.414756f
C1335 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1336 a_18882_32076# VPWR 0.436368f
C1337 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 5.19722f
C1338 a_18882_28204# VPWR 0.36179f
C1339 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S 0.363295f
C1340 VPWR clk 0.645958f
C1341 a_7670_42408# SUNSAR_CAPT8B_CV_0.XD09.XA2.Y 0.100131f
C1342 a_8802_36828# VPWR 0.396052f
C1343 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VPWR 0.405511f
C1344 a_18902_43288# VPWR 0.394205f
C1345 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.CKN 0.200119f
C1346 a_15230_42408# VPWR 0.391292f
C1347 SUNSAR_SAR8B_CV_0.XA7.CEO SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.127551f
C1348 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARP 0.187721f
C1349 a_18882_35068# VPWR 0.394528f
C1350 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.145048f
C1351 a_8822_42760# VPWR 0.391454f
C1352 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.328435f
C1353 a_3762_26796# VPWR 0.442908f
C1354 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C1355 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP0.D VPWR 0.106927f
C1356 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y a_5150_41000# 0.156079f
C1357 a_18882_35948# VPWR 0.417826f
C1358 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y SUNSAR_CAPT8B_CV_0.XD09.XA4.A 0.301485f
C1359 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.327152f
C1360 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR 1.70987f
C1361 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR 11.751401f
C1362 a_13862_42408# VPWR 0.391292f
C1363 a_23942_40648# VPWR 0.489579f
C1364 SUNSAR_SAR8B_CV_0.XA1.XA10.Y a_6282_36300# 0.13402f
C1365 SUNSAR_SAR8B_CV_0.XA6.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.693521f
C1366 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP0.D VPWR 0.106927f
C1367 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.XA11.Y 0.293159f
C1368 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_8802_35420# 0.133834f
C1369 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.2165f
C1370 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VPWR 2.95296f
C1371 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y SUNSAR_CAPT8B_CV_0.XE10.XA1.Y 0.63636f
C1372 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C1373 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.SARP 5.22744f
C1374 a_15230_42760# SUNSAR_CAPT8B_CV_0.XG12.XA4.A 0.111734f
C1375 a_23942_43992# VPWR 0.388156f
C1376 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.D VPWR 0.104609f
C1377 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.649845f
C1378 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 27.1615f
C1379 SUNSAR_SAR8B_CV_0.XA5.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C1380 a_15230_43816# VPWR 0.391817f
C1381 a_23922_27148# VPWR 0.483246f
C1382 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.107427f
C1383 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA5.CEO 0.432008f
C1384 SUNSAR_SAR8B_CV_0.XA6.XA6.Y SUNSAR_SAR8B_CV_0.XA6.XA8.A 0.527529f
C1385 SUNSAR_SAR8B_CV_0.XA2.XA8.A a_7650_35420# 0.160931f
C1386 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y a_21422_41000# 0.115667f
C1387 a_15210_32076# VPWR 0.436368f
C1388 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VPWR 1.77563f
C1389 a_15210_28204# VPWR 0.361706f
C1390 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.316693f
C1391 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y 0.204048f
C1392 a_5130_36828# VPWR 0.395767f
C1393 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C1394 a_15230_43288# VPWR 0.394205f
C1395 TIE_L uo_out[3] 0.188109f
C1396 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y SUNSAR_CAPT8B_CV_0.XI14.XA4.A 0.744161f
C1397 SUNSAR_SAR8B_CV_0.XB1.CKN VPWR 2.34497f
C1398 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.787331f
C1399 a_15210_35068# VPWR 0.394528f
C1400 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VPWR 0.271482f
C1401 SUNSAR_SAR8B_CV_0.XA4.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C1402 a_13862_43816# VPWR 0.391817f
C1403 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y 0.375196f
C1404 SUNSAR_SAR8B_CV_0.XA4.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.158152f
C1405 SUNSAR_SAR8B_CV_0.XA0.XA11.Y a_2610_36828# 0.10248f
C1406 a_15210_35948# VPWR 0.417826f
C1407 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 27.1625f
C1408 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y a_20270_41000# 0.156079f
C1409 a_13842_32076# VPWR 0.436368f
C1410 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP0.D VPWR 0.106927f
C1411 a_13842_28204# VPWR 0.36179f
C1412 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON 0.702226f
C1413 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S 0.126806f
C1414 a_5150_41352# VPWR 0.394053f
C1415 a_3762_36828# VPWR 0.395857f
C1416 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.142061f
C1417 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR 4.36162f
C1418 SUNSAR_CAPT8B_CV_0.XI14.QN VPWR 0.901631f
C1419 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G SUNSAR_SAR8B_CV_0.XB2.XA1.Y 0.22339f
C1420 a_10190_42408# VPWR 0.391292f
C1421 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VPWR 2.50821f
C1422 a_20270_40648# VPWR 0.492579f
C1423 a_3782_44168# VPWR 0.3405f
C1424 a_13842_35068# VPWR 0.394528f
C1425 SUNSAR_SAR8B_CV_0.XA3.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C1426 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP0.D VPWR 0.106927f
C1427 a_13842_35948# VPWR 0.417826f
C1428 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1429 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C1430 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.15651f
C1431 a_22790_41880# SUNSAR_CAPT8B_CV_0.XA4.Y 0.111538f
C1432 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.301485f
C1433 SUNSAR_SAR8B_CV_0.DONE SUNSAR_SAR8B_CV_0.XA7.CEO 0.301665f
C1434 a_3782_41352# VPWR 0.394053f
C1435 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.327909f
C1436 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C1437 a_23922_34540# VPWR 0.502044f
C1438 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.D VPWR 0.104609f
C1439 SUNSAR_CAPT8B_CV_0.XH13.QN VPWR 0.901622f
C1440 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.649845f
C1441 SUNSAR_SAR8B_CV_0.XB1.XA1.Y SUNSAR_SAR8B_CV_0.XB1.M3.G 0.224309f
C1442 a_8822_42408# VPWR 0.391292f
C1443 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.419738f
C1444 SUNSAR_SAR8B_CV_0.XB2.M3.G VPWR 0.665006f
C1445 a_18902_40648# VPWR 0.491225f
C1446 SUNSAR_CAPT8B_CV_0.XA3.Y SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y 0.254583f
C1447 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.D VPWR 0.104609f
C1448 uo_out[0] uo_out[1] 0.366897f
C1449 SUNSAR_SAR8B_CV_0.XA2.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C1450 a_20250_27148# VPWR 0.470364f
C1451 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP0.D VPWR 0.106927f
C1452 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA4.XA11.Y 0.220689f
C1453 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.240612f
C1454 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.86675f
C1455 SUNSAR_CAPT8B_CV_0.XB07.QN uo_out[7] 0.263255f
C1456 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C1457 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VPWR 1.77562f
C1458 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.255261f
C1459 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON 0.702226f
C1460 SUNSAR_SAR8B_CV_0.XA6.ENO a_17730_28556# 0.132757f
C1461 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S 0.363295f
C1462 a_13862_42760# SUNSAR_CAPT8B_CV_0.XF11.XA4.A 0.113305f
C1463 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VPWR 0.714341f
C1464 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1465 SUNSAR_CAPT8B_CV_0.XG12.QN VPWR 0.901622f
C1466 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y SUNSAR_CAPT8B_CV_0.XC08.XA4.A 0.744161f
C1467 a_16542_4566# VPWR 0.413433f
C1468 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6519f
C1469 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VPWR 0.271482f
C1470 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.820808f
C1471 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.59087f
C1472 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.29297f
C1473 a_10190_43816# VPWR 0.391817f
C1474 a_18882_27148# VPWR 0.471462f
C1475 SUNSAR_SAR8B_CV_0.XA0.CMP_OP SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y 0.383512f
C1476 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C1477 a_10170_32076# VPWR 0.436368f
C1478 SUNSAR_SAR8B_CV_0.XA20.XA1.CK SUNSAR_SAR8B_CV_0.XA20.XA2.VMR 0.380687f
C1479 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VPWR 2.95303f
C1480 a_10170_28204# VPWR 0.361706f
C1481 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.267238f
C1482 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y 0.204048f
C1483 SUNSAR_CAPT8B_CV_0.XA4.MN0.S VPWR 0.635621f
C1484 SUNSAR_SAR8B_CV_0.XA7.CEO VPWR 1.1111f
C1485 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VPWR 1.77562f
C1486 SUNSAR_SAR8B_CV_0.XA1.ENO SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.164325f
C1487 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[6] 0.258218f
C1488 SUNSAR_CAPT8B_CV_0.XF11.QN VPWR 0.901622f
C1489 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 0.440586f
C1490 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.419738f
C1491 SUNSAR_SAR8B_CV_0.XA0.XA10.Y a_2610_36300# 0.13253f
C1492 a_10170_35068# VPWR 0.394528f
C1493 SUNSAR_SAR8B_CV_0.XA0.ENO SUNSAR_SAR8B_CV_0.XA0.CMP_OP 0.6934f
C1494 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.2622f
C1495 a_8822_43816# VPWR 0.391817f
C1496 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87301f
C1497 SUNSAR_SAR8B_CV_0.XA3.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.377598f
C1498 a_10170_35948# VPWR 0.417826f
C1499 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 13.6523f
C1500 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_6282_35420# 0.160931f
C1501 a_8802_32076# VPWR 0.436368f
C1502 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1503 a_8802_28204# VPWR 0.36179f
C1504 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON 0.702226f
C1505 SUNSAR_SAR8B_CV_0.XA5.ENO a_16362_28556# 0.135353f
C1506 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D 0.109021f
C1507 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VPWR 0.723713f
C1508 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VPWR 2.95308f
C1509 SUNSAR_CAPT8B_CV_0.XE10.QN VPWR 0.901622f
C1510 SUNSAR_SAR8B_CV_0.XB1.M3.G VPWR 0.665006f
C1511 a_15230_40648# VPWR 0.492579f
C1512 a_8802_35068# VPWR 0.394528f
C1513 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.88588f
C1514 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C1515 a_18902_41352# VPWR 0.394053f
C1516 a_8802_35948# VPWR 0.417826f
C1517 SUNSAR_SAR8B_CV_0.XA1.XA8.A a_5130_35420# 0.133834f
C1518 SUNSAR_SAR8B_CV_0.XA20.XA10.B SUNSAR_SAR8B_CV_0.XA20.XA1.CKN 0.126085f
C1519 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C1520 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP0.D VPWR 0.106927f
C1521 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.327152f
C1522 SUNSAR_SAR8B_CV_0.XA6.CEO VPWR 2.28789f
C1523 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C1524 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y SUNSAR_SAR8B_CV_0.DONE 0.227625f
C1525 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GNG 1.62434f
C1526 SUNSAR_CAPT8B_CV_0.XD09.QN VPWR 0.901622f
C1527 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y SUNSAR_CAPT8B_CV_0.XH13.XA4.A 0.744161f
C1528 SUNSAR_SAR8B_CV_0.XB2.XA3.B m3_24750_2768# 0.172147f
C1529 a_13862_40648# VPWR 0.491225f
C1530 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38576f
C1531 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C1532 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.D VPWR 0.104609f
C1533 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.431984f
C1534 a_15210_27148# VPWR 0.470364f
C1535 SUNSAR_SAR8B_CV_0.XA2.CEO SUNSAR_SAR8B_CV_0.XA3.XA11.Y 0.293159f
C1536 SUNSAR_SAR8B_CV_0.XA5.XA6.Y SUNSAR_SAR8B_CV_0.XA5.XA8.A 0.527529f
C1537 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y a_18902_41000# 0.15757f
C1538 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1615f
C1539 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP 0.11382f
C1540 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VPWR 2.95304f
C1541 TIE_L uo_out[1] 0.50141f
C1542 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON 0.702226f
C1543 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y 0.37807f
C1544 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VPWR 0.720096f
C1545 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR 0.112098f
C1546 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y ui_in[0] 0.172623f
C1547 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP0.D VPWR 0.106927f
C1548 SUNSAR_CAPT8B_CV_0.XC08.QN VPWR 0.901622f
C1549 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.D VPWR 0.104609f
C1550 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.B 0.146458f
C1551 ua[2] VGND 0.117454f
C1552 ua[3] VGND 0.117454f
C1553 ua[4] VGND 0.118698f
C1554 ua[5] VGND 0.120088f
C1555 ua[6] VGND 0.120088f
C1556 ua[7] VGND 0.111009f
C1557 ua[0] VGND 7.62793f
C1558 ua[1] VGND 6.98581f
C1559 ui_in[0] VGND 5.66164f
C1560 clk VGND 6.42293f
C1561 uo_out[0] VGND 2.81872f
C1562 uo_out[1] VGND 1.77173f
C1563 uo_out[2] VGND 1.57211f
C1564 uo_out[3] VGND 1.79184f
C1565 uo_out[4] VGND 1.64454f
C1566 uo_out[5] VGND 2.45226f
C1567 uo_out[6] VGND 2.74323f
C1568 uo_out[7] VGND 3.47431f
C1569 VPWR VGND 0.941568p
C1570 TIE_L1 VGND 1.5148f
C1571 TIE_L2 VGND 1.73849f
C1572 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93609f
C1573 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93609f
C1574 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.5533f
C1575 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.5533f
C1576 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.334839f
C1577 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.334839f
C1578 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.469f
C1579 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.469f
C1580 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43533f
C1581 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43533f
C1582 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67745f
C1583 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67745f
C1584 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.6684f
C1585 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.6684f
C1586 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.574499f
C1587 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.574499f
C1588 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33412f
C1589 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33412f
C1590 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.469f
C1591 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.469f
C1592 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43533f
C1593 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43533f
C1594 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67745f
C1595 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67745f
C1596 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.6684f
C1597 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.6684f
C1598 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.575099f
C1599 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.575099f
C1600 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33412f
C1601 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33412f
C1602 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.469f
C1603 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.469f
C1604 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43533f
C1605 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43533f
C1606 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67745f
C1607 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67745f
C1608 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.6684f
C1609 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.6684f
C1610 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.571799f
C1611 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.571799f
C1612 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33412f
C1613 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33412f
C1614 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.471901f
C1615 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.471901f
C1616 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.439809f
C1617 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44253f
C1618 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.3859f
C1619 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.38266f
C1620 a_15390_2630# VGND 0.542161f $ **FLOATING
C1621 a_13950_2630# VGND 0.427094f $ **FLOATING
C1622 a_12582_2630# VGND 0.426679f $ **FLOATING
C1623 a_11142_2630# VGND 0.543317f $ **FLOATING
C1624 a_15390_2982# VGND 0.491607f $ **FLOATING
C1625 a_13950_2982# VGND 0.352472f $ **FLOATING
C1626 a_12582_2982# VGND 0.352472f $ **FLOATING
C1627 a_11142_2982# VGND 0.490037f $ **FLOATING
C1628 a_15390_3334# VGND 0.374919f $ **FLOATING
C1629 a_13950_3334# VGND 0.352438f $ **FLOATING
C1630 a_12582_3334# VGND 0.352438f $ **FLOATING
C1631 a_11142_3334# VGND 0.374919f $ **FLOATING
C1632 a_13950_3686# VGND 0.352418f $ **FLOATING
C1633 a_12582_3686# VGND 0.352418f $ **FLOATING
C1634 SUNSAR_SAR8B_CV_0.XB2.XA3.B VGND 41.5268f
C1635 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.70146f
C1636 SUNSAR_SAR8B_CV_0.XB1.XA3.B VGND 41.5268f
C1637 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.70146f
C1638 a_15390_4038# VGND 0.397033f $ **FLOATING
C1639 a_13950_4038# VGND 0.354407f $ **FLOATING
C1640 a_12582_4038# VGND 0.354407f $ **FLOATING
C1641 a_11142_4038# VGND 0.397033f $ **FLOATING
C1642 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG VGND 37.7832f
C1643 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.38998f
C1644 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.D VGND 0.103625f
C1645 a_13950_4390# VGND 0.352432f $ **FLOATING
C1646 a_12582_4390# VGND 0.352432f $ **FLOATING
C1647 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.D VGND 0.103625f
C1648 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.38998f
C1649 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG VGND 37.7832f
C1650 SUNSAR_SAR8B_CV_0.XB2.M3.G VGND 3.1165f
C1651 a_15390_4566# VGND 0.389036f $ **FLOATING
C1652 SUNSAR_SAR8B_CV_0.XB1.M3.G VGND 3.07938f
C1653 a_11142_4566# VGND 0.389036f $ **FLOATING
C1654 SUNSAR_SAR8B_CV_0.XB2.XA1.Y VGND 0.970036f
C1655 a_13950_4742# VGND 0.352456f $ **FLOATING
C1656 a_12582_4742# VGND 0.352456f $ **FLOATING
C1657 SUNSAR_SAR8B_CV_0.XB2.XA1.MN0.G VGND 0.7964f
C1658 a_15390_4918# VGND 0.470144f $ **FLOATING
C1659 SUNSAR_SAR8B_CV_0.XB1.XA1.MN0.G VGND 0.7964f
C1660 SUNSAR_SAR8B_CV_0.XB1.XA1.Y VGND 0.970036f
C1661 a_11142_4918# VGND 0.471715f $ **FLOATING
C1662 a_13950_5094# VGND 0.353103f $ **FLOATING
C1663 a_12582_5094# VGND 0.353103f $ **FLOATING
C1664 a_15390_5270# VGND 0.492927f $ **FLOATING
C1665 a_11142_5270# VGND 0.491356f $ **FLOATING
C1666 SUNSAR_SAR8B_CV_0.XB2.XA2.MN0.G VGND 0.596866f
C1667 a_13950_5446# VGND 0.433341f $ **FLOATING
C1668 a_12582_5446# VGND 0.433756f $ **FLOATING
C1669 a_15390_5622# VGND 0.47219f $ **FLOATING
C1670 a_15390_5974# VGND 0.541341f $ **FLOATING
C1671 SUNSAR_SAR8B_CV_0.XB1.XA2.MN0.G VGND 0.596866f
C1672 a_11142_5622# VGND 0.47376f $ **FLOATING
C1673 a_11142_5974# VGND 0.540186f $ **FLOATING
C1674 a_22770_26796# VGND 0.529341f $ **FLOATING
C1675 a_21402_26796# VGND 0.531659f $ **FLOATING
C1676 a_17730_26796# VGND 0.530834f $ **FLOATING
C1677 a_16362_26796# VGND 0.531989f $ **FLOATING
C1678 a_12690_26796# VGND 0.530834f $ **FLOATING
C1679 a_11322_26796# VGND 0.531989f $ **FLOATING
C1680 a_7650_26796# VGND 0.530213f $ **FLOATING
C1681 a_6282_26796# VGND 0.530979f $ **FLOATING
C1682 a_2610_26796# VGND 0.531178f $ **FLOATING
C1683 a_22770_27148# VGND 0.499848f $ **FLOATING
C1684 a_21402_27148# VGND 0.467094f $ **FLOATING
C1685 a_17730_27148# VGND 0.471508f $ **FLOATING
C1686 a_16362_27148# VGND 0.467722f $ **FLOATING
C1687 a_12690_27148# VGND 0.471508f $ **FLOATING
C1688 a_11322_27148# VGND 0.467722f $ **FLOATING
C1689 a_7650_27148# VGND 0.470266f $ **FLOATING
C1690 a_6282_27148# VGND 0.465734f $ **FLOATING
C1691 a_2610_27148# VGND 0.47123f $ **FLOATING
C1692 a_21402_27500# VGND 0.385968f $ **FLOATING
C1693 a_17730_27500# VGND 0.387712f $ **FLOATING
C1694 a_16362_27500# VGND 0.386249f $ **FLOATING
C1695 a_12690_27500# VGND 0.387712f $ **FLOATING
C1696 a_11322_27500# VGND 0.386249f $ **FLOATING
C1697 a_7650_27500# VGND 0.38671f $ **FLOATING
C1698 a_6282_27500# VGND 0.384229f $ **FLOATING
C1699 a_2610_27500# VGND 0.387675f $ **FLOATING
C1700 a_21402_27852# VGND 0.370125f $ **FLOATING
C1701 a_17730_27852# VGND 0.370785f $ **FLOATING
C1702 a_16362_27852# VGND 0.368771f $ **FLOATING
C1703 a_12690_27852# VGND 0.370785f $ **FLOATING
C1704 a_11322_27852# VGND 0.368771f $ **FLOATING
C1705 a_7650_27852# VGND 0.369543f $ **FLOATING
C1706 a_6282_27852# VGND 0.366751f $ **FLOATING
C1707 a_2610_27852# VGND 0.370508f $ **FLOATING
C1708 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.D VGND 0.506947f
C1709 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.D VGND 0.502211f
C1710 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.D VGND 0.477244f
C1711 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.D VGND 0.502211f
C1712 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.D VGND 0.477244f
C1713 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.D VGND 0.502211f
C1714 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.D VGND 0.477244f
C1715 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.D VGND 0.502211f
C1716 a_21402_28204# VGND 0.405715f $ **FLOATING
C1717 a_17730_28204# VGND 0.406284f $ **FLOATING
C1718 a_16362_28204# VGND 0.406284f $ **FLOATING
C1719 a_12690_28204# VGND 0.406284f $ **FLOATING
C1720 a_11322_28204# VGND 0.406284f $ **FLOATING
C1721 a_7650_28204# VGND 0.405133f $ **FLOATING
C1722 a_6282_28204# VGND 0.404355f $ **FLOATING
C1723 a_2610_28204# VGND 0.406098f $ **FLOATING
C1724 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.D VGND 0.608956f
C1725 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.S VGND 0.741242f
C1726 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.S VGND 0.749251f
C1727 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.S VGND 0.735502f
C1728 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.S VGND 0.749251f
C1729 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.S VGND 0.735502f
C1730 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.S VGND 0.746591f
C1731 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.S VGND 0.73057f
C1732 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.S VGND 0.74895f
C1733 a_22770_28556# VGND 0.401649f $ **FLOATING
C1734 a_21402_28556# VGND 0.387558f $ **FLOATING
C1735 a_17730_28556# VGND 0.388127f $ **FLOATING
C1736 a_16362_28556# VGND 0.388127f $ **FLOATING
C1737 a_12690_28556# VGND 0.388127f $ **FLOATING
C1738 a_11322_28556# VGND 0.388127f $ **FLOATING
C1739 a_7650_28556# VGND 0.386976f $ **FLOATING
C1740 a_6282_28556# VGND 0.386198f $ **FLOATING
C1741 a_2610_28556# VGND 0.38794f $ **FLOATING
C1742 a_21402_28908# VGND 0.394283f $ **FLOATING
C1743 a_17730_28908# VGND 0.394852f $ **FLOATING
C1744 a_16362_28908# VGND 0.394852f $ **FLOATING
C1745 a_12690_28908# VGND 0.394852f $ **FLOATING
C1746 a_11322_28908# VGND 0.394852f $ **FLOATING
C1747 a_7650_28908# VGND 0.393701f $ **FLOATING
C1748 a_6282_28908# VGND 0.392923f $ **FLOATING
C1749 a_2610_28908# VGND 0.394666f $ **FLOATING
C1750 SUNSAR_SAR8B_CV_0.SARP VGND 70.097496f
C1751 a_21402_29612# VGND 0.395457f $ **FLOATING
C1752 a_17730_29612# VGND 0.396116f $ **FLOATING
C1753 a_16362_29612# VGND 0.395588f $ **FLOATING
C1754 a_12690_29612# VGND 0.396116f $ **FLOATING
C1755 a_11322_29612# VGND 0.395588f $ **FLOATING
C1756 a_7650_29612# VGND 0.394965f $ **FLOATING
C1757 a_6282_29612# VGND 0.393746f $ **FLOATING
C1758 a_2610_29612# VGND 0.395923f $ **FLOATING
C1759 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318647f
C1760 a_22770_29964# VGND 0.400512f $ **FLOATING
C1761 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.D VGND 0.103281f
C1762 SUNSAR_SAR8B_CV_0.XA7.XA1.XA2.Y VGND 1.27143f
C1763 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.D VGND 0.100021f
C1764 SUNSAR_SAR8B_CV_0.XA6.XA1.XA2.Y VGND 1.26503f
C1765 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.D VGND 0.100021f
C1766 SUNSAR_SAR8B_CV_0.XA5.XA1.XA2.Y VGND 1.26391f
C1767 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.D VGND 0.100021f
C1768 SUNSAR_SAR8B_CV_0.XA4.XA1.XA2.Y VGND 1.26503f
C1769 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.D VGND 0.100021f
C1770 SUNSAR_SAR8B_CV_0.XA3.XA1.XA2.Y VGND 1.26391f
C1771 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.D VGND 0.100021f
C1772 SUNSAR_SAR8B_CV_0.XA2.XA1.XA2.Y VGND 1.25938f
C1773 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.D VGND 0.100021f
C1774 SUNSAR_SAR8B_CV_0.XA1.XA1.XA2.Y VGND 1.25329f
C1775 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.D VGND 0.100021f
C1776 SUNSAR_SAR8B_CV_0.XA0.XA1.XA2.Y VGND 1.26407f
C1777 a_21402_30316# VGND 0.401758f $ **FLOATING
C1778 a_17730_30316# VGND 0.401074f $ **FLOATING
C1779 a_16362_30316# VGND 0.401074f $ **FLOATING
C1780 a_12690_30316# VGND 0.401074f $ **FLOATING
C1781 a_11322_30316# VGND 0.401074f $ **FLOATING
C1782 a_7650_30316# VGND 0.399923f $ **FLOATING
C1783 a_6282_30316# VGND 0.399145f $ **FLOATING
C1784 a_2610_30316# VGND 0.400881f $ **FLOATING
C1785 SUNSAR_SAR8B_CV_0.XA0.CMP_OP VGND 15.315499f
C1786 a_22770_30844# VGND 0.421853f $ **FLOATING
C1787 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON VGND 2.24318f
C1788 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON VGND 2.22194f
C1789 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON VGND 2.22198f
C1790 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON VGND 2.22194f
C1791 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON VGND 2.22198f
C1792 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON VGND 2.20909f
C1793 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON VGND 2.19751f
C1794 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON VGND 2.21827f
C1795 a_21402_31196# VGND 0.4255f $ **FLOATING
C1796 a_17730_31196# VGND 0.426069f $ **FLOATING
C1797 a_16362_31196# VGND 0.426069f $ **FLOATING
C1798 a_12690_31196# VGND 0.426069f $ **FLOATING
C1799 a_11322_31196# VGND 0.426069f $ **FLOATING
C1800 a_7650_31196# VGND 0.424917f $ **FLOATING
C1801 a_6282_31196# VGND 0.42414f $ **FLOATING
C1802 a_2610_31196# VGND 0.425876f $ **FLOATING
C1803 SUNSAR_SAR8B_CV_0.XA0.CMP_ON VGND 19.4783f
C1804 a_22770_31724# VGND 0.423601f $ **FLOATING
C1805 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.99939f
C1806 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.97987f
C1807 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.97901f
C1808 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.97987f
C1809 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.97901f
C1810 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.85828f
C1811 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.37577f
C1812 a_21402_32076# VGND 0.426091f $ **FLOATING
C1813 a_17730_32076# VGND 0.42666f $ **FLOATING
C1814 a_16362_32076# VGND 0.42666f $ **FLOATING
C1815 a_12690_32076# VGND 0.42666f $ **FLOATING
C1816 a_11322_32076# VGND 0.42666f $ **FLOATING
C1817 a_7650_32076# VGND 0.42666f $ **FLOATING
C1818 a_6282_32076# VGND 0.42666f $ **FLOATING
C1819 a_2610_32076# VGND 0.426468f $ **FLOATING
C1820 SUNSAR_SAR8B_CV_0.XA20.XA2.N1 VGND 1.55564f
C1821 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C1822 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP VGND 3.19736f
C1823 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP VGND 3.22974f
C1824 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP VGND 3.22835f
C1825 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP VGND 3.22974f
C1826 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP VGND 3.22835f
C1827 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP VGND 3.22678f
C1828 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP VGND 3.22545f
C1829 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP VGND 3.31413f
C1830 SUNSAR_SAR8B_CV_0.XA20.XA2.CO VGND 2.68549f
C1831 a_21402_32956# VGND 0.426069f $ **FLOATING
C1832 a_17730_32956# VGND 0.426069f $ **FLOATING
C1833 a_16362_32956# VGND 0.426069f $ **FLOATING
C1834 a_12690_32956# VGND 0.426069f $ **FLOATING
C1835 a_11322_32956# VGND 0.426069f $ **FLOATING
C1836 a_7650_32956# VGND 0.426069f $ **FLOATING
C1837 a_6282_32956# VGND 0.426069f $ **FLOATING
C1838 a_2610_32956# VGND 0.425876f $ **FLOATING
C1839 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR VGND 2.85099f
C1840 a_22770_33132# VGND 0.403395f $ **FLOATING
C1841 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 3.01164f
C1842 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.01628f
C1843 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.01641f
C1844 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.01628f
C1845 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.01641f
C1846 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.54669f
C1847 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.78758f
C1848 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 12.1041f
C1849 a_21402_33836# VGND 0.426756f $ **FLOATING
C1850 a_17730_33836# VGND 0.426756f $ **FLOATING
C1851 a_16362_33836# VGND 0.426756f $ **FLOATING
C1852 a_12690_33836# VGND 0.426756f $ **FLOATING
C1853 a_11322_33836# VGND 0.426756f $ **FLOATING
C1854 a_7650_33836# VGND 0.426756f $ **FLOATING
C1855 a_6282_33836# VGND 0.426756f $ **FLOATING
C1856 a_2610_33836# VGND 0.426472f $ **FLOATING
C1857 SUNSAR_SAR8B_CV_0.SARN VGND 71.1589f
C1858 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND 0.149691f
C1859 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.D VGND 0.515385f
C1860 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C1861 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND 0.149691f
C1862 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.72791f
C1863 a_22770_34540# VGND 0.39377f $ **FLOATING
C1864 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND 0.102f
C1865 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND 0.149691f
C1866 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 4.1719f
C1867 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND 0.149691f
C1868 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.27991f
C1869 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND 0.102f
C1870 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND 0.102f
C1871 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND 0.149691f
C1872 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.31299f
C1873 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND 0.149691f
C1874 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.68294f
C1875 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND 0.102f
C1876 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND 0.102f
C1877 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND 0.149691f
C1878 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 4.25175f
C1879 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND 0.149691f
C1880 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 10.150401f
C1881 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND 0.102f
C1882 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND 0.102f
C1883 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND 0.102f
C1884 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 8.127279f
C1885 a_21402_34716# VGND 0.39476f $ **FLOATING
C1886 a_17730_34716# VGND 0.39476f $ **FLOATING
C1887 a_16362_34716# VGND 0.39476f $ **FLOATING
C1888 a_12690_34716# VGND 0.39476f $ **FLOATING
C1889 a_11322_34716# VGND 0.39476f $ **FLOATING
C1890 a_7650_34716# VGND 0.39476f $ **FLOATING
C1891 a_6282_34716# VGND 0.39476f $ **FLOATING
C1892 a_2610_34716# VGND 0.394567f $ **FLOATING
C1893 SUNSAR_SAR8B_CV_0.XA20.XA1.CK VGND 4.75219f
C1894 a_22770_34892# VGND 0.394644f $ **FLOATING
C1895 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.67603f
C1896 SUNSAR_SAR8B_CV_0.XA6.ENO VGND 4.51439f
C1897 SUNSAR_SAR8B_CV_0.XA5.ENO VGND 4.46191f
C1898 SUNSAR_SAR8B_CV_0.XA4.ENO VGND 4.27708f
C1899 SUNSAR_SAR8B_CV_0.XA3.ENO VGND 4.50282f
C1900 SUNSAR_SAR8B_CV_0.XA2.ENO VGND 4.42572f
C1901 SUNSAR_SAR8B_CV_0.XA1.ENO VGND 4.44437f
C1902 SUNSAR_SAR8B_CV_0.XA0.ENO VGND 4.39222f
C1903 a_21402_35068# VGND 0.389563f $ **FLOATING
C1904 a_17730_35068# VGND 0.389563f $ **FLOATING
C1905 a_16362_35068# VGND 0.389563f $ **FLOATING
C1906 a_12690_35068# VGND 0.389563f $ **FLOATING
C1907 a_11322_35068# VGND 0.389563f $ **FLOATING
C1908 a_7650_35068# VGND 0.389563f $ **FLOATING
C1909 a_6282_35068# VGND 0.389563f $ **FLOATING
C1910 a_2610_35068# VGND 0.38937f $ **FLOATING
C1911 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN VGND 4.54316f
C1912 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C1913 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C1914 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C1915 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C1916 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C1917 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C1918 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557214f
C1919 a_22770_35420# VGND 0.395535f $ **FLOATING
C1920 a_21402_35420# VGND 0.389041f $ **FLOATING
C1921 a_17730_35420# VGND 0.388925f $ **FLOATING
C1922 a_16362_35420# VGND 0.389297f $ **FLOATING
C1923 a_12690_35420# VGND 0.388925f $ **FLOATING
C1924 a_11322_35420# VGND 0.389297f $ **FLOATING
C1925 a_7650_35420# VGND 0.388925f $ **FLOATING
C1926 a_6282_35420# VGND 0.389297f $ **FLOATING
C1927 a_2610_35420# VGND 0.389015f $ **FLOATING
C1928 SUNSAR_SAR8B_CV_0.XA20.XA10.A VGND 1.07685f
C1929 SUNSAR_SAR8B_CV_0.XA7.XA9.MN0.D VGND 0.112889f
C1930 SUNSAR_SAR8B_CV_0.XA7.XA8.A VGND 1.50901f
C1931 SUNSAR_SAR8B_CV_0.XA7.XA6.Y VGND 1.53168f
C1932 SUNSAR_SAR8B_CV_0.XA6.XA8.A VGND 1.50964f
C1933 SUNSAR_SAR8B_CV_0.XA6.XA9.MN0.D VGND 0.112889f
C1934 SUNSAR_SAR8B_CV_0.XA6.XA6.Y VGND 1.54335f
C1935 SUNSAR_SAR8B_CV_0.XA5.XA9.MN0.D VGND 0.112889f
C1936 SUNSAR_SAR8B_CV_0.XA5.XA8.A VGND 1.51005f
C1937 SUNSAR_SAR8B_CV_0.XA5.XA6.Y VGND 1.53305f
C1938 SUNSAR_SAR8B_CV_0.XA4.XA8.A VGND 1.50964f
C1939 SUNSAR_SAR8B_CV_0.XA4.XA9.MN0.D VGND 0.112889f
C1940 SUNSAR_SAR8B_CV_0.XA4.XA6.Y VGND 1.54335f
C1941 SUNSAR_SAR8B_CV_0.XA3.XA9.MN0.D VGND 0.112889f
C1942 SUNSAR_SAR8B_CV_0.XA3.XA8.A VGND 1.51005f
C1943 SUNSAR_SAR8B_CV_0.XA3.XA6.Y VGND 1.53305f
C1944 SUNSAR_SAR8B_CV_0.XA2.XA8.A VGND 1.50964f
C1945 SUNSAR_SAR8B_CV_0.XA2.XA9.MN0.D VGND 0.112889f
C1946 SUNSAR_SAR8B_CV_0.XA2.XA6.Y VGND 1.54335f
C1947 SUNSAR_SAR8B_CV_0.XA1.XA9.MN0.D VGND 0.112889f
C1948 SUNSAR_SAR8B_CV_0.XA1.XA8.A VGND 1.51005f
C1949 SUNSAR_SAR8B_CV_0.XA1.XA6.Y VGND 1.53305f
C1950 SUNSAR_SAR8B_CV_0.XA0.XA8.A VGND 1.51935f
C1951 SUNSAR_SAR8B_CV_0.XA0.XA9.MN0.D VGND 0.112889f
C1952 SUNSAR_SAR8B_CV_0.XA0.XA6.Y VGND 1.61753f
C1953 a_22770_35948# VGND 0.414038f $ **FLOATING
C1954 a_21402_35948# VGND 0.390722f $ **FLOATING
C1955 a_17730_35948# VGND 0.391291f $ **FLOATING
C1956 a_16362_35948# VGND 0.391291f $ **FLOATING
C1957 a_12690_35948# VGND 0.391291f $ **FLOATING
C1958 a_11322_35948# VGND 0.391291f $ **FLOATING
C1959 a_7650_35948# VGND 0.391291f $ **FLOATING
C1960 a_6282_35948# VGND 0.391291f $ **FLOATING
C1961 a_2610_35948# VGND 0.391099f $ **FLOATING
C1962 SUNSAR_SAR8B_CV_0.XA20.XA10.B VGND 0.789814f
C1963 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C1964 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C1965 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C1966 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C1967 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C1968 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C1969 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C1970 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.895311f
C1971 a_22770_36300# VGND 0.472701f $ **FLOATING
C1972 a_21402_36300# VGND 0.393831f $ **FLOATING
C1973 a_17730_36300# VGND 0.394738f $ **FLOATING
C1974 a_16362_36300# VGND 0.3944f $ **FLOATING
C1975 a_12690_36300# VGND 0.394718f $ **FLOATING
C1976 a_11322_36300# VGND 0.3944f $ **FLOATING
C1977 a_7650_36300# VGND 0.394715f $ **FLOATING
C1978 a_6282_36300# VGND 0.3944f $ **FLOATING
C1979 a_2610_36300# VGND 0.394523f $ **FLOATING
C1980 a_22770_36652# VGND 0.542245f $ **FLOATING
C1981 SUNSAR_SAR8B_CV_0.XA7.XA10.Y VGND 0.881626f
C1982 SUNSAR_SAR8B_CV_0.XA6.XA10.Y VGND 0.884627f
C1983 SUNSAR_SAR8B_CV_0.XA5.XA10.Y VGND 0.877071f
C1984 SUNSAR_SAR8B_CV_0.XA4.XA10.Y VGND 0.884604f
C1985 SUNSAR_SAR8B_CV_0.XA3.XA10.Y VGND 0.877059f
C1986 SUNSAR_SAR8B_CV_0.XA2.XA10.Y VGND 0.884603f
C1987 SUNSAR_SAR8B_CV_0.XA1.XA10.Y VGND 0.877071f
C1988 SUNSAR_SAR8B_CV_0.XA0.XA10.Y VGND 0.892649f
C1989 SUNSAR_SAR8B_CV_0.XB1.TIE_L VGND 32.9183f
C1990 a_21402_36828# VGND 0.414041f $ **FLOATING
C1991 a_17730_36828# VGND 0.413952f $ **FLOATING
C1992 a_16362_36828# VGND 0.413659f $ **FLOATING
C1993 a_12690_36828# VGND 0.413942f $ **FLOATING
C1994 a_11322_36828# VGND 0.413658f $ **FLOATING
C1995 a_7650_36828# VGND 0.413944f $ **FLOATING
C1996 a_6282_36828# VGND 0.413659f $ **FLOATING
C1997 a_2610_36828# VGND 0.413594f $ **FLOATING
C1998 SUNSAR_SAR8B_CV_0.XA7.XA11.Y VGND 1.08552f
C1999 SUNSAR_SAR8B_CV_0.XA7.CEO VGND 2.06017f
C2000 SUNSAR_SAR8B_CV_0.XA6.XA11.Y VGND 1.10839f
C2001 SUNSAR_SAR8B_CV_0.XA6.CEO VGND 1.45333f
C2002 SUNSAR_SAR8B_CV_0.XA5.XA11.Y VGND 1.06778f
C2003 SUNSAR_SAR8B_CV_0.XA5.CEO VGND 1.71757f
C2004 SUNSAR_SAR8B_CV_0.XA4.XA11.Y VGND 1.10834f
C2005 SUNSAR_SAR8B_CV_0.XA4.CEO VGND 1.52588f
C2006 SUNSAR_SAR8B_CV_0.XA3.XA11.Y VGND 1.06777f
C2007 SUNSAR_SAR8B_CV_0.XA3.CEO VGND 1.71756f
C2008 SUNSAR_SAR8B_CV_0.XA2.XA11.Y VGND 1.10835f
C2009 SUNSAR_SAR8B_CV_0.XA2.CEO VGND 1.52589f
C2010 SUNSAR_SAR8B_CV_0.XA1.XA11.Y VGND 1.06778f
C2011 SUNSAR_SAR8B_CV_0.XA1.CEO VGND 1.71756f
C2012 SUNSAR_SAR8B_CV_0.XA0.XA11.Y VGND 1.11927f
C2013 SUNSAR_SAR8B_CV_0.XA0.CEO VGND 1.53308f
C2014 a_21402_37180# VGND 0.47501f $ **FLOATING
C2015 a_17730_37180# VGND 0.474809f $ **FLOATING
C2016 a_16362_37180# VGND 0.476355f $ **FLOATING
C2017 a_12690_37180# VGND 0.47479f $ **FLOATING
C2018 a_11322_37180# VGND 0.476354f $ **FLOATING
C2019 a_7650_37180# VGND 0.474794f $ **FLOATING
C2020 a_6282_37180# VGND 0.476355f $ **FLOATING
C2021 a_2610_37180# VGND 0.474277f $ **FLOATING
C2022 a_21402_37532# VGND 0.546649f $ **FLOATING
C2023 a_17730_37532# VGND 0.548986f $ **FLOATING
C2024 a_16362_37532# VGND 0.547631f $ **FLOATING
C2025 a_12690_37532# VGND 0.548815f $ **FLOATING
C2026 a_11322_37532# VGND 0.547631f $ **FLOATING
C2027 a_7650_37532# VGND 0.548857f $ **FLOATING
C2028 a_6282_37532# VGND 0.547634f $ **FLOATING
C2029 a_2610_37532# VGND 0.546853f $ **FLOATING
C2030 a_22790_40296# VGND 0.546732f $ **FLOATING
C2031 a_21422_40296# VGND 0.54563f $ **FLOATING
C2032 a_17750_40296# VGND 0.546813f $ **FLOATING
C2033 a_16382_40296# VGND 0.547966f $ **FLOATING
C2034 a_12710_40296# VGND 0.546813f $ **FLOATING
C2035 a_11342_40296# VGND 0.547969f $ **FLOATING
C2036 a_7670_40296# VGND 0.54681f $ **FLOATING
C2037 a_6302_40296# VGND 0.547966f $ **FLOATING
C2038 a_2630_40296# VGND 0.54539f $ **FLOATING
C2039 a_22790_40648# VGND 0.492438f $ **FLOATING
C2040 a_21422_40648# VGND 0.49034f $ **FLOATING
C2041 a_17750_40648# VGND 0.492453f $ **FLOATING
C2042 a_16382_40648# VGND 0.490883f $ **FLOATING
C2043 a_12710_40648# VGND 0.492453f $ **FLOATING
C2044 a_11342_40648# VGND 0.490883f $ **FLOATING
C2045 a_7670_40648# VGND 0.492453f $ **FLOATING
C2046 a_6302_40648# VGND 0.490883f $ **FLOATING
C2047 a_2630_40648# VGND 0.492826f $ **FLOATING
C2048 SUNSAR_SAR8B_CV_0.DONE VGND 20.737402f
C2049 a_22790_41000# VGND 0.388777f $ **FLOATING
C2050 a_21422_41000# VGND 0.388174f $ **FLOATING
C2051 a_17750_41000# VGND 0.388174f $ **FLOATING
C2052 a_16382_41000# VGND 0.388174f $ **FLOATING
C2053 a_12710_41000# VGND 0.388174f $ **FLOATING
C2054 a_11342_41000# VGND 0.388174f $ **FLOATING
C2055 a_7670_41000# VGND 0.388174f $ **FLOATING
C2056 a_6302_41000# VGND 0.388174f $ **FLOATING
C2057 a_2630_41000# VGND 0.388638f $ **FLOATING
C2058 a_22790_41352# VGND 0.374594f $ **FLOATING
C2059 a_21422_41352# VGND 0.393558f $ **FLOATING
C2060 a_17750_41352# VGND 0.393558f $ **FLOATING
C2061 a_16382_41352# VGND 0.393558f $ **FLOATING
C2062 a_12710_41352# VGND 0.393558f $ **FLOATING
C2063 a_11342_41352# VGND 0.393558f $ **FLOATING
C2064 a_7670_41352# VGND 0.393558f $ **FLOATING
C2065 a_6302_41352# VGND 0.393558f $ **FLOATING
C2066 a_2630_41352# VGND 0.394022f $ **FLOATING
C2067 SUNSAR_CAPT8B_CV_0.XA4.MN0.S VGND 0.803097f
C2068 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.D VGND 0.107737f
C2069 SUNSAR_SAR8B_CV_0.D<0> VGND 5.87227f
C2070 SUNSAR_SAR8B_CV_0.D<1> VGND 13.789701f
C2071 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN0.D VGND 0.107643f
C2072 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN0.D VGND 0.107643f
C2073 SUNSAR_SAR8B_CV_0.D<2> VGND 12.5832f
C2074 SUNSAR_SAR8B_CV_0.D<3> VGND 11.4395f
C2075 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN0.D VGND 0.107643f
C2076 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN0.D VGND 0.107643f
C2077 SUNSAR_SAR8B_CV_0.D<4> VGND 11.8306f
C2078 SUNSAR_SAR8B_CV_0.D<5> VGND 12.7012f
C2079 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN0.D VGND 0.107643f
C2080 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN0.D VGND 0.107643f
C2081 SUNSAR_SAR8B_CV_0.D<6> VGND 12.0145f
C2082 SUNSAR_SAR8B_CV_0.D<7> VGND 17.833302f
C2083 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN0.D VGND 0.107643f
C2084 a_22790_41880# VGND 0.394408f $ **FLOATING
C2085 a_21422_41880# VGND 0.395138f $ **FLOATING
C2086 a_17750_41880# VGND 0.395707f $ **FLOATING
C2087 a_16382_41880# VGND 0.395707f $ **FLOATING
C2088 a_12710_41880# VGND 0.395707f $ **FLOATING
C2089 a_11342_41880# VGND 0.395707f $ **FLOATING
C2090 a_7670_41880# VGND 0.395707f $ **FLOATING
C2091 a_6302_41880# VGND 0.395707f $ **FLOATING
C2092 a_2630_41880# VGND 0.396052f $ **FLOATING
C2093 SUNSAR_CAPT8B_CV_0.SUNSAR_IVX1_CV_0.Y VGND 1.96193f
C2094 a_22790_42408# VGND 0.410698f $ **FLOATING
C2095 a_21422_42408# VGND 0.389697f $ **FLOATING
C2096 a_17750_42408# VGND 0.390266f $ **FLOATING
C2097 a_16382_42408# VGND 0.390266f $ **FLOATING
C2098 a_12710_42408# VGND 0.390266f $ **FLOATING
C2099 a_11342_42408# VGND 0.390266f $ **FLOATING
C2100 a_7670_42408# VGND 0.390266f $ **FLOATING
C2101 a_6302_42408# VGND 0.390266f $ **FLOATING
C2102 a_2630_42408# VGND 0.390612f $ **FLOATING
C2103 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C2104 SUNSAR_CAPT8B_CV_0.XI14.XA3.Y VGND 1.28758f
C2105 SUNSAR_CAPT8B_CV_0.XH13.XA3.Y VGND 1.27933f
C2106 SUNSAR_CAPT8B_CV_0.XG12.XA3.Y VGND 1.27933f
C2107 SUNSAR_CAPT8B_CV_0.XF11.XA3.Y VGND 1.27933f
C2108 SUNSAR_CAPT8B_CV_0.XE10.XA3.Y VGND 1.27933f
C2109 SUNSAR_CAPT8B_CV_0.XD09.XA3.Y VGND 1.27933f
C2110 SUNSAR_CAPT8B_CV_0.XC08.XA3.Y VGND 1.27933f
C2111 SUNSAR_CAPT8B_CV_0.XB07.XA3.Y VGND 1.29578f
C2112 a_22790_42760# VGND 0.378208f $ **FLOATING
C2113 a_21422_42760# VGND 0.393027f $ **FLOATING
C2114 a_17750_42760# VGND 0.393596f $ **FLOATING
C2115 a_16382_42760# VGND 0.393596f $ **FLOATING
C2116 a_12710_42760# VGND 0.393596f $ **FLOATING
C2117 a_11342_42760# VGND 0.393596f $ **FLOATING
C2118 a_7670_42760# VGND 0.393596f $ **FLOATING
C2119 a_6302_42760# VGND 0.393596f $ **FLOATING
C2120 a_2630_42760# VGND 0.393942f $ **FLOATING
C2121 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 24.712801f
C2122 SUNSAR_SAR8B_CV_0.EN VGND 11.0158f
C2123 a_22790_43112# VGND 0.388427f $ **FLOATING
C2124 SUNSAR_CAPT8B_CV_0.XI14.XA4.A VGND 1.29446f
C2125 SUNSAR_CAPT8B_CV_0.XH13.XA4.A VGND 1.29655f
C2126 SUNSAR_CAPT8B_CV_0.XG12.XA4.A VGND 1.29655f
C2127 SUNSAR_CAPT8B_CV_0.XF11.XA4.A VGND 1.29655f
C2128 SUNSAR_CAPT8B_CV_0.XE10.XA4.A VGND 1.29655f
C2129 SUNSAR_CAPT8B_CV_0.XD09.XA4.A VGND 1.29655f
C2130 SUNSAR_CAPT8B_CV_0.XC08.XA4.A VGND 1.29655f
C2131 SUNSAR_CAPT8B_CV_0.XB07.XA4.A VGND 1.29893f
C2132 SUNSAR_CAPT8B_CV_0.XA4.Y VGND 2.38165f
C2133 a_21422_43288# VGND 0.394124f $ **FLOATING
C2134 a_17750_43288# VGND 0.394693f $ **FLOATING
C2135 a_16382_43288# VGND 0.394693f $ **FLOATING
C2136 a_12710_43288# VGND 0.394693f $ **FLOATING
C2137 a_11342_43288# VGND 0.394693f $ **FLOATING
C2138 a_7670_43288# VGND 0.394693f $ **FLOATING
C2139 a_6302_43288# VGND 0.394693f $ **FLOATING
C2140 a_2630_43288# VGND 0.395039f $ **FLOATING
C2141 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN0.D VGND 0.103608f
C2142 SUNSAR_CAPT8B_CV_0.XA3.Y VGND 1.65429f
C2143 a_22790_43640# VGND 0.387806f $ **FLOATING
C2144 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN0.D VGND 0.112889f
C2145 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y VGND 2.60322f
C2146 SUNSAR_CAPT8B_CV_0.XI14.XA2.Y VGND 1.6954f
C2147 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN0.D VGND 0.112889f
C2148 SUNSAR_CAPT8B_CV_0.XH13.XA2.Y VGND 1.69797f
C2149 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y VGND 2.58593f
C2150 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN0.D VGND 0.112889f
C2151 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y VGND 2.6374f
C2152 SUNSAR_CAPT8B_CV_0.XG12.XA2.Y VGND 1.69797f
C2153 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN0.D VGND 0.112889f
C2154 SUNSAR_CAPT8B_CV_0.XF11.XA2.Y VGND 1.69797f
C2155 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y VGND 2.63726f
C2156 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN0.D VGND 0.112889f
C2157 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y VGND 2.59274f
C2158 SUNSAR_CAPT8B_CV_0.XE10.XA2.Y VGND 1.69797f
C2159 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN0.D VGND 0.112889f
C2160 SUNSAR_CAPT8B_CV_0.XD09.XA2.Y VGND 1.69797f
C2161 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y VGND 2.5926f
C2162 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN0.D VGND 0.112889f
C2163 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y VGND 2.6374f
C2164 SUNSAR_CAPT8B_CV_0.XC08.XA2.Y VGND 1.69797f
C2165 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN0.D VGND 0.112889f
C2166 SUNSAR_CAPT8B_CV_0.XB07.XA2.Y VGND 1.69726f
C2167 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y VGND 2.70316f
C2168 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.891538f
C2169 a_21422_43816# VGND 0.390629f $ **FLOATING
C2170 a_17750_43816# VGND 0.391198f $ **FLOATING
C2171 a_16382_43816# VGND 0.391198f $ **FLOATING
C2172 a_12710_43816# VGND 0.391198f $ **FLOATING
C2173 a_11342_43816# VGND 0.391198f $ **FLOATING
C2174 a_7670_43816# VGND 0.391198f $ **FLOATING
C2175 a_6302_43816# VGND 0.391198f $ **FLOATING
C2176 a_2630_43816# VGND 0.391544f $ **FLOATING
C2177 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 26.6958f
C2178 a_22790_43992# VGND 0.384235f $ **FLOATING
C2179 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.26356f
C2180 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.26291f
C2181 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.26291f
C2182 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.26291f
C2183 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26291f
C2184 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C2185 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C2186 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C2187 SUNSAR_CAPT8B_CV_0.XA2.MN0.G VGND 0.651712f
C2188 a_21422_44168# VGND 0.425534f $ **FLOATING
C2189 a_17750_44168# VGND 0.425449f $ **FLOATING
C2190 a_16382_44168# VGND 0.425864f $ **FLOATING
C2191 a_12710_44168# VGND 0.425449f $ **FLOATING
C2192 a_11342_44168# VGND 0.425864f $ **FLOATING
C2193 a_7670_44168# VGND 0.425449f $ **FLOATING
C2194 a_6302_44168# VGND 0.425864f $ **FLOATING
C2195 a_2630_44168# VGND 0.426034f $ **FLOATING
C2196 TIE_L VGND 6.84182f
C2197 a_22790_44344# VGND 0.423601f $ **FLOATING
.ends

