magic
tech sky130A
magscale 1 2
timestamp 1710669355
<< metal3 >>
rect -1986 17492 1986 17520
rect -1986 13868 1902 17492
rect 1966 13868 1986 17492
rect -1986 13840 1986 13868
rect -1986 13572 1986 13600
rect -1986 9948 1902 13572
rect 1966 9948 1986 13572
rect -1986 9920 1986 9948
rect -1986 9652 1986 9680
rect -1986 6028 1902 9652
rect 1966 6028 1986 9652
rect -1986 6000 1986 6028
rect -1986 5732 1986 5760
rect -1986 2108 1902 5732
rect 1966 2108 1986 5732
rect -1986 2080 1986 2108
rect -1986 1812 1986 1840
rect -1986 -1812 1902 1812
rect 1966 -1812 1986 1812
rect -1986 -1840 1986 -1812
rect -1986 -2108 1986 -2080
rect -1986 -5732 1902 -2108
rect 1966 -5732 1986 -2108
rect -1986 -5760 1986 -5732
rect -1986 -6028 1986 -6000
rect -1986 -9652 1902 -6028
rect 1966 -9652 1986 -6028
rect -1986 -9680 1986 -9652
rect -1986 -9948 1986 -9920
rect -1986 -13572 1902 -9948
rect 1966 -13572 1986 -9948
rect -1986 -13600 1986 -13572
rect -1986 -13868 1986 -13840
rect -1986 -17492 1902 -13868
rect 1966 -17492 1986 -13868
rect -1986 -17520 1986 -17492
<< via3 >>
rect 1902 13868 1966 17492
rect 1902 9948 1966 13572
rect 1902 6028 1966 9652
rect 1902 2108 1966 5732
rect 1902 -1812 1966 1812
rect 1902 -5732 1966 -2108
rect 1902 -9652 1966 -6028
rect 1902 -13572 1966 -9948
rect 1902 -17492 1966 -13868
<< mimcap >>
rect -1946 17440 1654 17480
rect -1946 13920 -1906 17440
rect 1614 13920 1654 17440
rect -1946 13880 1654 13920
rect -1946 13520 1654 13560
rect -1946 10000 -1906 13520
rect 1614 10000 1654 13520
rect -1946 9960 1654 10000
rect -1946 9600 1654 9640
rect -1946 6080 -1906 9600
rect 1614 6080 1654 9600
rect -1946 6040 1654 6080
rect -1946 5680 1654 5720
rect -1946 2160 -1906 5680
rect 1614 2160 1654 5680
rect -1946 2120 1654 2160
rect -1946 1760 1654 1800
rect -1946 -1760 -1906 1760
rect 1614 -1760 1654 1760
rect -1946 -1800 1654 -1760
rect -1946 -2160 1654 -2120
rect -1946 -5680 -1906 -2160
rect 1614 -5680 1654 -2160
rect -1946 -5720 1654 -5680
rect -1946 -6080 1654 -6040
rect -1946 -9600 -1906 -6080
rect 1614 -9600 1654 -6080
rect -1946 -9640 1654 -9600
rect -1946 -10000 1654 -9960
rect -1946 -13520 -1906 -10000
rect 1614 -13520 1654 -10000
rect -1946 -13560 1654 -13520
rect -1946 -13920 1654 -13880
rect -1946 -17440 -1906 -13920
rect 1614 -17440 1654 -13920
rect -1946 -17480 1654 -17440
<< mimcapcontact >>
rect -1906 13920 1614 17440
rect -1906 10000 1614 13520
rect -1906 6080 1614 9600
rect -1906 2160 1614 5680
rect -1906 -1760 1614 1760
rect -1906 -5680 1614 -2160
rect -1906 -9600 1614 -6080
rect -1906 -13520 1614 -10000
rect -1906 -17440 1614 -13920
<< metal4 >>
rect -198 17441 -94 17640
rect 1882 17492 1986 17640
rect -1907 17440 1615 17441
rect -1907 13920 -1906 17440
rect 1614 13920 1615 17440
rect -1907 13919 1615 13920
rect -198 13521 -94 13919
rect 1882 13868 1902 17492
rect 1966 13868 1986 17492
rect 1882 13572 1986 13868
rect -1907 13520 1615 13521
rect -1907 10000 -1906 13520
rect 1614 10000 1615 13520
rect -1907 9999 1615 10000
rect -198 9601 -94 9999
rect 1882 9948 1902 13572
rect 1966 9948 1986 13572
rect 1882 9652 1986 9948
rect -1907 9600 1615 9601
rect -1907 6080 -1906 9600
rect 1614 6080 1615 9600
rect -1907 6079 1615 6080
rect -198 5681 -94 6079
rect 1882 6028 1902 9652
rect 1966 6028 1986 9652
rect 1882 5732 1986 6028
rect -1907 5680 1615 5681
rect -1907 2160 -1906 5680
rect 1614 2160 1615 5680
rect -1907 2159 1615 2160
rect -198 1761 -94 2159
rect 1882 2108 1902 5732
rect 1966 2108 1986 5732
rect 1882 1812 1986 2108
rect -1907 1760 1615 1761
rect -1907 -1760 -1906 1760
rect 1614 -1760 1615 1760
rect -1907 -1761 1615 -1760
rect -198 -2159 -94 -1761
rect 1882 -1812 1902 1812
rect 1966 -1812 1986 1812
rect 1882 -2108 1986 -1812
rect -1907 -2160 1615 -2159
rect -1907 -5680 -1906 -2160
rect 1614 -5680 1615 -2160
rect -1907 -5681 1615 -5680
rect -198 -6079 -94 -5681
rect 1882 -5732 1902 -2108
rect 1966 -5732 1986 -2108
rect 1882 -6028 1986 -5732
rect -1907 -6080 1615 -6079
rect -1907 -9600 -1906 -6080
rect 1614 -9600 1615 -6080
rect -1907 -9601 1615 -9600
rect -198 -9999 -94 -9601
rect 1882 -9652 1902 -6028
rect 1966 -9652 1986 -6028
rect 1882 -9948 1986 -9652
rect -1907 -10000 1615 -9999
rect -1907 -13520 -1906 -10000
rect 1614 -13520 1615 -10000
rect -1907 -13521 1615 -13520
rect -198 -13919 -94 -13521
rect 1882 -13572 1902 -9948
rect 1966 -13572 1986 -9948
rect 1882 -13868 1986 -13572
rect -1907 -13920 1615 -13919
rect -1907 -17440 -1906 -13920
rect 1614 -17440 1615 -13920
rect -1907 -17441 1615 -17440
rect -198 -17640 -94 -17441
rect 1882 -17492 1902 -13868
rect 1966 -17492 1986 -13868
rect 1882 -17640 1986 -17492
<< properties >>
string FIXED_BBOX -1986 13840 1694 17520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17.999 l 17.999 val 661.674 carea 2.00 cperi 0.19 nx 1 ny 9 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
