* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[1] uio_oe[2]
*+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[1] uio_out[2] uio_out[3]
*+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7] uio_oe[0] ui_in[0]
*+ uo_out[6] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3] uio_out[0]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t7 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t8 VGND.t27 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR.t28 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA0.XA11.A VPWR.t212 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t0 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t10 VPWR.t22 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND.t486 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA4.CP0.t1 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND.t153 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t5 VPWR.t558 VPWR.t557 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND.t540 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t8 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR.t213 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND.t499 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t1 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t29 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t8 VPWR.t593 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR.t589 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t5 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND.t66 VGND.t63 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR.t77 VPWR.t74 VPWR.t76 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.D<3>.t8 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND.t518 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t23 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t3 VPWR.t543 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND.t464 clk.t0 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR.t570 SUNSAR_SAR8B_CV_0.XA3.CN1.t8 SUNSAR_SAR8B_CV_0.D<4>.t7 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND.t69 VGND.t67 VGND.t68 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR.t84 VPWR.t82 VPWR.t83 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND.t12 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND.t476 SUNSAR_SAR8B_CV_0.D<7>.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t0 VGND.t475 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5>.t4 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t9 VPWR.t432 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t59 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1.t1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t2 VGND.t424 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR.t11 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR.t489 SUNSAR_SAR8B_CV_0.XA6.CN1.t8 SUNSAR_SAR8B_CV_0.D<1>.t6 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND.t421 SUNSAR_SAR8B_CV_0.XA6.CN1.t10 SUNSAR_SAR8B_CV_0.D<1>.t1 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1.t4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t4 VPWR.t494 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA6.A VGND.t21 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VPWR.t216 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR.t224 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND.t491 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t1 VGND.t490 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t7 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t9 VPWR.t458 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VGND.t166 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t13 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR.t468 SUNSAR_SAR8B_CV_0.XA6.CP0.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t5 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5>.t5 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t10 VPWR.t433 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND.t442 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA5.CN1.t1 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR.t511 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA5.CN1.t6 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VPWR.t501 SUNSAR_SAR8B_CV_0.DONE.t11 tt_um_TT06_SAR_done_0.x3.MP1.G VPWR.t500 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X51 VGND.t388 SUNSAR_SAR8B_CV_0.XA7.CP0.t8 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X52 SUNSAR_SAR8B_CV_0.XB1.CKN.t0 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t2 VGND.t352 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 VPWR.t542 SUNSAR_SAR8B_CV_0.EN.t57 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_SAR8B_CV_0.XA7.CN1.t2 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t5 VGND.t425 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR.t237 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X56 VPWR.t455 SUNSAR_SAR8B_CV_0.XA7.CP0.t10 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP.t11 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X58 SUNSAR_SAR8B_CV_0.XA7.CN1.t6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t6 VPWR.t495 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND.t176 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<7>.t12 VGND.t480 VGND.t479 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR.t242 VPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X63 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<1>.t11 VPWR.t513 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X65 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VGND.t180 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X66 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR.t247 VPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t19 VGND.t436 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t19 VGND.t549 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t33 VPWR.t531 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VPWR.t248 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR.t225 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X72 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X74 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND.t191 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t35 VGND.t529 VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X76 VGND.t396 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X77 ua[1].t4 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP.t3 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X78 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t55 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X79 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR.t253 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t0 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND.t182 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S uo_out[3].t2 VGND.t379 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t9 SUNSAR_SAR8B_CV_0.XA6.XA9.B VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND.t193 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t2 VGND.t385 VGND.t384 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t13 VGND.t431 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.ENO.t2 VGND.t359 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t17 VPWR.t504 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X88 VPWR.t255 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.t1 VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t21 VPWR.t529 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X90 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND.t197 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND.t198 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t3 VPWR.t435 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X93 VGND.t135 VGND.t132 VGND.t134 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND.t115 VGND.t113 VGND.t114 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X95 VGND.t337 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA3.CP0.t1 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X96 VPWR.t123 VPWR.t120 VPWR.t122 VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X97 ua[1].t8 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t6 SUNSAR_SAR8B_CV_0.SARN VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X98 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP.t13 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X99 VPWR.t261 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X100 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t53 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X101 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t23 SUNSAR_SAR8B_CV_0.XA3.EN VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND.t201 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t21 VGND.t437 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR.t262 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X106 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t0 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t5 VGND.t401 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X107 uo_out[0].t0 SUNSAR_CAPT8B_CV_0.XI14.QN VGND.t158 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X108 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t1 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t6 VPWR.t485 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R8 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X109 VGND.t37 VGND.t34 VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND.t90 VGND.t87 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 VGND.t62 VGND.t60 VGND.t61 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND.t202 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t1 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t11 VGND.t393 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X114 VPWR.t446 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t10 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t3 VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X115 VPWR.t147 VPWR.t144 VPWR.t146 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X116 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA11.A VPWR.t263 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND.t204 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X118 VGND.t23 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X119 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND.t195 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X120 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X121 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t13 VGND.t510 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X122 VGND.t322 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t0 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<6>.t8 VPWR.t413 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X124 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t3 SUNSAR_SAR8B_CV_0.D<7>.t13 VPWR.t576 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X125 VGND.t122 VGND.t119 VGND.t121 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t33 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t1 SUNSAR_SAR8B_CV_0.XA3.CP0.t10 VGND.t343 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.D<2>.t8 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t2 VGND.t443 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X130 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t8 VPWR.t487 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X131 VPWR.t403 SUNSAR_SAR8B_CV_0.XA4.CN1.t8 SUNSAR_SAR8B_CV_0.D<3>.t0 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X132 VGND.t327 SUNSAR_SAR8B_CV_0.XA4.CN1.t10 SUNSAR_SAR8B_CV_0.D<3>.t2 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR.t268 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X134 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X135 VGND.t141 VGND.t139 VGND.t140 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X136 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t27 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X137 VPWR.t448 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t11 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t4 VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VGND.t319 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA3.CN1.t1 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 VPWR.t274 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t5 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t11 VPWR.t587 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.EN.t31 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 VPWR.t599 SUNSAR_SAR8B_CV_0.XA4.CP0.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t5 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X146 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t5 SUNSAR_SAR8B_CV_0.D<7>.t15 VPWR.t577 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X147 VGND.t33 VGND.t30 VGND.t32 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X148 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND.t205 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X149 VPWR.t395 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA3.CN1.t2 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X150 VGND.t112 VGND.t109 VGND.t111 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VPWR.t266 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t1 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t4 VPWR.t400 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA1.ENO.t3 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X155 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<3>.t9 VPWR.t579 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VGND.t170 VGND.t169 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 VGND.t159 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA6.CN1.t1 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X158 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA1.ENO.t4 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND.t155 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R10 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X160 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR.t214 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR.t270 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VPWR.t304 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X163 VGND.t457 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t0 VGND.t456 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t51 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X166 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t5 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t12 VGND.t382 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X167 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t9 SUNSAR_SAR8B_CV_0.XA4.XA9.B VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 VPWR.t409 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA6.CP0.t1 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X169 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.ENO.t2 VGND.t330 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t21 VGND.t550 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 VPWR.t460 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t12 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t5 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t5 VPWR.t401 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X174 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.ENO.t4 VPWR.t407 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X175 VPWR.t143 VPWR.t140 VPWR.t142 VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X176 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X177 VGND.t297 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA7.CP0.t0 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X178 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t15 VPWR.t526 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X181 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND.t175 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X182 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t4 VPWR.t457 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X183 VGND.t73 VGND.t70 VGND.t72 VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 VPWR.t358 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA7.CP0.t2 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X185 VGND.t138 VGND.t136 VGND.t137 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X186 ua[1].t0 SUNSAR_SAR8B_CV_0.XB1.CKN.t4 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t2 VPWR.t472 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t49 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X188 VPWR.t132 VPWR.t130 VPWR.t131 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t21 SUNSAR_SAR8B_CV_0.XA1.EN VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t15 VGND.t433 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 VGND.t47 VGND.t45 VGND.t46 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X193 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t25 VGND.t553 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X194 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X195 VGND.t516 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t21 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR.t307 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 VPWR.t236 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X198 SUNSAR_SAR8B_CV_0.XA5.ENO.t1 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND.t250 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X199 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t0 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t14 VGND.t495 VGND.t494 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 VPWR.t312 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R13 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X201 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND.t179 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t4 SUNSAR_SAR8B_CV_0.XA6.CP0.t11 VPWR.t470 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP.t15 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X205 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t5 VGND.t397 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X206 VGND.t417 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.D<7>.t2 VGND.t416 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R14 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X207 VGND.t59 VGND.t56 VGND.t58 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND.t253 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 VPWR.t220 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA6.CN1.t2 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t3 VGND.t306 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.D<4>.t9 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X212 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.t0 SUNSAR_SAR8B_CV_0.XB1.CKN.t5 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X213 VGND.t213 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R15 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X214 VGND.t108 VGND.t105 VGND.t107 VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t31 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X216 uo_out[5].t1 SUNSAR_CAPT8B_CV_0.XD09.QN VPWR.t271 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t31 VGND.t526 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.XA3.CP0.t2 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t5 VGND.t338 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 SUNSAR_SAR8B_CV_0.D<6>.t0 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t11 VGND.t468 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.D<6>.t7 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t13 VPWR.t569 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X221 VPWR.t173 VPWR.t171 VPWR.t172 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t15 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R16 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X223 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP.t10 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t2 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t10 VPWR.t385 VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X225 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND.t256 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND.t257 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X228 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t6 VGND.t398 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X229 VGND.t439 SUNSAR_SAR8B_CV_0.XA5.CN1.t11 SUNSAR_SAR8B_CV_0.D<2>.t0 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X230 VPWR.t387 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t11 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t4 VPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR.t319 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X232 VPWR.t508 SUNSAR_SAR8B_CV_0.XA5.CN1.t12 SUNSAR_SAR8B_CV_0.D<2>.t7 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X233 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND.t177 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X235 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X236 VPWR.t604 VGND.t2 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X237 VPWR.t43 VPWR.t40 VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VPWR.t313 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X239 VPWR.t267 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t29 VGND.t524 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t4 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t15 VGND.t26 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA1.ENO.t5 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t2 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t14 VPWR.t24 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.D<7>.t3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t5 VPWR.t479 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X246 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.EN.t29 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND.t452 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 VGND.t285 SUNSAR_SAR8B_CV_0.XA5.CP0.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t2 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.XA3.CP0.t0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t6 VGND.t339 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 VPWR.t346 SUNSAR_SAR8B_CV_0.XA5.CP0.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t4 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 SUNSAR_SAR8B_CV_0.D<6>.t2 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t14 VGND.t469 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.D<6>.t4 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t8 VPWR.t566 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 VGND.t309 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA4.CN1.t1 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X253 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t47 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND.t255 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X255 ua[0].t6 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.EN.t19 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t0 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t6 VPWR.t560 VPWR.t559 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND.t190 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t0 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t4 VGND.t307 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR.t252 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VPWR.t249 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X263 VPWR.t538 SUNSAR_SAR8B_CV_0.EN.t45 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S uo_out[0].t2 VGND.t341 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X266 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<2>.t11 VGND.t163 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X268 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<2>.t10 VPWR.t223 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 VPWR.t582 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA4.CP0.t5 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X270 ua[0].t1 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t7 SUNSAR_SAR8B_CV_0.SARP.t6 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_SAR8B_CV_0.D<7>.t5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t7 VPWR.t481 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.ENO.t4 VPWR.t436 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t28 VGND.t537 VGND.t536 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND.t199 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X275 VGND.t86 VGND.t84 VGND.t85 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X276 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND.t260 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 VPWR.t585 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t6 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X278 uio_oe[0].t0 tt_um_TT06_SAR_done_0.x4.MP0.G VPWR.t330 VPWR.t329 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR.t322 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R17 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X280 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t27 VPWR.t530 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X282 VPWR.t565 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t9 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t19 VGND.t514 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X284 VPWR.t96 VPWR.t93 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t9 SUNSAR_SAR8B_CV_0.XA5.XA9.B VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R18 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R19 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X286 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VGND.t244 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t25 VGND.t373 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t1 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR.t332 VPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t2 VGND.t294 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t43 VPWR.t537 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X292 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t4 VPWR.t354 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR.t327 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X294 VPWR.t308 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t31 VGND.t378 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t5 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t12 VGND.t314 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t60 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X300 uio_out[0].t1 tt_um_TT06_SAR_done_0.x3.MP1.G VPWR.t235 VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t17 SUNSAR_SAR8B_CV_0.XA1.ENO.t1 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t4 SUNSAR_SAR8B_CV_0.XA4.CP0.t12 VPWR.t601 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t2 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t6 VGND.t459 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR.t462 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t0 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VGND.t449 SUNSAR_SAR8B_CV_0.XA7.CN1.t14 SUNSAR_SAR8B_CV_0.D<0>.t1 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND.t150 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X307 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND.t152 VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X308 SUNSAR_SAR8B_CV_0.XA6.CP0.t3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t5 VPWR.t411 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X309 VPWR.t515 SUNSAR_SAR8B_CV_0.XA7.CN1.t8 SUNSAR_SAR8B_CV_0.D<0>.t6 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X310 VPWR.t375 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA4.CN1.t2 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X311 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP.t9 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X312 VPWR.t139 VPWR.t136 VPWR.t138 VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X313 VPWR.t230 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X314 VGND.t156 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA6.XA11.A VPWR.t250 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X316 uo_out[7].t1 SUNSAR_CAPT8B_CV_0.XB07.QN VPWR.t251 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t27 VGND.t522 VGND.t521 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X318 VPWR.t483 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t8 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 ua[1].t1 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP.t0 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR.t168 VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X321 VPWR.t191 VPWR.t189 VPWR.t190 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X322 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t37 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<1>.t10 VPWR.t512 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X324 VGND.t44 VGND.t42 VGND.t43 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t2 VGND.t455 VGND.t454 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR.t572 SUNSAR_SAR8B_CV_0.XA3.CN1.t12 SUNSAR_SAR8B_CV_0.D<4>.t6 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 VGND.t541 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t11 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X328 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B SUNSAR_SAR8B_CV_0.XB2.CKN.t3 VGND.t301 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t10 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XA6.CP0.t4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t6 VPWR.t412 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 VPWR.t316 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.D<5>.t2 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t14 VGND.t356 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X333 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.EN.t41 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR.t336 VPWR.t335 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X337 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND.t18 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X338 VGND.t423 SUNSAR_SAR8B_CV_0.XA6.CN1.t13 SUNSAR_SAR8B_CV_0.D<1>.t3 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t25 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<5>.t11 VGND.t462 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X341 VPWR.t423 SUNSAR_SAR8B_CV_0.XA3.CP0.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t7 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X342 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.EN.t39 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND.t157 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X344 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t3 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t8 VGND.t392 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X346 ua[1].t9 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t9 SUNSAR_SAR8B_CV_0.SARN VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X347 SUNSAR_SAR8B_CV_0.D<4>.t0 SUNSAR_SAR8B_CV_0.XA3.CN1.t13 VGND.t473 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X348 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t2 VGND.t498 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X349 VPWR.t527 SUNSAR_SAR8B_CV_0.EN.t17 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t8 VPWR.t592 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R23 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X351 VGND.t405 SUNSAR_SAR8B_CV_0.XA6.CP0.t14 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t3 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X352 VPWR.t556 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t4 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR.t555 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<4>.t11 VGND.t463 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND.t194 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_SAR8B_CV_0.D<5>.t0 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t15 VGND.t357 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<4>.t10 VPWR.t549 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 VPWR.t39 VPWR.t36 VPWR.t38 VPWR.t37 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X359 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND.t216 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X360 VGND.t406 SUNSAR_SAR8B_CV_0.XB1.CKN.t2 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND.t174 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t2 VGND.t400 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.ENO.t6 VGND.t331 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R24 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X364 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X365 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR.t334 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X366 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.ENO.t7 VPWR.t408 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t2 SUNSAR_SAR8B_CV_0.XA3.CP0.t14 VGND.t344 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X368 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t37 VPWR.t534 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t9 VGND.t430 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R25 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X370 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<1>.t8 VGND.t446 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X371 VGND.t290 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA5.CP0.t1 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X372 SUNSAR_SAR8B_CV_0.D<4>.t3 SUNSAR_SAR8B_CV_0.XA3.CN1.t14 VGND.t474 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R26 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X373 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t9 SUNSAR_SAR8B_CV_0.XA3.XA9.B VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X374 VGND.t29 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t6 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X375 VPWR.t348 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA5.CP0.t2 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X376 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t0 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t9 VGND.t501 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X377 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VGND.t183 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X378 VPWR.t25 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t12 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t3 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X379 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t6 VPWR.t590 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND.t164 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X381 VPWR.t159 VPWR.t156 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X382 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND.t386 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S uo_out[5].t2 VPWR.t356 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X384 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t5 VGND.t346 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X385 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R27 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X386 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t2 VPWR.t424 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X387 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND.t212 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 VPWR.t602 VGND.t0 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X389 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X390 VGND.t101 VGND.t99 VGND.t100 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X391 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t25 VGND.t520 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t23 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X393 VPWR.t204 VPWR.t202 VPWR.t203 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X394 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X395 VGND.t51 VGND.t48 VGND.t50 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t28 VGND.t376 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t5 VGND.t358 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE.t17 VGND.t512 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND.t217 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X400 VPWR.t546 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t4 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR.t278 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X402 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND.t200 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XA4.CP0.t6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t6 VPWR.t583 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X404 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t13 VGND.t364 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X407 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t3 SUNSAR_SAR8B_CV_0.XA5.CP0.t13 VGND.t288 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA4.XA11.A VPWR.t303 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t7 SUNSAR_SAR8B_CV_0.XA5.CP0.t14 VPWR.t361 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X410 VPWR.t514 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t9 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t11 VGND.t363 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t0 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t7 VGND.t380 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R29 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R30 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X413 SUNSAR_SAR8B_CV_0.EN.t1 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t11 VPWR.t595 VPWR.t594 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X414 VPWR.t553 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t2 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR.t552 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 VGND.t349 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA5.CN1.t0 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X416 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<3>.t10 VPWR.t580 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X417 VPWR.t425 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA5.CN1.t7 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X418 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t16 VGND.t369 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X419 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.DONE.t7 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X420 uo_out[6].t0 SUNSAR_CAPT8B_CV_0.XC08.QN VGND.t248 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X421 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0].t0 VPWR.t20 VPWR.t19 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X422 uo_out[6].t1 SUNSAR_CAPT8B_CV_0.XC08.QN VPWR.t309 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X423 SUNSAR_SAR8B_CV_0.XA4.CP0.t7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t2 VPWR.t581 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X424 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t4 SUNSAR_SAR8B_CV_0.D<7>.t14 VGND.t482 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X425 VGND.t76 VGND.t74 VGND.t75 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X426 VPWR.t35 VPWR.t33 VPWR.t34 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X427 VPWR.t163 VPWR.t160 VPWR.t162 VPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X428 VPWR.t431 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t8 SUNSAR_SAR8B_CV_0.D<5>.t7 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R31 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X429 VGND.t426 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA7.CN1.t0 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND.t207 VGND.t206 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 VGND.t329 SUNSAR_SAR8B_CV_0.XA4.CN1.t13 SUNSAR_SAR8B_CV_0.D<3>.t5 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.D<1>.t5 SUNSAR_SAR8B_CV_0.XA6.CN1.t14 VPWR.t491 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X433 VPWR.t496 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA7.CN1.t7 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X434 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t10 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X435 VGND.t546 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t16 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X436 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t1 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR.t311 VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X437 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR.t306 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t3 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t12 VGND.t493 VGND.t492 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R32 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X440 VPWR.t32 VPWR.t29 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X441 VPWR.t606 VGND.t4 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X442 VGND.t535 SUNSAR_SAR8B_CV_0.XA4.CP0.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t3 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X443 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t7 SUNSAR_SAR8B_CV_0.XA6.CP0.t15 VPWR.t471 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 VPWR.t181 VPWR.t178 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t3 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t14 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t6 SUNSAR_SAR8B_CV_0.D<7>.t16 VGND.t484 VGND.t483 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X447 VGND.t545 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X449 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R34 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X450 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t11 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X452 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t6 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X453 SUNSAR_SAR8B_CV_0.D<1>.t4 SUNSAR_SAR8B_CV_0.XA6.CN1.t15 VPWR.t492 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X454 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X455 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP.t8 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X457 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.ENO.t5 VPWR.t437 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X458 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t7 VGND.t324 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X459 VPWR.t521 SUNSAR_SAR8B_CV_0.EN.t4 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 VPWR.t66 VPWR.t63 VPWR.t65 VPWR.t64 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X462 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X463 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<3>.t11 VGND.t485 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 VPWR.t415 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA3.CP0.t7 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R35 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X465 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND.t210 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VGND.t243 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t14 VGND.t544 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X468 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S uo_out[7].t2 VPWR.t367 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 SUNSAR_SAR8B_CV_0.XB2.CKN.t1 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t3 VPWR.t428 VPWR.t427 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X470 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t20 VPWR.t528 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X471 SUNSAR_SAR8B_CV_0.XA3.CN1.t4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t6 VGND.t321 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X472 uo_out[0].t1 SUNSAR_CAPT8B_CV_0.XI14.QN VPWR.t217 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X473 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND.t178 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X474 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t7 VGND.t507 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 VGND.t332 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA6.CP0.t0 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R36 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X477 VPWR.t177 VPWR.t174 VPWR.t176 VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X478 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR.t239 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X479 VPWR.t104 VPWR.t101 VPWR.t103 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X480 VGND.t394 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t14 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t0 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X481 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t8 VGND.t325 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X482 SUNSAR_SAR8B_CV_0.XB2.CKN.t0 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t4 VGND.t353 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t15 VGND.t368 VGND.t367 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t6 VGND.t391 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP.t14 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X486 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t8 VPWR.t498 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR.t257 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 VGND.t261 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X489 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t2 VPWR.t519 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X491 VGND.t125 VGND.t123 VGND.t124 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X492 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X493 ua[0].t5 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X494 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t14 VGND.t366 VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA3.CN1.t0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t2 VGND.t318 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X496 VGND.t342 SUNSAR_SAR8B_CV_0.XA3.CP0.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t3 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t4 SUNSAR_SAR8B_CV_0.XA3.CP0.t12 VPWR.t422 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X498 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t8 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X499 VPWR.t488 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t4 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X500 VGND.t445 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t7 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R37 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X501 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X502 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t8 SUNSAR_SAR8B_CV_0.XA7.EN VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X503 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND.t245 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.D<0>.t10 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X505 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR.t256 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X506 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t4 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t15 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA5.CP0.t0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t2 VGND.t289 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X508 SUNSAR_SAR8B_CV_0.XA5.CP0.t6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t8 VPWR.t351 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 VPWR.t397 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA3.CN1.t6 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R38 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X510 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND.t267 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X511 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t1 SUNSAR_SAR8B_CV_0.XA6.CP0.t13 VGND.t404 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X512 VPWR.t151 VPWR.t148 VPWR.t150 VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X513 VPWR.t155 VPWR.t152 VPWR.t154 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X514 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA11.A VPWR.t328 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X515 VGND.t515 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t20 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X516 VPWR.t26 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t9 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X517 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t2 VGND.t502 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X519 VPWR.t574 SUNSAR_SAR8B_CV_0.D<7>.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t1 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X520 VGND.t161 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA6.CN1.t4 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X521 VPWR.t184 VPWR.t182 VPWR.t183 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X522 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<2>.t9 VPWR.t218 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND.t224 VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 SUNSAR_SAR8B_CV_0.D<3>.t6 SUNSAR_SAR8B_CV_0.XA4.CN1.t14 VPWR.t405 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X525 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VPWR.t284 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X526 ua[0].t3 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t4 SUNSAR_SAR8B_CV_0.SARP.t4 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X527 VGND.t539 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t30 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X528 SUNSAR_SAR8B_CV_0.XA5.CP0.t7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t9 VGND.t292 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 VPWR.t607 VGND.t5 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X530 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR.t326 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.CP0.t4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t6 VPWR.t349 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X532 VGND.t94 VGND.t91 VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R39 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X533 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t26 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t2 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t7 VGND.t284 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S VGND.t186 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X536 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t5 VGND.t308 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X537 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t7 SUNSAR_SAR8B_CV_0.XA4.CP0.t8 VPWR.t598 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t28 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X540 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND.t215 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X541 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t44 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.D<3>.t7 SUNSAR_SAR8B_CV_0.XA4.CN1.t15 VPWR.t406 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X544 SUNSAR_SAR8B_CV_0.D<7>.t0 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t2 VGND.t413 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X545 VPWR.t525 SUNSAR_SAR8B_CV_0.EN.t12 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND.t220 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t3 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t5 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X548 VPWR.t402 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t7 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO.t2 VGND.t280 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO.t3 VPWR.t341 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA5.ENO.t8 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA6.CN1.t0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t2 VPWR.t219 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R41 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X553 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X554 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VGND.t184 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA5.ENO.t5 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X557 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t40 VPWR.t536 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X558 ua[1].t6 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t2 SUNSAR_SAR8B_CV_0.SARN VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 VPWR.t88 VPWR.t85 VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X560 VGND.t488 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA4.CP0.t3 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X561 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t24 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X562 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR.t286 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 VGND.t497 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t2 VGND.t496 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X564 SUNSAR_SAR8B_CV_0.D<7>.t7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t9 VGND.t419 VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X565 ua[1].t3 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP.t2 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 VPWR.t5 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t0 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X567 SUNSAR_SAR8B_CV_0.XA7.ENO.t1 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND.t229 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X568 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S uo_out[6].t2 VGND.t282 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 VPWR.t47 VPWR.t44 VPWR.t46 VPWR.t45 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X570 VPWR.t288 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X571 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t18 VGND.t548 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X572 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S uo_out[6].t3 VPWR.t343 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X573 VPWR.t469 SUNSAR_SAR8B_CV_0.XA6.CP0.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t6 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X574 SUNSAR_SAR8B_CV_0.XA6.CN1.t6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t8 VPWR.t222 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X575 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t10 VPWR.t499 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_CAPT8B_CV_0.XA2.MP0.G SUNSAR_CAPT8B_CV_0.XA2.MP0.G VPWR.t290 VPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X578 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t36 VPWR.t533 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X579 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X580 VGND.t98 VGND.t95 VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X581 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t0 VPWR.t199 VPWR.t201 VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X582 ua[1].t7 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t3 SUNSAR_SAR8B_CV_0.SARN VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X583 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S SUNSAR_CAPT8B_CV_0.XA6.A VPWR.t16 VPWR.t15 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X584 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t2 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t9 VPWR.t444 VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t22 SUNSAR_SAR8B_CV_0.XA5.EN VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND.t265 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X587 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR.t337 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X588 SUNSAR_SAR8B_CV_0.XA3.CP0.t6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t9 VPWR.t418 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X589 VPWR.t603 VGND.t1 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X590 ua[1].t5 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XA3.B.t3 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X591 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t1 SUNSAR_SAR8B_CV_0.XA4.CP0.t13 VGND.t533 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X592 VPWR.t188 VPWR.t185 VPWR.t187 VPWR.t186 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X593 VPWR.t167 VPWR.t164 VPWR.t166 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X594 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA11.A VPWR.t318 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X595 VGND.t399 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t6 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R42 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X596 VGND.t450 SUNSAR_SAR8B_CV_0.XA7.CN1.t15 SUNSAR_SAR8B_CV_0.D<0>.t3 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X598 SUNSAR_SAR8B_CV_0.XA6.CP0.t7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t9 VGND.t335 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VPWR.t518 SUNSAR_SAR8B_CV_0.XA7.CN1.t13 SUNSAR_SAR8B_CV_0.D<0>.t4 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 VGND.t311 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA4.CN1.t4 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X601 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<4>.t8 VPWR.t484 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X602 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R43 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X603 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X604 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND.t185 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X605 VPWR.t285 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X606 uo_out[7].t0 SUNSAR_CAPT8B_CV_0.XB07.QN VGND.t189 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.D<5>.t10 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VGND.t519 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t24 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X609 VGND.t165 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X610 VGND.t340 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA3.CP0.t3 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 SUNSAR_SAR8B_CV_0.XA3.CP0.t5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t4 VPWR.t416 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 VGND.t390 SUNSAR_SAR8B_CV_0.XA7.CP0.t13 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X613 VGND.t470 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t15 SUNSAR_SAR8B_CV_0.D<6>.t3 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X614 VGND.t131 VGND.t129 VGND.t130 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t9 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X616 uo_out[1].t1 SUNSAR_CAPT8B_CV_0.XH13.QN VPWR.t279 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t22 VGND.t517 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X618 VPWR.t478 SUNSAR_SAR8B_CV_0.XA7.CP0.t14 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X619 VPWR.t567 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t10 SUNSAR_SAR8B_CV_0.D<6>.t6 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.D<2>.t3 SUNSAR_SAR8B_CV_0.XA5.CN1.t15 VGND.t441 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X621 VPWR.t389 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t15 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t4 VPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.D<2>.t5 SUNSAR_SAR8B_CV_0.XA5.CN1.t8 VPWR.t506 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t22 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X624 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S uo_out[0].t3 VPWR.t419 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB1.CKN.t7 VGND.t408 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X626 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND.t218 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA6.CP0.t6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t8 VGND.t334 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 VPWR.t371 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t7 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR.t370 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR.t277 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X631 VGND.t525 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t30 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<0>.t11 VGND.t293 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VPWR.t315 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t1 SUNSAR_SAR8B_CV_0.XA5.CP0.t9 VGND.t286 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 VPWR.t480 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.D<7>.t4 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA5.ENO.t3 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X637 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t6 SUNSAR_SAR8B_CV_0.XA5.CP0.t15 VPWR.t362 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND.t233 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_SAR8B_CV_0.XA4.CN1.t0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t2 VPWR.t374 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X640 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.XA3.ENO.t6 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR.t292 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R44 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X642 VPWR.t207 VPWR.t205 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_SAR8B_CV_0.D<2>.t2 SUNSAR_SAR8B_CV_0.XA5.CN1.t13 VGND.t440 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X644 SUNSAR_SAR8B_CV_0.D<2>.t4 SUNSAR_SAR8B_CV_0.XA5.CN1.t10 VPWR.t507 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X645 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA3.ENO.t7 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t18 VGND.t513 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X647 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X648 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA9.B VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X649 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X650 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR.t240 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X652 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t54 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X653 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t7 VGND.t295 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R46 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X654 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t12 VGND.t542 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X656 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X657 VGND.t283 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t5 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t0 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X658 VPWR.t600 SUNSAR_SAR8B_CV_0.XA4.CP0.t11 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t6 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 SUNSAR_SAR8B_CV_0.XA4.CN1.t6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t8 VPWR.t377 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t30 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X661 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VPWR.t245 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X663 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t1 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t8 VPWR.t373 VPWR.t372 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X664 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X665 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X666 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND.t237 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R48 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X667 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR.t297 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X669 VPWR.t452 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t16 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t1 VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X670 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t2 VGND.t409 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t20 VPWR.t505 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t18 VGND.t370 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X674 VPWR.t100 VPWR.t97 VPWR.t99 VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X675 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t46 VPWR.t539 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X676 VPWR.t551 clk.t1 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR.t550 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VPWR.t273 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 VGND.t461 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t1 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t9 VGND.t361 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X680 VPWR.t81 VPWR.t78 VPWR.t80 VPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X681 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t12 SUNSAR_SAR8B_CV_0.XA5.ENO.t0 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X682 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND.t221 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X683 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR.t282 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X684 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB1.TIE_L.t8 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X685 SUNSAR_SAR8B_CV_0.XA4.CP0.t2 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t9 VGND.t489 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X686 VPWR.t410 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA6.CP0.t2 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X687 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VPWR.t14 VPWR.t13 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X688 VPWR.t129 VPWR.t127 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 VGND.t145 VGND.t142 VGND.t144 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X690 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND.t242 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X691 VPWR.t58 VPWR.t55 VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t9 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X693 VGND.t531 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t36 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X694 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t0 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND.t270 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X695 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VPWR.t227 VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R49 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X696 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t7 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t16 VPWR.t391 VPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X697 uo_out[3].t1 SUNSAR_CAPT8B_CV_0.XF11.QN VPWR.t283 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t14 VGND.t511 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X699 VPWR.t467 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t8 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X700 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X701 SUNSAR_SAR8B_CV_0.D<4>.t5 SUNSAR_SAR8B_CV_0.XA3.CN1.t15 VPWR.t573 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.XA4.CP0.t0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t5 VGND.t487 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR.t258 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X704 VPWR.t434 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t12 SUNSAR_SAR8B_CV_0.D<5>.t6 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X705 VGND.t354 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t11 SUNSAR_SAR8B_CV_0.D<5>.t1 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X706 VGND.t552 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t24 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X707 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t20 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t8 VPWR.t564 VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X709 VGND.t429 SUNSAR_SAR8B_CV_0.DONE.t6 tt_um_TT06_SAR_done_0.x3.MP1.G VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X710 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR.t275 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VPWR.t333 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 VPWR.t293 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X713 SUNSAR_SAR8B_CV_0.D<1>.t0 SUNSAR_SAR8B_CV_0.XA6.CN1.t9 VGND.t420 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X714 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA3.ENO.t8 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X715 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X716 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t5 SUNSAR_SAR8B_CV_0.XA3.CP0.t11 VPWR.t421 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X717 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X718 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X719 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO.t4 VGND.t281 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X720 SUNSAR_SAR8B_CV_0.XB1.CKN.t1 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t5 VPWR.t430 VPWR.t429 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X721 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t5 VPWR.t477 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X722 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND.t246 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO.t5 VPWR.t342 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 ua[0].t2 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t10 SUNSAR_SAR8B_CV_0.SARP.t7 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 VPWR.t461 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t4 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R51 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X726 VPWR.t605 VGND.t3 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X727 VGND.t472 SUNSAR_SAR8B_CV_0.XA3.CN1.t11 SUNSAR_SAR8B_CV_0.D<4>.t1 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X728 SUNSAR_SAR8B_CV_0.D<4>.t4 SUNSAR_SAR8B_CV_0.XA3.CN1.t10 VPWR.t571 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X729 VGND.t298 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA7.CP0.t3 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X730 VGND.t500 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t2 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X731 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t1 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND.t274 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X732 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t0 SUNSAR_SAR8B_CV_0.XA6.CP0.t12 VGND.t403 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 VPWR.t359 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA7.CP0.t4 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X734 VPWR.t591 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t4 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X735 ua[0].t7 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR.t287 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 SUNSAR_SAR8B_CV_0.XA5.CN1.t3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t9 VGND.t351 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X738 SUNSAR_SAR8B_CV_0.XA5.CN1.t5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t8 VPWR.t426 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR.t272 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X740 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X741 SUNSAR_SAR8B_CV_0.D<1>.t2 SUNSAR_SAR8B_CV_0.XA6.CN1.t11 VGND.t422 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X742 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<5>.t9 VPWR.t548 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 VGND.t55 VGND.t52 VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X745 VPWR.t62 VPWR.t59 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X746 VPWR.t73 VPWR.t70 VPWR.t72 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X747 ua[0].t0 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t5 SUNSAR_SAR8B_CV_0.SARP.t5 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VPWR.t231 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X749 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR.t12 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X751 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X752 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t14 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X753 SUNSAR_SAR8B_CV_0.DONE.t0 SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND.t240 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R53 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X754 VGND.t41 VGND.t38 VGND.t40 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X755 SUNSAR_SAR8B_CV_0.DONE.t1 SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR.t298 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S uo_out[7].t3 VGND.t305 VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t9 SUNSAR_SAR8B_CV_0.XA2.XA9.B VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 VGND.t287 SUNSAR_SAR8B_CV_0.XA5.CP0.t12 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t0 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X759 SUNSAR_SAR8B_CV_0.XA5.CN1.t2 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t7 VGND.t350 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X760 VPWR.t364 SUNSAR_SAR8B_CV_0.XB2.CKN.t2 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 VPWR.t347 SUNSAR_SAR8B_CV_0.XA5.CP0.t11 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t5 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X762 SUNSAR_SAR8B_CV_0.XA5.CN1.t4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t3 VPWR.t510 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X763 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0.t15 VGND.t411 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X765 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S uo_out[1].t2 VPWR.t340 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X766 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0.t12 VPWR.t456 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X767 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t38 VPWR.t535 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X768 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t3 VPWR.t466 VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 VGND.t383 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t13 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t6 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R54 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X770 VPWR.t325 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X771 VGND.t427 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA7.CN1.t3 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 VGND.t303 SUNSAR_SAR8B_CV_0.XB2.CKN.t7 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X773 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t34 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X774 VPWR.t493 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA7.CN1.t5 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t24 SUNSAR_SAR8B_CV_0.XA3.ENO.t1 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 VPWR.t584 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA4.CP0.t4 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X777 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t20 VGND.t372 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X778 VPWR.t112 VPWR.t109 VPWR.t111 VPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X779 VGND.t80 VGND.t77 VGND.t79 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X780 VPWR.t115 VPWR.t113 VPWR.t114 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t26 VGND.t374 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X782 VGND.t381 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t8 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R55 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X783 VGND.t238 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 VPWR.t394 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t8 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X786 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X787 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t16 VPWR.t597 VPWR.t596 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X788 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t10 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.D<6>.t11 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X790 VPWR.t578 SUNSAR_SAR8B_CV_0.D<7>.t17 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X791 uo_out[2].t0 SUNSAR_CAPT8B_CV_0.XG12.QN VGND.t231 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X792 VPWR.t211 VPWR.t208 VPWR.t210 VPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X793 VGND.t478 SUNSAR_SAR8B_CV_0.D<7>.t10 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t2 VGND.t477 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t22 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 uo_out[2].t1 SUNSAR_CAPT8B_CV_0.XG12.QN VPWR.t291 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t1 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t42 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X798 VPWR.t7 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.D<3>.t1 SUNSAR_SAR8B_CV_0.XA4.CN1.t9 VGND.t326 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X800 VPWR.t490 SUNSAR_SAR8B_CV_0.XA6.CN1.t12 SUNSAR_SAR8B_CV_0.D<1>.t7 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X802 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t7 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t14 VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND.t266 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 VPWR.t532 SUNSAR_SAR8B_CV_0.EN.t35 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 VGND.t543 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t13 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 VPWR.t588 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t4 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X809 SUNSAR_SAR8B_CV_0.EN.t0 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t6 VGND.t506 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X810 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND.t203 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VPWR.t264 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t0 SUNSAR_SAR8B_CV_0.XA4.CP0.t9 VGND.t532 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X813 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X814 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0].t1 VGND.t24 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.XA3.CN1.t7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t9 VPWR.t398 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X816 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t17 VGND.t547 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X817 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t8 VPWR.t523 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X818 SUNSAR_SAR8B_CV_0.D<3>.t3 SUNSAR_SAR8B_CV_0.XA4.CN1.t11 VGND.t328 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X819 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<7>.t11 VPWR.t575 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VGND.t323 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t4 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X821 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND.t236 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X822 VGND.t104 VGND.t102 VGND.t103 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X823 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR.t296 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X824 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X825 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR.t8 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VPWR.t244 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA6.CN1.t7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t9 VGND.t162 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X828 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t0 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND.t249 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X829 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X830 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X831 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t8 SUNSAR_SAR8B_CV_0.XA0.XA9.B VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X832 VPWR.t465 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t7 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X833 ua[1].t2 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP.t1 VGND.t192 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X834 VPWR.t383 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t9 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t1 VPWR.t382 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X835 VGND.t118 VGND.t116 VGND.t117 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X836 VPWR.t420 SUNSAR_SAR8B_CV_0.XA3.CP0.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t6 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X837 VGND.t320 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA3.CN1.t3 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X838 SUNSAR_SAR8B_CV_0.XA3.CN1.t5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t7 VPWR.t396 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X839 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.ENO.t2 VGND.t316 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.ENO.t8 VPWR.t393 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S uo_out[3].t3 VPWR.t438 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R57 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X842 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X843 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND.t228 VGND.t227 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X844 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t3 VPWR.t453 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X845 VPWR.t119 VPWR.t116 VPWR.t118 VPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XA7.CP0.t7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t9 VGND.t300 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R58 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X847 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t7 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X848 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR.t260 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X849 VPWR.t50 VPWR.t48 VPWR.t49 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X850 VGND.t402 SUNSAR_SAR8B_CV_0.XA6.CP0.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t2 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA7.CP0.t6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t8 VPWR.t360 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X852 SUNSAR_SAR8B_CV_0.XA6.CN1.t3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t5 VGND.t160 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X853 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t18 VGND.t435 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X854 VPWR.t608 VGND.t6 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X855 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND.t234 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t10 VGND.t362 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA11.A VPWR.t294 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X858 VPWR.t610 VGND.t8 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X859 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t12 VPWR.t502 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR.t10 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR.t302 VPWR.t301 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X862 SUNSAR_SAR8B_CV_0.XA1.ENO.t0 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND.t171 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X864 VPWR.t233 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t4 VGND.t504 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t27 VGND.t375 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X867 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<0>.t9 VPWR.t353 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X868 uo_out[5].t0 SUNSAR_CAPT8B_CV_0.XD09.QN VGND.t211 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND.t276 VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t6 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t10 VPWR.t459 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VGND.t291 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA5.CP0.t3 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X872 VPWR.t350 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA5.CP0.t5 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X873 SUNSAR_SAR8B_CV_0.XA7.CP0.t5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t7 VGND.t299 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X874 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND.t241 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X875 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR.t265 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X876 SUNSAR_SAR8B_CV_0.XA7.CP0.t1 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t3 VPWR.t357 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 VPWR.t92 VPWR.t89 VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X878 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP.t17 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X879 VGND.t149 VGND.t146 VGND.t148 VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 VPWR.t399 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t1 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VGND.t315 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t13 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t6 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR.t276 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X883 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t1 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X884 uo_out[4].t0 SUNSAR_CAPT8B_CV_0.XE10.QN VGND.t235 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 VPWR.t198 VPWR.t195 VPWR.t197 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X886 VGND.t232 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X887 VGND.t503 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t3 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VPWR.t324 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.t0 VPWR.t323 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP.t12 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X890 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t16 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 uo_out[4].t1 SUNSAR_CAPT8B_CV_0.XE10.QN VPWR.t295 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X892 VPWR.t18 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t8 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X893 VPWR.t404 SUNSAR_SAR8B_CV_0.XA4.CN1.t12 SUNSAR_SAR8B_CV_0.D<3>.t4 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X894 VPWR.t194 VPWR.t192 VPWR.t193 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X895 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t32 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X896 VPWR.t442 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t6 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t2 VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X897 VGND.t467 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t9 SUNSAR_SAR8B_CV_0.D<6>.t1 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 VGND.t551 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t23 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X899 VPWR.t568 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t12 SUNSAR_SAR8B_CV_0.D<6>.t5 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X901 uo_out[1].t0 SUNSAR_CAPT8B_CV_0.XH13.QN VGND.t219 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X902 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP.t16 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X903 VGND.t251 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X905 VPWR.t300 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R60 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X906 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t26 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X909 VGND.t28 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t11 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t5 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X910 VPWR.t23 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t1 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R61 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X911 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t32 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X912 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND.t254 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X913 VGND.t415 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.D<7>.t1 VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X914 tt_um_TT06_SAR_done_0.x4.MP0.G tt_um_TT06_SAR_done_0.x4.MP0.G VGND.t269 VGND.t268 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X915 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VPWR.t232 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA4.CN1.t7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t9 VGND.t312 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X917 VPWR.t221 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA6.CN1.t5 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R62 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X918 VPWR.t541 SUNSAR_SAR8B_CV_0.EN.t56 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X920 VPWR.t369 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t6 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t3 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t8 VPWR.t381 VPWR.t380 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X923 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<6>.t10 VGND.t336 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X924 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X925 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<6>.t9 VPWR.t414 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X926 VPWR.t544 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t6 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND.t252 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X928 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X929 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND.t259 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X930 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X931 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR.t321 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X932 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X933 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X934 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t3 VPWR.t520 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X935 uio_out[0].t0 tt_um_TT06_SAR_done_0.x3.MP1.G VGND.t173 VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X936 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t2 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VPWR.t281 VPWR.t280 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X937 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t34 VGND.t527 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t52 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X939 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR.t238 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X940 VPWR.t135 VPWR.t133 VPWR.t134 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X941 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t8 SUNSAR_SAR8B_CV_0.XA1.XA9.B VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X942 VGND.t534 SUNSAR_SAR8B_CV_0.XA4.CP0.t14 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t2 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XA4.CN1.t3 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t5 VGND.t310 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X944 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VGND.t181 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X945 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S uo_out[2].t2 VGND.t277 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X946 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S uo_out[2].t3 VPWR.t338 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X947 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t7 VGND.t313 VGND.t143 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X948 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t6 VPWR.t379 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X949 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t16 VPWR.t503 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X950 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR.t269 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X951 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN.t26 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X953 VPWR.t609 VGND.t7 sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X954 VGND.t128 VGND.t126 VGND.t127 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X955 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t7 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t9 VPWR.t586 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.ENO.t3 VGND.t360 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X957 VPWR.t417 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA3.CP0.t4 VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t1 SUNSAR_SAR8B_CV_0.XB1.CKN.t3 VGND.t407 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X959 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR.t243 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND.t214 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X961 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t4 VPWR.t463 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X962 VPWR.t482 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.D<7>.t6 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X963 SUNSAR_SAR8B_CV_0.D<0>.t2 SUNSAR_SAR8B_CV_0.XA7.CN1.t11 VGND.t448 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X964 VPWR.t108 VPWR.t105 VPWR.t107 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X965 VGND.t348 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t11 SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA2.XA11.A VPWR.t314 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X967 VGND.t333 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA6.CP0.t5 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.D<0>.t5 SUNSAR_SAR8B_CV_0.XA7.CN1.t10 VPWR.t516 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 TIE_L SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND.t230 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X970 VPWR.t378 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t8 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X971 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND.t239 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X972 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<0>.t8 VPWR.t352 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X974 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR.t299 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R65 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X975 VPWR.t126 VPWR.t124 VPWR.t125 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X976 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE.t28 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND.t523 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<5>.t8 VPWR.t547 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X978 ua[0].t9 SUNSAR_SAR8B_CV_0.XB2.CKN.t5 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA3.ENO.t0 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND.t247 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X980 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VGND.t20 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0.t11 VGND.t389 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X982 uo_out[3].t0 SUNSAR_CAPT8B_CV_0.XF11.QN VGND.t222 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.D<1>.t9 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X984 VGND.t505 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t5 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X985 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0.t9 VPWR.t454 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X986 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t7 VPWR.t464 VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X987 VGND.t438 SUNSAR_SAR8B_CV_0.XA5.CN1.t9 SUNSAR_SAR8B_CV_0.D<2>.t1 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X988 VPWR.t509 SUNSAR_SAR8B_CV_0.XA5.CN1.t14 SUNSAR_SAR8B_CV_0.D<2>.t6 VPWR.t17 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.D<0>.t0 SUNSAR_SAR8B_CV_0.XA7.CN1.t9 VGND.t447 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 ua[0].t4 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_SAR8B_CV_0.D<0>.t7 SUNSAR_SAR8B_CV_0.XA7.CN1.t12 VPWR.t517 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t10 VGND.t465 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X993 VGND.t355 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t13 SUNSAR_SAR8B_CV_0.D<5>.t3 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X994 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t0 SUNSAR_SAR8B_CV_0.EN.t58 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR.t9 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X995 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t6 VPWR.t355 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t0 SUNSAR_SAR8B_CV_0.EN.t18 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X997 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND.t272 VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X999 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1000 VPWR.t376 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA4.CN1.t5 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1001 VPWR.t475 SUNSAR_SAR8B_CV_0.XB1.CKN.t6 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR.t474 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1002 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VPWR.t317 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 ua[0].t8 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1004 VPWR.t522 SUNSAR_SAR8B_CV_0.EN.t5 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1005 VGND.t395 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t2 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.t1 SUNSAR_SAR8B_CV_0.XB2.CKN.t4 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 VGND.t471 SUNSAR_SAR8B_CV_0.XA3.CN1.t9 SUNSAR_SAR8B_CV_0.D<4>.t2 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R67 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1008 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S uo_out[5].t3 VGND.t296 VGND.t133 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 VPWR.t554 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t3 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND.t226 VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1013 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.ENO.t6 VGND.t317 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1014 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.ENO.t7 VPWR.t392 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R68 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1016 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.CKN.t6 VGND.t302 VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN.t9 VPWR.t524 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1018 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1019 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR.t259 VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1020 VGND.t345 SUNSAR_SAR8B_CV_0.XA3.CP0.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t0 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1021 VGND.t444 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t6 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1022 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN.t50 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t19 VGND.t371 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 VPWR.t486 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t2 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1025 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN.t48 VPWR.t540 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VGND.t168 VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S uo_out[4].t2 VGND.t278 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND.t19 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S uo_out[4].t3 VPWR.t339 VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t29 VGND.t377 VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VPWR.t305 VPWR.t27 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1033 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t30 SUNSAR_SAR8B_CV_0.XA7.ENO.t0 VPWR.t71 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1034 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1035 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND.t154 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1036 VGND.t83 VGND.t81 VGND.t82 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1037 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t9 VGND.t508 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1038 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t0 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t7 VPWR.t562 VPWR.t561 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1039 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR.t215 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1040 VPWR.t69 VPWR.t67 VPWR.t68 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1041 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S uo_out[1].t3 VGND.t279 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1042 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND.t273 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1043 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t11 VGND.t466 VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1044 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t0 SUNSAR_SAR8B_CV_0.DONE.t3 VGND.t410 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1045 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND.t258 VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1046 VPWR.t345 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t6 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t1 VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1047 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t1 SUNSAR_SAR8B_CV_0.DONE.t4 VPWR.t476 VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1048 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR.t320 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1049 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND.t264 VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1050 VGND.t432 SUNSAR_SAR8B_CV_0.DONE.t14 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1051 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t7 VPWR.t545 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1052 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1053 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE.t12 VGND.t509 VGND.t31 sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1054 VPWR.t54 VPWR.t51 VPWR.t53 VPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t11 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t9 1060.4
R70 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t14 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t15 1060.4
R71 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t10 1060.4
R72 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t12 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t13 1060.4
R73 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n1 568.956
R74 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t11 568.956
R75 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t15 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n3 568.956
R76 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t14 568.956
R77 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t8 568.956
R78 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t10 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n6 568.956
R79 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t12 568.956
R80 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t13 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n0 568.956
R81 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n11 292.5
R82 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n17 292.5
R83 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 197.272
R84 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n15 112.829
R85 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n16 111.059
R86 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n8 92.5005
R87 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n12 81.5064
R88 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t2 63.8431
R89 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t1 63.8431
R90 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t4 63.8431
R91 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t3 63.8431
R92 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n14 53.4593
R93 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t7 38.8894
R94 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t5 38.8894
R95 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t6 38.8894
R96 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t0 38.8894
R97 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n10 37.5726
R98 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n13 29.5534
R99 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.5854
R100 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n1 20.3299
R101 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R102 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R103 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n0 20.3299
R104 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n2 20.3299
R105 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R106 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R107 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R108 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n5 20.3299
R109 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n4 20.3299
R110 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R111 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R112 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n0 20.3299
R113 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n7 20.3299
R114 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n9 20.3299
R115 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 20.3299
R116 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n18 20.3299
R117 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 17.6946
R118 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 17.6946
R119 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 10.3476
R120 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.168144
R121 VGND.n1971 VGND.n1970 21703.2
R122 VGND.t143 VGND.n2332 14478.2
R123 VGND.t120 VGND.t49 13996.1
R124 VGND.t64 VGND.t57 13996.1
R125 VGND.t133 VGND.t88 13996.1
R126 VGND.t9 VGND.n1034 12001.4
R127 VGND.n1035 VGND.t428 11148.4
R128 VGND.n1971 VGND.n1034 8907.51
R129 VGND.n2436 VGND.n667 8835.2
R130 VGND.n1972 VGND.n1020 8520.99
R131 VGND.n1020 VGND.t35 7833.63
R132 VGND.n1617 VGND.n1033 6617.6
R133 VGND.n2727 VGND.n2726 6617.6
R134 VGND.n1084 VGND.n1035 5329.03
R135 VGND.t39 VGND.n80 5108.47
R136 VGND.n2726 VGND.n2725 1923.29
R137 VGND.n2726 VGND.n82 1921.57
R138 VGND.n2525 VGND.n159 1401.45
R139 VGND.n2525 VGND.n2524 1396.14
R140 VGND.n1970 VGND.n1033 1198.89
R141 VGND.n1983 VGND.n667 1078.7
R142 VGND.n2509 VGND.n2508 1073.01
R143 VGND.n1972 VGND.n1971 1009.66
R144 VGND.n2437 VGND.n81 957.933
R145 VGND.n1973 VGND.n1972 954.444
R146 VGND.n2605 VGND.n80 924.966
R147 VGND.n2438 VGND.n667 809.029
R148 VGND.n1969 VGND.t9 764.909
R149 VGND.n1969 VGND.t49 764.909
R150 VGND.n1617 VGND.t120 764.909
R151 VGND.n1617 VGND.t64 764.909
R152 VGND.n2436 VGND.t57 764.909
R153 VGND.n2436 VGND.t88 764.909
R154 VGND.n2372 VGND.t133 764.909
R155 VGND.n2372 VGND.t143 764.909
R156 VGND.n1972 VGND.n1033 678.889
R157 VGND.n2507 VGND 672.929
R158 VGND.n2435 VGND 663.399
R159 VGND.n1616 VGND 663.399
R160 VGND VGND.n1085 663.399
R161 VGND.n2443 VGND.n542 661.385
R162 VGND.n665 VGND.n664 660.793
R163 VGND.n2499 VGND.n2498 660.793
R164 VGND.n2197 VGND.n50 660.793
R165 VGND.n1274 VGND.n668 660.793
R166 VGND.n1903 VGND.n1444 660.793
R167 VGND VGND.n2501 658.184
R168 VGND VGND.n581 658.184
R169 VGND.n573 VGND 658.184
R170 VGND.n2500 VGND.t35 620.771
R171 VGND.n2438 VGND.t262 620.771
R172 VGND.n2438 VGND.t192 620.771
R173 VGND.n666 VGND.t39 620.771
R174 VGND.n2371 VGND 592.822
R175 VGND.n2331 VGND 592.822
R176 VGND.n1032 VGND.n1031 590.216
R177 VGND.n2724 VGND.n2723 590.216
R178 VGND.n1071 VGND.n1044 590.216
R179 VGND VGND.n708 587.607
R180 VGND VGND.n698 587.607
R181 VGND VGND.n1618 587.607
R182 VGND.n1019 VGND 587.607
R183 VGND VGND.n2373 587.607
R184 VGND VGND.n788 587.607
R185 VGND VGND.n2728 587.607
R186 VGND.n2604 VGND 587.607
R187 VGND VGND.n1038 587.607
R188 VGND.n1276 VGND.n1275 585
R189 VGND.n1278 VGND.n1277 585
R190 VGND.n1280 VGND.n1279 585
R191 VGND.n1282 VGND.n1281 585
R192 VGND.n1284 VGND.n1283 585
R193 VGND.n1286 VGND.n1285 585
R194 VGND.n1288 VGND.n1287 585
R195 VGND.n1290 VGND.n1289 585
R196 VGND.n1292 VGND.n1291 585
R197 VGND.n1294 VGND.n1293 585
R198 VGND.n1296 VGND.n1295 585
R199 VGND.n1298 VGND.n1297 585
R200 VGND.n1300 VGND.n1299 585
R201 VGND.n1302 VGND.n1301 585
R202 VGND.n1304 VGND.n1303 585
R203 VGND.n1306 VGND.n1305 585
R204 VGND.n1308 VGND.n1307 585
R205 VGND.n1310 VGND.n1309 585
R206 VGND.n1312 VGND.n1311 585
R207 VGND.n1314 VGND.n1313 585
R208 VGND.n1316 VGND.n1315 585
R209 VGND.n1318 VGND.n1317 585
R210 VGND.n1320 VGND.n1319 585
R211 VGND.n1322 VGND.n1321 585
R212 VGND.n1324 VGND.n1323 585
R213 VGND.n1326 VGND.n1325 585
R214 VGND.n1328 VGND.n1327 585
R215 VGND.n1330 VGND.n1329 585
R216 VGND.n1332 VGND.n1331 585
R217 VGND.n1334 VGND.n1333 585
R218 VGND.n1336 VGND.n1335 585
R219 VGND.n1338 VGND.n1337 585
R220 VGND.n1340 VGND.n1339 585
R221 VGND.n1342 VGND.n1341 585
R222 VGND.n1344 VGND.n1343 585
R223 VGND.n1346 VGND.n1345 585
R224 VGND.n1348 VGND.n1347 585
R225 VGND.n1350 VGND.n1349 585
R226 VGND.n1352 VGND.n1351 585
R227 VGND.n1354 VGND.n1353 585
R228 VGND.n1356 VGND.n1355 585
R229 VGND.n1358 VGND.n1357 585
R230 VGND.n1360 VGND.n1359 585
R231 VGND.n1362 VGND.n1361 585
R232 VGND.n1364 VGND.n1363 585
R233 VGND.n1366 VGND.n1365 585
R234 VGND.n1368 VGND.n1367 585
R235 VGND.n1370 VGND.n1369 585
R236 VGND.n1372 VGND.n1371 585
R237 VGND.n1374 VGND.n1373 585
R238 VGND.n1376 VGND.n1375 585
R239 VGND.n1378 VGND.n1377 585
R240 VGND.n1380 VGND.n1379 585
R241 VGND.n1382 VGND.n1381 585
R242 VGND.n1384 VGND.n1383 585
R243 VGND.n1386 VGND.n1385 585
R244 VGND.n1388 VGND.n1387 585
R245 VGND.n1390 VGND.n1389 585
R246 VGND.n1392 VGND.n1391 585
R247 VGND.n2437 VGND.n698 585
R248 VGND.n1902 VGND.n1901 585
R249 VGND.n1900 VGND.n1445 585
R250 VGND.n1898 VGND.n1897 585
R251 VGND.n1896 VGND.n1446 585
R252 VGND.n1895 VGND.n1894 585
R253 VGND.n1892 VGND.n1891 585
R254 VGND.n1890 VGND.n1889 585
R255 VGND.n1888 VGND.n1887 585
R256 VGND.n1886 VGND.n1885 585
R257 VGND.n1884 VGND.n1883 585
R258 VGND.n1882 VGND.n1881 585
R259 VGND.n1880 VGND.n1450 585
R260 VGND.n1878 VGND.n1877 585
R261 VGND.n1876 VGND.n1451 585
R262 VGND.n1875 VGND.n1874 585
R263 VGND.n1872 VGND.n1452 585
R264 VGND.n1870 VGND.n1869 585
R265 VGND.n1868 VGND.n1453 585
R266 VGND.n1867 VGND.n1866 585
R267 VGND.n1864 VGND.n1863 585
R268 VGND.n1862 VGND.n1861 585
R269 VGND.n1860 VGND.n1859 585
R270 VGND.n1858 VGND.n1857 585
R271 VGND.n1856 VGND.n1855 585
R272 VGND.n1854 VGND.n1853 585
R273 VGND.n1852 VGND.n1457 585
R274 VGND.n1850 VGND.n1849 585
R275 VGND.n1848 VGND.n1458 585
R276 VGND.n1847 VGND.n1846 585
R277 VGND.n1844 VGND.n1843 585
R278 VGND.n1842 VGND.n1841 585
R279 VGND.n1840 VGND.n1839 585
R280 VGND.n1838 VGND.n1837 585
R281 VGND.n1836 VGND.n1835 585
R282 VGND.n1834 VGND.n1833 585
R283 VGND.n1832 VGND.n1462 585
R284 VGND.n1830 VGND.n1829 585
R285 VGND.n1828 VGND.n1463 585
R286 VGND.n1827 VGND.n1826 585
R287 VGND.n1824 VGND.n1823 585
R288 VGND.n1822 VGND.n1821 585
R289 VGND.n1820 VGND.n1819 585
R290 VGND.n1818 VGND.n1817 585
R291 VGND.n1816 VGND.n1815 585
R292 VGND.n1814 VGND.n1813 585
R293 VGND.n1812 VGND.n1811 585
R294 VGND.n1810 VGND.n1809 585
R295 VGND.n1808 VGND.n1807 585
R296 VGND.n1806 VGND.n1805 585
R297 VGND.n1804 VGND.n1803 585
R298 VGND.n1802 VGND.n1801 585
R299 VGND.n1800 VGND.n1799 585
R300 VGND.n1798 VGND.n1797 585
R301 VGND.n1796 VGND.n1795 585
R302 VGND.n1794 VGND.n1793 585
R303 VGND.n1792 VGND.n1791 585
R304 VGND.n1790 VGND.n1789 585
R305 VGND.n1788 VGND.n1787 585
R306 VGND.n1786 VGND.n1785 585
R307 VGND.n1784 VGND.n1783 585
R308 VGND.n1784 VGND.n667 585
R309 VGND.n1973 VGND.n1032 585
R310 VGND.n1977 VGND.n1976 585
R311 VGND.n1976 VGND.n1975 585
R312 VGND.n1978 VGND.n1021 585
R313 VGND.n1974 VGND.n1021 585
R314 VGND.n1981 VGND.n1980 585
R315 VGND.n1982 VGND.n1981 585
R316 VGND.n1979 VGND.n1022 585
R317 VGND.n887 VGND.n885 585
R318 VGND.n1986 VGND.n1985 585
R319 VGND.n888 VGND.n886 585
R320 VGND.n917 VGND.n916 585
R321 VGND.n919 VGND.n918 585
R322 VGND.n921 VGND.n920 585
R323 VGND.n923 VGND.n922 585
R324 VGND.n925 VGND.n924 585
R325 VGND.n927 VGND.n926 585
R326 VGND.n929 VGND.n928 585
R327 VGND.n931 VGND.n930 585
R328 VGND.n933 VGND.n932 585
R329 VGND.n935 VGND.n934 585
R330 VGND.n937 VGND.n936 585
R331 VGND.n939 VGND.n938 585
R332 VGND.n941 VGND.n940 585
R333 VGND.n943 VGND.n942 585
R334 VGND.n945 VGND.n944 585
R335 VGND.n947 VGND.n946 585
R336 VGND.n949 VGND.n948 585
R337 VGND.n951 VGND.n950 585
R338 VGND.n953 VGND.n952 585
R339 VGND.n955 VGND.n954 585
R340 VGND.n957 VGND.n956 585
R341 VGND.n959 VGND.n958 585
R342 VGND.n961 VGND.n960 585
R343 VGND.n963 VGND.n962 585
R344 VGND.n965 VGND.n964 585
R345 VGND.n967 VGND.n966 585
R346 VGND.n969 VGND.n968 585
R347 VGND.n971 VGND.n970 585
R348 VGND.n973 VGND.n972 585
R349 VGND.n975 VGND.n974 585
R350 VGND.n977 VGND.n976 585
R351 VGND.n979 VGND.n978 585
R352 VGND.n981 VGND.n980 585
R353 VGND.n983 VGND.n982 585
R354 VGND.n985 VGND.n984 585
R355 VGND.n987 VGND.n986 585
R356 VGND.n989 VGND.n988 585
R357 VGND.n991 VGND.n990 585
R358 VGND.n993 VGND.n992 585
R359 VGND.n995 VGND.n994 585
R360 VGND.n997 VGND.n996 585
R361 VGND.n999 VGND.n998 585
R362 VGND.n1001 VGND.n1000 585
R363 VGND.n1003 VGND.n1002 585
R364 VGND.n1005 VGND.n1004 585
R365 VGND.n1007 VGND.n1006 585
R366 VGND.n1009 VGND.n1008 585
R367 VGND.n1011 VGND.n1010 585
R368 VGND.n1013 VGND.n1012 585
R369 VGND.n1014 VGND.n915 585
R370 VGND.n1016 VGND.n1015 585
R371 VGND.n1018 VGND.n882 585
R372 VGND.n1983 VGND.n1019 585
R373 VGND.n1098 VGND.n1097 585
R374 VGND.n1967 VGND.n1966 585
R375 VGND.n1965 VGND.n1096 585
R376 VGND.n1964 VGND.n1963 585
R377 VGND.n1962 VGND.n1961 585
R378 VGND.n1960 VGND.n1959 585
R379 VGND.n1958 VGND.n1957 585
R380 VGND.n1956 VGND.n1955 585
R381 VGND.n1954 VGND.n1953 585
R382 VGND.n1952 VGND.n1951 585
R383 VGND.n1950 VGND.n1949 585
R384 VGND.n1948 VGND.n1947 585
R385 VGND.n1946 VGND.n1945 585
R386 VGND.n1944 VGND.n1943 585
R387 VGND.n1942 VGND.n1941 585
R388 VGND.n1940 VGND.n1939 585
R389 VGND.n1938 VGND.n1937 585
R390 VGND.n1936 VGND.n1935 585
R391 VGND.n1934 VGND.n1933 585
R392 VGND.n1932 VGND.n1931 585
R393 VGND.n1930 VGND.n1929 585
R394 VGND.n1928 VGND.n1086 585
R395 VGND.n1969 VGND.n1086 585
R396 VGND.n1615 VGND.n1579 585
R397 VGND.n1614 VGND.n1578 585
R398 VGND.n1617 VGND.n1578 585
R399 VGND.n1613 VGND.n1612 585
R400 VGND.n1611 VGND.n1610 585
R401 VGND.n1609 VGND.n1608 585
R402 VGND.n1607 VGND.n1606 585
R403 VGND.n1605 VGND.n1604 585
R404 VGND.n1603 VGND.n1602 585
R405 VGND.n1601 VGND.n1600 585
R406 VGND.n1599 VGND.n1598 585
R407 VGND.n1597 VGND.n1596 585
R408 VGND.n1595 VGND.n1594 585
R409 VGND.n1593 VGND.n1592 585
R410 VGND.n1591 VGND.n1590 585
R411 VGND.n1589 VGND.n1588 585
R412 VGND.n1587 VGND.n1586 585
R413 VGND.n1585 VGND.n1584 585
R414 VGND.n1583 VGND.n1582 585
R415 VGND.n1581 VGND.n1580 585
R416 VGND.n1568 VGND.n1567 585
R417 VGND.n1618 VGND.n1617 585
R418 VGND.n2434 VGND.n710 585
R419 VGND.n2433 VGND.n709 585
R420 VGND.n2436 VGND.n709 585
R421 VGND.n2432 VGND.n2431 585
R422 VGND.n2430 VGND.n2429 585
R423 VGND.n2428 VGND.n2427 585
R424 VGND.n2426 VGND.n2425 585
R425 VGND.n2424 VGND.n2423 585
R426 VGND.n2422 VGND.n2421 585
R427 VGND.n2420 VGND.n2419 585
R428 VGND.n2418 VGND.n2417 585
R429 VGND.n2416 VGND.n2415 585
R430 VGND.n2414 VGND.n2413 585
R431 VGND.n2412 VGND.n2411 585
R432 VGND.n2410 VGND.n2409 585
R433 VGND.n2408 VGND.n2407 585
R434 VGND.n2406 VGND.n2405 585
R435 VGND.n2404 VGND.n2403 585
R436 VGND.n2402 VGND.n2401 585
R437 VGND.n2400 VGND.n2399 585
R438 VGND.n2398 VGND.n2397 585
R439 VGND.n2436 VGND.n708 585
R440 VGND.n2372 VGND.n2371 585
R441 VGND.n2370 VGND.n2333 585
R442 VGND.n2369 VGND.n2368 585
R443 VGND.n2367 VGND.n2366 585
R444 VGND.n2365 VGND.n2364 585
R445 VGND.n2363 VGND.n2362 585
R446 VGND.n2361 VGND.n2360 585
R447 VGND.n2359 VGND.n2358 585
R448 VGND.n2357 VGND.n2356 585
R449 VGND.n2355 VGND.n2354 585
R450 VGND.n2353 VGND.n2352 585
R451 VGND.n2351 VGND.n2350 585
R452 VGND.n2349 VGND.n2348 585
R453 VGND.n2347 VGND.n2346 585
R454 VGND.n2345 VGND.n2344 585
R455 VGND.n2343 VGND.n2342 585
R456 VGND.n2341 VGND.n2340 585
R457 VGND.n2339 VGND.n2338 585
R458 VGND.n2337 VGND.n2336 585
R459 VGND.n2335 VGND.n2334 585
R460 VGND.n758 VGND.n757 585
R461 VGND.n2373 VGND.n2372 585
R462 VGND.n2196 VGND.n2195 585
R463 VGND.n2194 VGND.n2193 585
R464 VGND.n2192 VGND.n2191 585
R465 VGND.n2190 VGND.n2189 585
R466 VGND.n2188 VGND.n2187 585
R467 VGND.n2186 VGND.n2185 585
R468 VGND.n2184 VGND.n2183 585
R469 VGND.n2182 VGND.n2181 585
R470 VGND.n2180 VGND.n2179 585
R471 VGND.n2178 VGND.n2177 585
R472 VGND.n2176 VGND.n2175 585
R473 VGND.n2174 VGND.n2173 585
R474 VGND.n2172 VGND.n2171 585
R475 VGND.n2170 VGND.n2169 585
R476 VGND.n2168 VGND.n2167 585
R477 VGND.n2166 VGND.n2165 585
R478 VGND.n2164 VGND.n2163 585
R479 VGND.n2162 VGND.n2161 585
R480 VGND.n2160 VGND.n2159 585
R481 VGND.n2158 VGND.n2157 585
R482 VGND.n2156 VGND.n2155 585
R483 VGND.n2154 VGND.n2153 585
R484 VGND.n2152 VGND.n2151 585
R485 VGND.n2150 VGND.n2149 585
R486 VGND.n2148 VGND.n2147 585
R487 VGND.n2146 VGND.n2145 585
R488 VGND.n2144 VGND.n2143 585
R489 VGND.n2142 VGND.n2141 585
R490 VGND.n2140 VGND.n2139 585
R491 VGND.n2138 VGND.n2137 585
R492 VGND.n2136 VGND.n2135 585
R493 VGND.n2134 VGND.n2133 585
R494 VGND.n2132 VGND.n2131 585
R495 VGND.n2130 VGND.n2129 585
R496 VGND.n2128 VGND.n2127 585
R497 VGND.n2126 VGND.n2125 585
R498 VGND.n2124 VGND.n2123 585
R499 VGND.n2122 VGND.n2121 585
R500 VGND.n2120 VGND.n2119 585
R501 VGND.n2118 VGND.n2117 585
R502 VGND.n2116 VGND.n2115 585
R503 VGND.n2114 VGND.n2113 585
R504 VGND.n2112 VGND.n2111 585
R505 VGND.n2110 VGND.n2109 585
R506 VGND.n2108 VGND.n2107 585
R507 VGND.n2106 VGND.n2105 585
R508 VGND.n2104 VGND.n2103 585
R509 VGND.n2102 VGND.n2101 585
R510 VGND.n2100 VGND.n2099 585
R511 VGND.n2098 VGND.n2097 585
R512 VGND.n2096 VGND.n2095 585
R513 VGND.n2094 VGND.n2093 585
R514 VGND.n2092 VGND.n2091 585
R515 VGND.n2090 VGND.n2089 585
R516 VGND.n2088 VGND.n2087 585
R517 VGND.n2086 VGND.n2085 585
R518 VGND.n2084 VGND.n2083 585
R519 VGND.n2082 VGND.n2081 585
R520 VGND.n49 VGND.n48 585
R521 VGND.n2728 VGND.n2727 585
R522 VGND.n2332 VGND.n2331 585
R523 VGND.n2330 VGND.n769 585
R524 VGND.n771 VGND.n769 585
R525 VGND.n2329 VGND.n2328 585
R526 VGND.n2328 VGND.n2327 585
R527 VGND.n774 VGND.n770 585
R528 VGND.n2326 VGND.n770 585
R529 VGND.n2324 VGND.n2323 585
R530 VGND.n2325 VGND.n2324 585
R531 VGND.n2322 VGND.n773 585
R532 VGND.n773 VGND.n772 585
R533 VGND.n2321 VGND.n2320 585
R534 VGND.n2320 VGND.n2319 585
R535 VGND.n777 VGND.n775 585
R536 VGND.n2318 VGND.n775 585
R537 VGND.n2316 VGND.n2315 585
R538 VGND.n2317 VGND.n2316 585
R539 VGND.n2314 VGND.n776 585
R540 VGND.n779 VGND.n776 585
R541 VGND.n2313 VGND.n2312 585
R542 VGND.n2312 VGND.n2311 585
R543 VGND.n782 VGND.n778 585
R544 VGND.n2310 VGND.n778 585
R545 VGND.n2308 VGND.n2307 585
R546 VGND.n2309 VGND.n2308 585
R547 VGND.n2306 VGND.n781 585
R548 VGND.n781 VGND.n780 585
R549 VGND.n2305 VGND.n2304 585
R550 VGND.n2304 VGND.n2303 585
R551 VGND.n785 VGND.n783 585
R552 VGND.n2302 VGND.n783 585
R553 VGND.n2300 VGND.n2299 585
R554 VGND.n2301 VGND.n2300 585
R555 VGND.n2298 VGND.n784 585
R556 VGND.n787 VGND.n784 585
R557 VGND.n2297 VGND.n2296 585
R558 VGND.n2296 VGND.n2295 585
R559 VGND.n789 VGND.n786 585
R560 VGND.n2294 VGND.n786 585
R561 VGND.n2292 VGND.n2291 585
R562 VGND.n2293 VGND.n2292 585
R563 VGND.n788 VGND.n82 585
R564 VGND.n2725 VGND.n2724 585
R565 VGND.n2722 VGND.n83 585
R566 VGND.n85 VGND.n83 585
R567 VGND.n2721 VGND.n2720 585
R568 VGND.n2720 VGND.n2719 585
R569 VGND.n87 VGND.n84 585
R570 VGND.n2718 VGND.n84 585
R571 VGND.n2716 VGND.n2715 585
R572 VGND.n2717 VGND.n2716 585
R573 VGND.n2714 VGND.n86 585
R574 VGND.n90 VGND.n86 585
R575 VGND.n2713 VGND.n2712 585
R576 VGND.n2712 VGND.n2711 585
R577 VGND.n89 VGND.n88 585
R578 VGND.n2710 VGND.n89 585
R579 VGND.n2708 VGND.n2707 585
R580 VGND.n2709 VGND.n2708 585
R581 VGND.n2706 VGND.n92 585
R582 VGND.n92 VGND.n91 585
R583 VGND.n2705 VGND.n2704 585
R584 VGND.n2704 VGND.n2703 585
R585 VGND.n95 VGND.n93 585
R586 VGND.n2702 VGND.n93 585
R587 VGND.n2700 VGND.n2699 585
R588 VGND.n2701 VGND.n2700 585
R589 VGND.n2698 VGND.n94 585
R590 VGND.n97 VGND.n94 585
R591 VGND.n2697 VGND.n2696 585
R592 VGND.n2696 VGND.n2695 585
R593 VGND.n99 VGND.n96 585
R594 VGND.n2694 VGND.n96 585
R595 VGND.n2692 VGND.n2691 585
R596 VGND.n2693 VGND.n2692 585
R597 VGND.n2690 VGND.n98 585
R598 VGND.n101 VGND.n98 585
R599 VGND.n2689 VGND.n2688 585
R600 VGND.n2688 VGND.n2687 585
R601 VGND.n104 VGND.n100 585
R602 VGND.n2686 VGND.n100 585
R603 VGND.n2684 VGND.n2683 585
R604 VGND.n2685 VGND.n2684 585
R605 VGND.n2682 VGND.n103 585
R606 VGND.n103 VGND.n102 585
R607 VGND.n2681 VGND.n2680 585
R608 VGND.n2680 VGND.n2679 585
R609 VGND.n107 VGND.n105 585
R610 VGND.n2678 VGND.n105 585
R611 VGND.n2676 VGND.n2675 585
R612 VGND.n2677 VGND.n2676 585
R613 VGND.n2674 VGND.n106 585
R614 VGND.n109 VGND.n106 585
R615 VGND.n2673 VGND.n2672 585
R616 VGND.n2672 VGND.n2671 585
R617 VGND.n111 VGND.n108 585
R618 VGND.n2670 VGND.n108 585
R619 VGND.n2668 VGND.n2667 585
R620 VGND.n2669 VGND.n2668 585
R621 VGND.n2666 VGND.n110 585
R622 VGND.n114 VGND.n110 585
R623 VGND.n2665 VGND.n2664 585
R624 VGND.n2664 VGND.n2663 585
R625 VGND.n113 VGND.n112 585
R626 VGND.n2662 VGND.n113 585
R627 VGND.n2660 VGND.n2659 585
R628 VGND.n2661 VGND.n2660 585
R629 VGND.n2658 VGND.n115 585
R630 VGND.n117 VGND.n115 585
R631 VGND.n2657 VGND.n2656 585
R632 VGND.n2656 VGND.n2655 585
R633 VGND.n119 VGND.n116 585
R634 VGND.n2654 VGND.n116 585
R635 VGND.n2652 VGND.n2651 585
R636 VGND.n2653 VGND.n2652 585
R637 VGND.n2650 VGND.n118 585
R638 VGND.n121 VGND.n118 585
R639 VGND.n2649 VGND.n2648 585
R640 VGND.n2648 VGND.n2647 585
R641 VGND.n124 VGND.n120 585
R642 VGND.n2646 VGND.n120 585
R643 VGND.n2644 VGND.n2643 585
R644 VGND.n2645 VGND.n2644 585
R645 VGND.n2642 VGND.n123 585
R646 VGND.n123 VGND.n122 585
R647 VGND.n2641 VGND.n2640 585
R648 VGND.n2640 VGND.n2639 585
R649 VGND.n128 VGND.n125 585
R650 VGND.n2638 VGND.n125 585
R651 VGND.n2636 VGND.n2635 585
R652 VGND.n2637 VGND.n2636 585
R653 VGND.n2634 VGND.n127 585
R654 VGND.n127 VGND.n126 585
R655 VGND.n2633 VGND.n2632 585
R656 VGND.n2632 VGND.n2631 585
R657 VGND.n132 VGND.n129 585
R658 VGND.n2630 VGND.n129 585
R659 VGND.n2628 VGND.n2627 585
R660 VGND.n2629 VGND.n2628 585
R661 VGND.n2626 VGND.n131 585
R662 VGND.n131 VGND.n130 585
R663 VGND.n2625 VGND.n2624 585
R664 VGND.n2624 VGND.n2623 585
R665 VGND.n134 VGND.n133 585
R666 VGND.n2622 VGND.n134 585
R667 VGND.n2620 VGND.n2619 585
R668 VGND.n2621 VGND.n2620 585
R669 VGND.n2618 VGND.n136 585
R670 VGND.n136 VGND.n135 585
R671 VGND.n2617 VGND.n2616 585
R672 VGND.n2616 VGND.n2615 585
R673 VGND.n138 VGND.n137 585
R674 VGND.n2614 VGND.n138 585
R675 VGND.n2612 VGND.n2611 585
R676 VGND.n2613 VGND.n2612 585
R677 VGND.n2610 VGND.n140 585
R678 VGND.n140 VGND.n139 585
R679 VGND.n2609 VGND.n2608 585
R680 VGND.n2608 VGND.n2607 585
R681 VGND.n142 VGND.n141 585
R682 VGND.n2606 VGND.n142 585
R683 VGND.n2605 VGND.n2604 585
R684 VGND.n2442 VGND.n2441 585
R685 VGND.n2440 VGND.n543 585
R686 VGND.n551 VGND.n544 585
R687 VGND.n553 VGND.n552 585
R688 VGND.n555 VGND.n554 585
R689 VGND.n557 VGND.n556 585
R690 VGND.n559 VGND.n558 585
R691 VGND.n561 VGND.n560 585
R692 VGND.n563 VGND.n562 585
R693 VGND.n565 VGND.n564 585
R694 VGND.n567 VGND.n566 585
R695 VGND.n569 VGND.n568 585
R696 VGND.n570 VGND.n550 585
R697 VGND.n572 VGND.n571 585
R698 VGND.n2496 VGND.n540 585
R699 VGND.n2495 VGND.n539 585
R700 VGND.n2500 VGND.n539 585
R701 VGND.n2494 VGND.n2493 585
R702 VGND.n2492 VGND.n2491 585
R703 VGND.n2490 VGND.n2489 585
R704 VGND.n2488 VGND.n2487 585
R705 VGND.n2486 VGND.n2485 585
R706 VGND.n2484 VGND.n2483 585
R707 VGND.n2482 VGND.n2481 585
R708 VGND.n2480 VGND.n2479 585
R709 VGND.n2478 VGND.n2477 585
R710 VGND.n2476 VGND.n2475 585
R711 VGND.n2474 VGND.n2473 585
R712 VGND.n2472 VGND.n2471 585
R713 VGND.n2470 VGND.n2469 585
R714 VGND.n2468 VGND.n2467 585
R715 VGND.n531 VGND.n530 585
R716 VGND.n600 VGND.n583 585
R717 VGND.n601 VGND.n582 585
R718 VGND.n666 VGND.n582 585
R719 VGND.n603 VGND.n602 585
R720 VGND.n614 VGND.n613 585
R721 VGND.n616 VGND.n615 585
R722 VGND.n618 VGND.n617 585
R723 VGND.n620 VGND.n619 585
R724 VGND.n622 VGND.n621 585
R725 VGND.n624 VGND.n623 585
R726 VGND.n626 VGND.n625 585
R727 VGND.n628 VGND.n627 585
R728 VGND.n630 VGND.n629 585
R729 VGND.n632 VGND.n631 585
R730 VGND.n634 VGND.n633 585
R731 VGND.n636 VGND.n635 585
R732 VGND.n638 VGND.n637 585
R733 VGND.n640 VGND.n639 585
R734 VGND.n1044 VGND.n1043 585
R735 VGND.n1072 VGND.n1042 585
R736 VGND.n1042 VGND.n1041 585
R737 VGND.n1074 VGND.n1073 585
R738 VGND.n1075 VGND.n1074 585
R739 VGND.n1040 VGND.n1039 585
R740 VGND.n1076 VGND.n1040 585
R741 VGND.n1079 VGND.n1078 585
R742 VGND.n1078 VGND.n1077 585
R743 VGND.n1080 VGND.n1037 585
R744 VGND.n1037 VGND.n1036 585
R745 VGND.n1082 VGND.n1081 585
R746 VGND.n1083 VGND.n1082 585
R747 VGND.n1038 VGND.n1035 585
R748 VGND.n1070 VGND.t109 568.956
R749 VGND.n663 VGND.t126 568.956
R750 VGND.n642 VGND.t102 568.956
R751 VGND.n611 VGND.t38 568.956
R752 VGND.n2465 VGND.t34 568.956
R753 VGND.n2445 VGND.t42 568.956
R754 VGND.n2503 VGND.t45 568.956
R755 VGND.n2602 VGND.t105 568.956
R756 VGND.n2080 VGND.t113 568.956
R757 VGND.n2198 VGND.t81 568.956
R758 VGND.n47 VGND.t67 568.956
R759 VGND.n2375 VGND.t132 568.956
R760 VGND.n756 VGND.t142 568.956
R761 VGND.n1927 VGND.t48 568.956
R762 VGND.n1146 VGND.t116 568.956
R763 VGND.n2029 VGND.t136 568.956
R764 VGND.n1273 VGND.t95 568.956
R765 VGND.n1202 VGND.t60 568.956
R766 VGND.n1394 VGND.t30 568.956
R767 VGND.n2395 VGND.t87 568.956
R768 VGND.n1676 VGND.t56 568.956
R769 VGND.n1238 VGND.t129 568.956
R770 VGND.n1782 VGND.t74 568.956
R771 VGND.n1538 VGND.t91 568.956
R772 VGND.n1443 VGND.t99 568.956
R773 VGND.n1645 VGND.t63 568.956
R774 VGND.n1647 VGND.t119 568.956
R775 VGND.n1904 VGND.t123 568.956
R776 VGND.n1030 VGND.t52 568.956
R777 VGND.n2031 VGND.t77 568.956
R778 VGND.n1988 VGND.t84 568.956
R779 VGND.n2730 VGND.t139 568.956
R780 VGND.n2289 VGND.t146 568.956
R781 VGND.n2534 VGND.t70 568.956
R782 VGND.n2727 VGND.n80 531.433
R783 VGND.n1983 VGND.n1020 496.974
R784 VGND.n2500 VGND.t262 413.848
R785 VGND.t192 VGND.n666 413.848
R786 VGND.n527 VGND.n526 389.514
R787 VGND.n1983 VGND.t11 375.652
R788 VGND.n1983 VGND.t78 375.652
R789 VGND.n2437 VGND.t96 345.601
R790 VGND.n2437 VGND.t31 345.601
R791 VGND.n667 VGND.t92 345.601
R792 VGND.n667 VGND.t22 345.601
R793 VGND.n2727 VGND.t16 345.601
R794 VGND.n2727 VGND.t25 345.601
R795 VGND.n2497 VGND.n2443 316.988
R796 VGND.n2443 VGND.n541 316.988
R797 VGND.n2508 VGND.n2507 315.18
R798 VGND.n1043 VGND.n1034 289.387
R799 VGND.n2438 VGND.n2437 269.676
R800 VGND.n2437 VGND.n668 257.212
R801 VGND.n2437 VGND.n669 257.212
R802 VGND.n2437 VGND.n670 257.212
R803 VGND.n2437 VGND.n671 257.212
R804 VGND.n2437 VGND.n672 257.212
R805 VGND.n2437 VGND.n673 257.212
R806 VGND.n2437 VGND.n674 257.212
R807 VGND.n2437 VGND.n675 257.212
R808 VGND.n2437 VGND.n676 257.212
R809 VGND.n2437 VGND.n677 257.212
R810 VGND.n2437 VGND.n678 257.212
R811 VGND.n2437 VGND.n679 257.212
R812 VGND.n2437 VGND.n680 257.212
R813 VGND.n2437 VGND.n681 257.212
R814 VGND.n2437 VGND.n682 257.212
R815 VGND.n2437 VGND.n683 257.212
R816 VGND.n2437 VGND.n684 257.212
R817 VGND.n2437 VGND.n685 257.212
R818 VGND.n2437 VGND.n686 257.212
R819 VGND.n2437 VGND.n687 257.212
R820 VGND.n2437 VGND.n688 257.212
R821 VGND.n2437 VGND.n689 257.212
R822 VGND.n2437 VGND.n690 257.212
R823 VGND.n2437 VGND.n691 257.212
R824 VGND.n2437 VGND.n692 257.212
R825 VGND.n2437 VGND.n693 257.212
R826 VGND.n2437 VGND.n694 257.212
R827 VGND.n2437 VGND.n695 257.212
R828 VGND.n2437 VGND.n696 257.212
R829 VGND.n2437 VGND.n697 257.212
R830 VGND.n1444 VGND.n667 257.212
R831 VGND.n1899 VGND.n667 257.212
R832 VGND.n1893 VGND.n667 257.212
R833 VGND.n1447 VGND.n667 257.212
R834 VGND.n1448 VGND.n667 257.212
R835 VGND.n1449 VGND.n667 257.212
R836 VGND.n1879 VGND.n667 257.212
R837 VGND.n1873 VGND.n667 257.212
R838 VGND.n1871 VGND.n667 257.212
R839 VGND.n1865 VGND.n667 257.212
R840 VGND.n1454 VGND.n667 257.212
R841 VGND.n1455 VGND.n667 257.212
R842 VGND.n1456 VGND.n667 257.212
R843 VGND.n1851 VGND.n667 257.212
R844 VGND.n1845 VGND.n667 257.212
R845 VGND.n1459 VGND.n667 257.212
R846 VGND.n1460 VGND.n667 257.212
R847 VGND.n1461 VGND.n667 257.212
R848 VGND.n1831 VGND.n667 257.212
R849 VGND.n1825 VGND.n667 257.212
R850 VGND.n1464 VGND.n667 257.212
R851 VGND.n1465 VGND.n667 257.212
R852 VGND.n1466 VGND.n667 257.212
R853 VGND.n1467 VGND.n667 257.212
R854 VGND.n1468 VGND.n667 257.212
R855 VGND.n1469 VGND.n667 257.212
R856 VGND.n1470 VGND.n667 257.212
R857 VGND.n1471 VGND.n667 257.212
R858 VGND.n1472 VGND.n667 257.212
R859 VGND.n1473 VGND.n667 257.212
R860 VGND.n1983 VGND.n889 257.212
R861 VGND.n1984 VGND.n1983 257.212
R862 VGND.n1983 VGND.n890 257.212
R863 VGND.n1983 VGND.n891 257.212
R864 VGND.n1983 VGND.n892 257.212
R865 VGND.n1983 VGND.n893 257.212
R866 VGND.n1983 VGND.n894 257.212
R867 VGND.n1983 VGND.n895 257.212
R868 VGND.n1983 VGND.n896 257.212
R869 VGND.n1983 VGND.n897 257.212
R870 VGND.n1983 VGND.n898 257.212
R871 VGND.n1983 VGND.n899 257.212
R872 VGND.n1983 VGND.n900 257.212
R873 VGND.n1983 VGND.n901 257.212
R874 VGND.n1983 VGND.n902 257.212
R875 VGND.n1983 VGND.n903 257.212
R876 VGND.n1983 VGND.n904 257.212
R877 VGND.n1983 VGND.n905 257.212
R878 VGND.n1983 VGND.n906 257.212
R879 VGND.n1983 VGND.n907 257.212
R880 VGND.n1983 VGND.n908 257.212
R881 VGND.n1983 VGND.n909 257.212
R882 VGND.n1983 VGND.n910 257.212
R883 VGND.n1983 VGND.n911 257.212
R884 VGND.n1983 VGND.n912 257.212
R885 VGND.n1983 VGND.n913 257.212
R886 VGND.n1983 VGND.n914 257.212
R887 VGND.n1983 VGND.n1017 257.212
R888 VGND.n1969 VGND.n1085 257.212
R889 VGND.n1969 VGND.n1968 257.212
R890 VGND.n1969 VGND.n1095 257.212
R891 VGND.n1969 VGND.n1094 257.212
R892 VGND.n1969 VGND.n1093 257.212
R893 VGND.n1969 VGND.n1092 257.212
R894 VGND.n1969 VGND.n1091 257.212
R895 VGND.n1969 VGND.n1090 257.212
R896 VGND.n1969 VGND.n1089 257.212
R897 VGND.n1969 VGND.n1088 257.212
R898 VGND.n1969 VGND.n1087 257.212
R899 VGND.n1617 VGND.n1616 257.212
R900 VGND.n1617 VGND.n1569 257.212
R901 VGND.n1617 VGND.n1570 257.212
R902 VGND.n1617 VGND.n1571 257.212
R903 VGND.n1617 VGND.n1572 257.212
R904 VGND.n1617 VGND.n1573 257.212
R905 VGND.n1617 VGND.n1574 257.212
R906 VGND.n1617 VGND.n1575 257.212
R907 VGND.n1617 VGND.n1576 257.212
R908 VGND.n1617 VGND.n1577 257.212
R909 VGND.n2436 VGND.n2435 257.212
R910 VGND.n2436 VGND.n699 257.212
R911 VGND.n2436 VGND.n700 257.212
R912 VGND.n2436 VGND.n701 257.212
R913 VGND.n2436 VGND.n702 257.212
R914 VGND.n2436 VGND.n703 257.212
R915 VGND.n2436 VGND.n704 257.212
R916 VGND.n2436 VGND.n705 257.212
R917 VGND.n2436 VGND.n706 257.212
R918 VGND.n2436 VGND.n707 257.212
R919 VGND.n2372 VGND.n759 257.212
R920 VGND.n2372 VGND.n760 257.212
R921 VGND.n2372 VGND.n761 257.212
R922 VGND.n2372 VGND.n762 257.212
R923 VGND.n2372 VGND.n763 257.212
R924 VGND.n2372 VGND.n764 257.212
R925 VGND.n2372 VGND.n765 257.212
R926 VGND.n2372 VGND.n766 257.212
R927 VGND.n2372 VGND.n767 257.212
R928 VGND.n2372 VGND.n768 257.212
R929 VGND.n2727 VGND.n50 257.212
R930 VGND.n2727 VGND.n51 257.212
R931 VGND.n2727 VGND.n52 257.212
R932 VGND.n2727 VGND.n53 257.212
R933 VGND.n2727 VGND.n54 257.212
R934 VGND.n2727 VGND.n55 257.212
R935 VGND.n2727 VGND.n56 257.212
R936 VGND.n2727 VGND.n57 257.212
R937 VGND.n2727 VGND.n58 257.212
R938 VGND.n2727 VGND.n59 257.212
R939 VGND.n2727 VGND.n60 257.212
R940 VGND.n2727 VGND.n61 257.212
R941 VGND.n2727 VGND.n62 257.212
R942 VGND.n2727 VGND.n63 257.212
R943 VGND.n2727 VGND.n64 257.212
R944 VGND.n2727 VGND.n65 257.212
R945 VGND.n2727 VGND.n66 257.212
R946 VGND.n2727 VGND.n67 257.212
R947 VGND.n2727 VGND.n68 257.212
R948 VGND.n2727 VGND.n69 257.212
R949 VGND.n2727 VGND.n70 257.212
R950 VGND.n2727 VGND.n71 257.212
R951 VGND.n2727 VGND.n72 257.212
R952 VGND.n2727 VGND.n73 257.212
R953 VGND.n2727 VGND.n74 257.212
R954 VGND.n2727 VGND.n75 257.212
R955 VGND.n2727 VGND.n76 257.212
R956 VGND.n2727 VGND.n77 257.212
R957 VGND.n2727 VGND.n78 257.212
R958 VGND.n2727 VGND.n79 257.212
R959 VGND.n2438 VGND.n542 257.212
R960 VGND.n2439 VGND.n2438 257.212
R961 VGND.n2438 VGND.n545 257.212
R962 VGND.n2438 VGND.n546 257.212
R963 VGND.n2438 VGND.n547 257.212
R964 VGND.n2438 VGND.n548 257.212
R965 VGND.n2438 VGND.n549 257.212
R966 VGND.n2438 VGND.n573 257.212
R967 VGND.n2500 VGND.n2499 257.212
R968 VGND.n2500 VGND.n532 257.212
R969 VGND.n2500 VGND.n533 257.212
R970 VGND.n2500 VGND.n534 257.212
R971 VGND.n2500 VGND.n535 257.212
R972 VGND.n2500 VGND.n536 257.212
R973 VGND.n2500 VGND.n537 257.212
R974 VGND.n2500 VGND.n538 257.212
R975 VGND.n2501 VGND.n2500 257.212
R976 VGND.n666 VGND.n665 257.212
R977 VGND.n666 VGND.n574 257.212
R978 VGND.n666 VGND.n575 257.212
R979 VGND.n666 VGND.n576 257.212
R980 VGND.n666 VGND.n577 257.212
R981 VGND.n666 VGND.n578 257.212
R982 VGND.n666 VGND.n579 257.212
R983 VGND.n666 VGND.n580 257.212
R984 VGND.n666 VGND.n581 257.212
R985 VGND.n524 VGND.n159 234.508
R986 VGND.n525 VGND.n524 234.508
R987 VGND.n526 VGND.n525 234.508
R988 VGND.n2524 VGND.n160 233.371
R989 VGND.n169 VGND.n160 233.371
R990 VGND.n2509 VGND.n169 233.371
R991 VGND.n1075 VGND.n1041 231.511
R992 VGND.n1077 VGND.n1076 231.511
R993 VGND.n1083 VGND.n1036 231.511
R994 VGND.n2719 VGND.n85 231.441
R995 VGND.n2718 VGND.n2717 231.441
R996 VGND.n2711 VGND.n2710 231.441
R997 VGND.n2709 VGND.n91 231.441
R998 VGND.n2702 VGND.n2701 231.441
R999 VGND.n2695 VGND.n97 231.441
R1000 VGND.n2694 VGND.n2693 231.441
R1001 VGND.n2685 VGND.n102 231.441
R1002 VGND.n2671 VGND.n109 231.441
R1003 VGND.n2663 VGND.n2662 231.441
R1004 VGND.n2654 VGND.n2653 231.441
R1005 VGND.n2645 VGND.n122 231.441
R1006 VGND.n2637 VGND.n126 231.441
R1007 VGND.n2629 VGND.n130 231.441
R1008 VGND.n2623 VGND.n2622 231.441
R1009 VGND.n2621 VGND.n135 231.441
R1010 VGND.n2615 VGND.n2614 231.441
R1011 VGND.n2613 VGND.n139 231.441
R1012 VGND.n2607 VGND.n2606 231.441
R1013 VGND.n2327 VGND.n771 230.065
R1014 VGND.n2325 VGND.n772 230.065
R1015 VGND.n2318 VGND.n2317 230.065
R1016 VGND.n2311 VGND.n779 230.065
R1017 VGND.n2309 VGND.n780 230.065
R1018 VGND.n2302 VGND.n2301 230.065
R1019 VGND.n2295 VGND.n787 230.065
R1020 VGND.n2294 VGND.n2293 230.065
R1021 VGND.n1922 VGND.n1121 227.434
R1022 VGND.n2285 VGND.n2284 227.434
R1023 VGND.n1694 VGND.n1693 225.392
R1024 VGND.n2385 VGND.n2384 225.392
R1025 VGND.n1975 VGND.n1974 195.556
R1026 VGND.n1970 VGND.n1969 190
R1027 VGND.n583 VGND.n582 160.519
R1028 VGND.n602 VGND.n582 160.519
R1029 VGND.n615 VGND.n614 160.519
R1030 VGND.n619 VGND.n618 160.519
R1031 VGND.n623 VGND.n622 160.519
R1032 VGND.n627 VGND.n626 160.519
R1033 VGND.n631 VGND.n630 160.519
R1034 VGND.n635 VGND.n634 160.519
R1035 VGND.n639 VGND.n638 160.519
R1036 VGND.n540 VGND.n539 160.519
R1037 VGND.n2493 VGND.n539 160.519
R1038 VGND.n2491 VGND.n2490 160.519
R1039 VGND.n2487 VGND.n2486 160.519
R1040 VGND.n2483 VGND.n2482 160.519
R1041 VGND.n2479 VGND.n2478 160.519
R1042 VGND.n2475 VGND.n2474 160.519
R1043 VGND.n2471 VGND.n2470 160.519
R1044 VGND.n2467 VGND.n531 160.519
R1045 VGND.n2441 VGND.n2440 160.519
R1046 VGND.n552 VGND.n544 160.519
R1047 VGND.n556 VGND.n555 160.519
R1048 VGND.n560 VGND.n559 160.519
R1049 VGND.n564 VGND.n563 160.519
R1050 VGND.n568 VGND.n567 160.519
R1051 VGND.n572 VGND.n550 160.519
R1052 VGND.n2331 VGND.n769 160.519
R1053 VGND.n2328 VGND.n769 160.519
R1054 VGND.n2328 VGND.n770 160.519
R1055 VGND.n2324 VGND.n770 160.519
R1056 VGND.n2324 VGND.n773 160.519
R1057 VGND.n2320 VGND.n773 160.519
R1058 VGND.n2320 VGND.n775 160.519
R1059 VGND.n2316 VGND.n775 160.519
R1060 VGND.n2316 VGND.n776 160.519
R1061 VGND.n2312 VGND.n776 160.519
R1062 VGND.n2312 VGND.n778 160.519
R1063 VGND.n2308 VGND.n778 160.519
R1064 VGND.n2308 VGND.n781 160.519
R1065 VGND.n2304 VGND.n781 160.519
R1066 VGND.n2304 VGND.n783 160.519
R1067 VGND.n2300 VGND.n783 160.519
R1068 VGND.n2300 VGND.n784 160.519
R1069 VGND.n2296 VGND.n784 160.519
R1070 VGND.n2296 VGND.n786 160.519
R1071 VGND.n2292 VGND.n786 160.519
R1072 VGND.n2292 VGND.n788 160.519
R1073 VGND.n2195 VGND.n2194 160.519
R1074 VGND.n2191 VGND.n2190 160.519
R1075 VGND.n2187 VGND.n2186 160.519
R1076 VGND.n2183 VGND.n2182 160.519
R1077 VGND.n2179 VGND.n2178 160.519
R1078 VGND.n2175 VGND.n2174 160.519
R1079 VGND.n2171 VGND.n2170 160.519
R1080 VGND.n2167 VGND.n2166 160.519
R1081 VGND.n2163 VGND.n2162 160.519
R1082 VGND.n2159 VGND.n2158 160.519
R1083 VGND.n2155 VGND.n2154 160.519
R1084 VGND.n2151 VGND.n2150 160.519
R1085 VGND.n2147 VGND.n2146 160.519
R1086 VGND.n2143 VGND.n2142 160.519
R1087 VGND.n2139 VGND.n2138 160.519
R1088 VGND.n2135 VGND.n2134 160.519
R1089 VGND.n2131 VGND.n2130 160.519
R1090 VGND.n2127 VGND.n2126 160.519
R1091 VGND.n2123 VGND.n2122 160.519
R1092 VGND.n2119 VGND.n2118 160.519
R1093 VGND.n2115 VGND.n2114 160.519
R1094 VGND.n2111 VGND.n2110 160.519
R1095 VGND.n2107 VGND.n2106 160.519
R1096 VGND.n2103 VGND.n2102 160.519
R1097 VGND.n2099 VGND.n2098 160.519
R1098 VGND.n2095 VGND.n2094 160.519
R1099 VGND.n2091 VGND.n2090 160.519
R1100 VGND.n2087 VGND.n2086 160.519
R1101 VGND.n2083 VGND.n2082 160.519
R1102 VGND.n2728 VGND.n49 160.519
R1103 VGND.n710 VGND.n709 160.519
R1104 VGND.n2431 VGND.n709 160.519
R1105 VGND.n2429 VGND.n2428 160.519
R1106 VGND.n2425 VGND.n2424 160.519
R1107 VGND.n2421 VGND.n2420 160.519
R1108 VGND.n2417 VGND.n2416 160.519
R1109 VGND.n2413 VGND.n2412 160.519
R1110 VGND.n2409 VGND.n2408 160.519
R1111 VGND.n2405 VGND.n2404 160.519
R1112 VGND.n2401 VGND.n2400 160.519
R1113 VGND.n2397 VGND.n708 160.519
R1114 VGND.n1579 VGND.n1578 160.519
R1115 VGND.n1612 VGND.n1578 160.519
R1116 VGND.n1610 VGND.n1609 160.519
R1117 VGND.n1606 VGND.n1605 160.519
R1118 VGND.n1602 VGND.n1601 160.519
R1119 VGND.n1598 VGND.n1597 160.519
R1120 VGND.n1594 VGND.n1593 160.519
R1121 VGND.n1590 VGND.n1589 160.519
R1122 VGND.n1586 VGND.n1585 160.519
R1123 VGND.n1582 VGND.n1581 160.519
R1124 VGND.n1618 VGND.n1568 160.519
R1125 VGND.n1967 VGND.n1097 160.519
R1126 VGND.n1963 VGND.n1096 160.519
R1127 VGND.n1961 VGND.n1960 160.519
R1128 VGND.n1957 VGND.n1956 160.519
R1129 VGND.n1953 VGND.n1952 160.519
R1130 VGND.n1949 VGND.n1948 160.519
R1131 VGND.n1945 VGND.n1944 160.519
R1132 VGND.n1941 VGND.n1940 160.519
R1133 VGND.n1937 VGND.n1936 160.519
R1134 VGND.n1933 VGND.n1932 160.519
R1135 VGND.n1929 VGND.n1086 160.519
R1136 VGND.n1277 VGND.n1276 160.519
R1137 VGND.n1281 VGND.n1280 160.519
R1138 VGND.n1285 VGND.n1284 160.519
R1139 VGND.n1289 VGND.n1288 160.519
R1140 VGND.n1293 VGND.n1292 160.519
R1141 VGND.n1297 VGND.n1296 160.519
R1142 VGND.n1301 VGND.n1300 160.519
R1143 VGND.n1305 VGND.n1304 160.519
R1144 VGND.n1309 VGND.n1308 160.519
R1145 VGND.n1313 VGND.n1312 160.519
R1146 VGND.n1317 VGND.n1316 160.519
R1147 VGND.n1321 VGND.n1320 160.519
R1148 VGND.n1325 VGND.n1324 160.519
R1149 VGND.n1329 VGND.n1328 160.519
R1150 VGND.n1333 VGND.n1332 160.519
R1151 VGND.n1337 VGND.n1336 160.519
R1152 VGND.n1341 VGND.n1340 160.519
R1153 VGND.n1345 VGND.n1344 160.519
R1154 VGND.n1349 VGND.n1348 160.519
R1155 VGND.n1353 VGND.n1352 160.519
R1156 VGND.n1357 VGND.n1356 160.519
R1157 VGND.n1361 VGND.n1360 160.519
R1158 VGND.n1365 VGND.n1364 160.519
R1159 VGND.n1369 VGND.n1368 160.519
R1160 VGND.n1373 VGND.n1372 160.519
R1161 VGND.n1377 VGND.n1376 160.519
R1162 VGND.n1381 VGND.n1380 160.519
R1163 VGND.n1385 VGND.n1384 160.519
R1164 VGND.n1389 VGND.n1388 160.519
R1165 VGND.n1391 VGND.n698 160.519
R1166 VGND.n1901 VGND.n1900 160.519
R1167 VGND.n1898 VGND.n1446 160.519
R1168 VGND.n1894 VGND.n1892 160.519
R1169 VGND.n1889 VGND.n1888 160.519
R1170 VGND.n1885 VGND.n1884 160.519
R1171 VGND.n1881 VGND.n1880 160.519
R1172 VGND.n1878 VGND.n1451 160.519
R1173 VGND.n1874 VGND.n1872 160.519
R1174 VGND.n1870 VGND.n1453 160.519
R1175 VGND.n1866 VGND.n1864 160.519
R1176 VGND.n1861 VGND.n1860 160.519
R1177 VGND.n1857 VGND.n1856 160.519
R1178 VGND.n1853 VGND.n1852 160.519
R1179 VGND.n1850 VGND.n1458 160.519
R1180 VGND.n1846 VGND.n1844 160.519
R1181 VGND.n1841 VGND.n1840 160.519
R1182 VGND.n1837 VGND.n1836 160.519
R1183 VGND.n1833 VGND.n1832 160.519
R1184 VGND.n1830 VGND.n1463 160.519
R1185 VGND.n1826 VGND.n1824 160.519
R1186 VGND.n1821 VGND.n1820 160.519
R1187 VGND.n1817 VGND.n1816 160.519
R1188 VGND.n1813 VGND.n1812 160.519
R1189 VGND.n1809 VGND.n1808 160.519
R1190 VGND.n1805 VGND.n1804 160.519
R1191 VGND.n1801 VGND.n1800 160.519
R1192 VGND.n1797 VGND.n1796 160.519
R1193 VGND.n1793 VGND.n1792 160.519
R1194 VGND.n1789 VGND.n1788 160.519
R1195 VGND.n1785 VGND.n1784 160.519
R1196 VGND.n1976 VGND.n1032 160.519
R1197 VGND.n1976 VGND.n1021 160.519
R1198 VGND.n1981 VGND.n1021 160.519
R1199 VGND.n1981 VGND.n1022 160.519
R1200 VGND.n1985 VGND.n887 160.519
R1201 VGND.n916 VGND.n888 160.519
R1202 VGND.n920 VGND.n919 160.519
R1203 VGND.n924 VGND.n923 160.519
R1204 VGND.n928 VGND.n927 160.519
R1205 VGND.n932 VGND.n931 160.519
R1206 VGND.n936 VGND.n935 160.519
R1207 VGND.n940 VGND.n939 160.519
R1208 VGND.n944 VGND.n943 160.519
R1209 VGND.n948 VGND.n947 160.519
R1210 VGND.n952 VGND.n951 160.519
R1211 VGND.n956 VGND.n955 160.519
R1212 VGND.n960 VGND.n959 160.519
R1213 VGND.n964 VGND.n963 160.519
R1214 VGND.n968 VGND.n967 160.519
R1215 VGND.n972 VGND.n971 160.519
R1216 VGND.n976 VGND.n975 160.519
R1217 VGND.n980 VGND.n979 160.519
R1218 VGND.n984 VGND.n983 160.519
R1219 VGND.n988 VGND.n987 160.519
R1220 VGND.n992 VGND.n991 160.519
R1221 VGND.n996 VGND.n995 160.519
R1222 VGND.n1000 VGND.n999 160.519
R1223 VGND.n1004 VGND.n1003 160.519
R1224 VGND.n1008 VGND.n1007 160.519
R1225 VGND.n1012 VGND.n1011 160.519
R1226 VGND.n1016 VGND.n915 160.519
R1227 VGND.n1019 VGND.n1018 160.519
R1228 VGND.n2371 VGND.n2333 160.519
R1229 VGND.n2368 VGND.n2367 160.519
R1230 VGND.n2364 VGND.n2363 160.519
R1231 VGND.n2360 VGND.n2359 160.519
R1232 VGND.n2356 VGND.n2355 160.519
R1233 VGND.n2352 VGND.n2351 160.519
R1234 VGND.n2348 VGND.n2347 160.519
R1235 VGND.n2344 VGND.n2343 160.519
R1236 VGND.n2340 VGND.n2339 160.519
R1237 VGND.n2336 VGND.n2335 160.519
R1238 VGND.n2373 VGND.n758 160.519
R1239 VGND.n2724 VGND.n83 160.519
R1240 VGND.n2720 VGND.n83 160.519
R1241 VGND.n2720 VGND.n84 160.519
R1242 VGND.n2716 VGND.n84 160.519
R1243 VGND.n2716 VGND.n86 160.519
R1244 VGND.n2712 VGND.n86 160.519
R1245 VGND.n2712 VGND.n89 160.519
R1246 VGND.n2708 VGND.n89 160.519
R1247 VGND.n2708 VGND.n92 160.519
R1248 VGND.n2704 VGND.n92 160.519
R1249 VGND.n2704 VGND.n93 160.519
R1250 VGND.n2700 VGND.n93 160.519
R1251 VGND.n2700 VGND.n94 160.519
R1252 VGND.n2696 VGND.n94 160.519
R1253 VGND.n2696 VGND.n96 160.519
R1254 VGND.n2692 VGND.n96 160.519
R1255 VGND.n2692 VGND.n98 160.519
R1256 VGND.n2688 VGND.n98 160.519
R1257 VGND.n2688 VGND.n100 160.519
R1258 VGND.n2684 VGND.n100 160.519
R1259 VGND.n2684 VGND.n103 160.519
R1260 VGND.n2680 VGND.n103 160.519
R1261 VGND.n2680 VGND.n105 160.519
R1262 VGND.n2676 VGND.n105 160.519
R1263 VGND.n2676 VGND.n106 160.519
R1264 VGND.n2672 VGND.n106 160.519
R1265 VGND.n2672 VGND.n108 160.519
R1266 VGND.n2668 VGND.n108 160.519
R1267 VGND.n2668 VGND.n110 160.519
R1268 VGND.n2664 VGND.n110 160.519
R1269 VGND.n2664 VGND.n113 160.519
R1270 VGND.n2660 VGND.n113 160.519
R1271 VGND.n2660 VGND.n115 160.519
R1272 VGND.n2656 VGND.n115 160.519
R1273 VGND.n2656 VGND.n116 160.519
R1274 VGND.n2652 VGND.n116 160.519
R1275 VGND.n2652 VGND.n118 160.519
R1276 VGND.n2648 VGND.n118 160.519
R1277 VGND.n2648 VGND.n120 160.519
R1278 VGND.n2644 VGND.n120 160.519
R1279 VGND.n2644 VGND.n123 160.519
R1280 VGND.n2640 VGND.n123 160.519
R1281 VGND.n2640 VGND.n125 160.519
R1282 VGND.n2636 VGND.n125 160.519
R1283 VGND.n2636 VGND.n127 160.519
R1284 VGND.n2632 VGND.n127 160.519
R1285 VGND.n2632 VGND.n129 160.519
R1286 VGND.n2628 VGND.n129 160.519
R1287 VGND.n2628 VGND.n131 160.519
R1288 VGND.n2624 VGND.n131 160.519
R1289 VGND.n2624 VGND.n134 160.519
R1290 VGND.n2620 VGND.n134 160.519
R1291 VGND.n2620 VGND.n136 160.519
R1292 VGND.n2616 VGND.n136 160.519
R1293 VGND.n2616 VGND.n138 160.519
R1294 VGND.n2612 VGND.n138 160.519
R1295 VGND.n2612 VGND.n140 160.519
R1296 VGND.n2608 VGND.n140 160.519
R1297 VGND.n2608 VGND.n142 160.519
R1298 VGND.n2604 VGND.n142 160.519
R1299 VGND.n1044 VGND.n1042 160.519
R1300 VGND.n1074 VGND.n1042 160.519
R1301 VGND.n1074 VGND.n1040 160.519
R1302 VGND.n1078 VGND.n1040 160.519
R1303 VGND.n1078 VGND.n1037 160.519
R1304 VGND.n1082 VGND.n1037 160.519
R1305 VGND.n1082 VGND.n1038 160.519
R1306 VGND.n1983 VGND.n1982 146.667
R1307 VGND.n2451 VGND.t37 136.786
R1308 VGND.n2447 VGND.t44 136.786
R1309 VGND.n2505 VGND.t47 136.786
R1310 VGND.n2463 VGND.t36 136.786
R1311 VGND.n2449 VGND.t182 136.786
R1312 VGND.n2452 VGND.t241 136.786
R1313 VGND.n2453 VGND.t302 136.786
R1314 VGND.n2456 VGND.t353 136.786
R1315 VGND.n529 VGND.t46 136.786
R1316 VGND.n2444 VGND.t43 136.786
R1317 VGND.n2597 VGND.t108 136.786
R1318 VGND.n739 VGND.t211 136.786
R1319 VGND.n740 VGND.t296 136.786
R1320 VGND.n742 VGND.t176 136.786
R1321 VGND.n744 VGND.t193 136.786
R1322 VGND.n746 VGND.t177 136.786
R1323 VGND.n748 VGND.t462 136.786
R1324 VGND.n750 VGND.t400 136.786
R1325 VGND.n752 VGND.t436 136.786
R1326 VGND.n1145 VGND.t117 136.786
R1327 VGND.n1124 VGND.t230 136.786
R1328 VGND.n1125 VGND.t270 136.786
R1329 VGND.n1127 VGND.t21 136.786
R1330 VGND.n1129 VGND.t506 136.786
R1331 VGND.n1131 VGND.t249 136.786
R1332 VGND.n1133 VGND.t165 136.786
R1333 VGND.n1135 VGND.t20 136.786
R1334 VGND.n1140 VGND.t166 136.786
R1335 VGND.n1142 VGND.t24 136.786
R1336 VGND.n1148 VGND.t118 136.786
R1337 VGND.n2024 VGND.t138 136.786
R1338 VGND.n1675 VGND.t58 136.786
R1339 VGND.n1659 VGND.t222 136.786
R1340 VGND.n1660 VGND.t379 136.786
R1341 VGND.n1662 VGND.t175 136.786
R1342 VGND.n1664 VGND.t179 136.786
R1343 VGND.n1666 VGND.t174 136.786
R1344 VGND.n1668 VGND.t485 136.786
R1345 VGND.n1670 VGND.t391 136.786
R1346 VGND.n1672 VGND.t433 136.786
R1347 VGND.n1678 VGND.t59 136.786
R1348 VGND.n1203 VGND.t97 136.786
R1349 VGND.n1271 VGND.t98 136.786
R1350 VGND.n1240 VGND.t131 136.786
R1351 VGND.n1237 VGND.t130 136.786
R1352 VGND.n1205 VGND.t157 136.786
R1353 VGND.n1206 VGND.t156 136.786
R1354 VGND.n1207 VGND.t242 136.786
R1355 VGND.n1208 VGND.t210 136.786
R1356 VGND.n1209 VGND.t266 136.786
R1357 VGND.n1210 VGND.t265 136.786
R1358 VGND.n1211 VGND.t184 136.786
R1359 VGND.n1214 VGND.t507 136.786
R1360 VGND.n1215 VGND.t535 136.786
R1361 VGND.n1218 VGND.t533 136.786
R1362 VGND.n1219 VGND.t488 136.786
R1363 VGND.n1222 VGND.t487 136.786
R1364 VGND.n1223 VGND.t329 136.786
R1365 VGND.n1226 VGND.t328 136.786
R1366 VGND.n1227 VGND.t311 136.786
R1367 VGND.n1230 VGND.t310 136.786
R1368 VGND.n1231 VGND.t362 136.786
R1369 VGND.n1232 VGND.t542 136.786
R1370 VGND.n1233 VGND.t183 136.786
R1371 VGND.n1234 VGND.t200 136.786
R1372 VGND.n1235 VGND.t551 136.786
R1373 VGND.n1236 VGND.t375 136.786
R1374 VGND.n1566 VGND.t121 136.786
R1375 VGND.n1550 VGND.t219 136.786
R1376 VGND.n1551 VGND.t279 136.786
R1377 VGND.n1553 VGND.t198 136.786
R1378 VGND.n1555 VGND.t204 136.786
R1379 VGND.n1557 VGND.t199 136.786
R1380 VGND.n1559 VGND.t446 136.786
R1381 VGND.n1561 VGND.t358 136.786
R1382 VGND.n1563 VGND.t437 136.786
R1383 VGND.n1649 VGND.t122 136.786
R1384 VGND.n1905 VGND.t125 136.786
R1385 VGND.n1533 VGND.t94 136.786
R1386 VGND.n1536 VGND.t93 136.786
R1387 VGND.n1474 VGND.t255 136.786
R1388 VGND.n1476 VGND.t213 136.786
R1389 VGND.n1478 VGND.t185 136.786
R1390 VGND.n1480 VGND.t164 136.786
R1391 VGND.n1482 VGND.t246 136.786
R1392 VGND.n1484 VGND.t245 136.786
R1393 VGND.n1486 VGND.t243 136.786
R1394 VGND.n1491 VGND.t520 136.786
R1395 VGND.n1493 VGND.t405 136.786
R1396 VGND.n1498 VGND.t404 136.786
R1397 VGND.n1500 VGND.t332 136.786
R1398 VGND.n1505 VGND.t334 136.786
R1399 VGND.n1507 VGND.t423 136.786
R1400 VGND.n1512 VGND.t422 136.786
R1401 VGND.n1514 VGND.t161 136.786
R1402 VGND.n1519 VGND.t160 136.786
R1403 VGND.n1521 VGND.t372 136.786
R1404 VGND.n1523 VGND.t548 136.786
R1405 VGND.n1525 VGND.t244 136.786
R1406 VGND.n1527 VGND.t150 136.786
R1407 VGND.n1529 VGND.t543 136.786
R1408 VGND.n1531 VGND.t374 136.786
R1409 VGND.n1907 VGND.t124 136.786
R1410 VGND.n1990 VGND.t86 136.786
R1411 VGND.n2027 VGND.t137 136.786
R1412 VGND.n1992 VGND.t12 136.786
R1413 VGND.n1994 VGND.t432 136.786
R1414 VGND.n1996 VGND.t512 136.786
R1415 VGND.n1998 VGND.t220 136.786
R1416 VGND.n2000 VGND.t307 136.786
R1417 VGND.n2002 VGND.t308 136.786
R1418 VGND.n2004 VGND.t466 136.786
R1419 VGND.n2006 VGND.t383 136.786
R1420 VGND.n2011 VGND.t382 136.786
R1421 VGND.n2013 VGND.t315 136.786
R1422 VGND.n2018 VGND.t314 136.786
R1423 VGND.n2020 VGND.t465 136.786
R1424 VGND.n2022 VGND.t306 136.786
R1425 VGND.n884 VGND.t85 136.786
R1426 VGND.n2377 VGND.t135 136.786
R1427 VGND.n12 VGND.t114 136.786
R1428 VGND.n13 VGND.t115 136.786
R1429 VGND.n2732 VGND.t141 136.786
R1430 VGND.n46 VGND.t140 136.786
R1431 VGND.n14 VGND.t254 136.786
R1432 VGND.n15 VGND.t232 136.786
R1433 VGND.n16 VGND.t253 136.786
R1434 VGND.n17 VGND.t19 136.786
R1435 VGND.n18 VGND.t18 136.786
R1436 VGND.n19 VGND.t17 136.786
R1437 VGND.n20 VGND.t180 136.786
R1438 VGND.n23 VGND.t508 136.786
R1439 VGND.n24 VGND.t395 136.786
R1440 VGND.n27 VGND.t393 136.786
R1441 VGND.n28 VGND.t396 136.786
R1442 VGND.n31 VGND.t398 136.786
R1443 VGND.n32 VGND.t355 136.786
R1444 VGND.n35 VGND.t357 136.786
R1445 VGND.n36 VGND.t322 136.786
R1446 VGND.n39 VGND.t325 136.786
R1447 VGND.n40 VGND.t376 136.786
R1448 VGND.n41 VGND.t550 136.786
R1449 VGND.n42 VGND.t181 136.786
R1450 VGND.n43 VGND.t214 136.786
R1451 VGND.n44 VGND.t546 136.786
R1452 VGND.n45 VGND.t364 136.786
R1453 VGND.n755 VGND.t134 136.786
R1454 VGND.n790 VGND.t189 136.786
R1455 VGND.n791 VGND.t305 136.786
R1456 VGND.n793 VGND.t228 136.786
R1457 VGND.n795 VGND.t276 136.786
R1458 VGND.n797 VGND.t226 136.786
R1459 VGND.n799 VGND.t480 136.786
R1460 VGND.n801 VGND.t385 136.786
R1461 VGND.n803 VGND.t435 136.786
R1462 VGND.n2287 VGND.t149 136.786
R1463 VGND.n805 VGND.t148 136.786
R1464 VGND.n2536 VGND.t73 136.786
R1465 VGND.n2600 VGND.t107 136.786
R1466 VGND.n2538 VGND.t272 136.786
R1467 VGND.n2540 VGND.t348 136.786
R1468 VGND.n2542 VGND.t152 136.786
R1469 VGND.n2544 VGND.t15 136.786
R1470 VGND.n2546 VGND.t207 136.786
R1471 VGND.n2548 VGND.t209 136.786
R1472 VGND.n2550 VGND.t170 136.786
R1473 VGND.n2555 VGND.t529 136.786
R1474 VGND.n2557 VGND.t491 136.786
R1475 VGND.n2562 VGND.t495 136.786
R1476 VGND.n2564 VGND.t457 136.786
R1477 VGND.n2569 VGND.t455 136.786
R1478 VGND.n2571 VGND.t476 136.786
R1479 VGND.n2576 VGND.t484 136.786
R1480 VGND.n2578 VGND.t417 136.786
R1481 VGND.n2583 VGND.t419 136.786
R1482 VGND.n2585 VGND.t368 136.786
R1483 VGND.n2587 VGND.t537 136.786
R1484 VGND.n2589 VGND.t168 136.786
R1485 VGND.n2591 VGND.t264 136.786
R1486 VGND.n2593 VGND.t539 136.786
R1487 VGND.n2595 VGND.t366 136.786
R1488 VGND.n2533 VGND.t72 136.786
R1489 VGND.n2203 VGND.t203 135.31
R1490 VGND.n2204 VGND.t238 135.31
R1491 VGND.n2205 VGND.t202 135.31
R1492 VGND.n2206 VGND.t259 135.31
R1493 VGND.n2207 VGND.t257 135.31
R1494 VGND.n2208 VGND.t258 135.31
R1495 VGND.n2209 VGND.t317 135.31
R1496 VGND.n2212 VGND.t527 135.31
R1497 VGND.n2213 VGND.t28 135.31
R1498 VGND.n2216 VGND.t27 135.31
R1499 VGND.n2217 VGND.t444 135.31
R1500 VGND.n2220 VGND.t443 135.31
R1501 VGND.n2221 VGND.t467 135.31
R1502 VGND.n2224 VGND.t469 135.31
R1503 VGND.n2225 VGND.t499 135.31
R1504 VGND.n2228 VGND.t501 135.31
R1505 VGND.n2229 VGND.t373 135.31
R1506 VGND.n2230 VGND.t549 135.31
R1507 VGND.n2231 VGND.t316 135.31
R1508 VGND.n2232 VGND.t171 135.31
R1509 VGND.n2233 VGND.t541 135.31
R1510 VGND.n2234 VGND.t378 135.31
R1511 VGND.n810 VGND.t248 135.31
R1512 VGND.n811 VGND.t282 135.31
R1513 VGND.n813 VGND.t237 135.31
R1514 VGND.n815 VGND.t221 135.31
R1515 VGND.n817 VGND.t236 135.31
R1516 VGND.n819 VGND.t336 135.31
R1517 VGND.n821 VGND.t313 135.31
R1518 VGND.n823 VGND.t409 135.31
R1519 VGND.n1161 VGND.t252 135.31
R1520 VGND.n1162 VGND.t251 135.31
R1521 VGND.n1163 VGND.t256 135.31
R1522 VGND.n1164 VGND.t273 135.31
R1523 VGND.n1165 VGND.t194 135.31
R1524 VGND.n1166 VGND.t195 135.31
R1525 VGND.n1167 VGND.t359 135.31
R1526 VGND.n1170 VGND.t509 135.31
R1527 VGND.n1171 VGND.t345 135.31
R1528 VGND.n1174 VGND.t343 135.31
R1529 VGND.n1175 VGND.t337 135.31
R1530 VGND.n1178 VGND.t339 135.31
R1531 VGND.n1179 VGND.t471 135.31
R1532 VGND.n1182 VGND.t474 135.31
R1533 VGND.n1183 VGND.t319 135.31
R1534 VGND.n1186 VGND.t318 135.31
R1535 VGND.n1187 VGND.t363 135.31
R1536 VGND.n1188 VGND.t553 135.31
R1537 VGND.n1189 VGND.t360 135.31
R1538 VGND.n1190 VGND.t247 135.31
R1539 VGND.n1191 VGND.t545 135.31
R1540 VGND.n1192 VGND.t369 135.31
R1541 VGND.n713 VGND.t235 135.31
R1542 VGND.n714 VGND.t278 135.31
R1543 VGND.n716 VGND.t191 135.31
R1544 VGND.n718 VGND.t201 135.31
R1545 VGND.n720 VGND.t190 135.31
R1546 VGND.n722 VGND.t463 135.31
R1547 VGND.n724 VGND.t346 135.31
R1548 VGND.n726 VGND.t431 135.31
R1549 VGND.n1715 VGND.t205 135.31
R1550 VGND.n1717 VGND.t23 135.31
R1551 VGND.n1719 VGND.t267 135.31
R1552 VGND.n1721 VGND.t260 135.31
R1553 VGND.n1723 VGND.t218 135.31
R1554 VGND.n1725 VGND.t217 135.31
R1555 VGND.n1727 VGND.t331 135.31
R1556 VGND.n1732 VGND.t514 135.31
R1557 VGND.n1734 VGND.t285 135.31
R1558 VGND.n1739 VGND.t288 135.31
R1559 VGND.n1741 VGND.t290 135.31
R1560 VGND.n1746 VGND.t292 135.31
R1561 VGND.n1748 VGND.t439 135.31
R1562 VGND.n1753 VGND.t440 135.31
R1563 VGND.n1755 VGND.t349 135.31
R1564 VGND.n1760 VGND.t350 135.31
R1565 VGND.n1762 VGND.t370 135.31
R1566 VGND.n1764 VGND.t544 135.31
R1567 VGND.n1766 VGND.t330 135.31
R1568 VGND.n1768 VGND.t250 135.31
R1569 VGND.n1770 VGND.t552 135.31
R1570 VGND.n1772 VGND.t361 135.31
R1571 VGND.n1621 VGND.t231 135.31
R1572 VGND.n1622 VGND.t277 135.31
R1573 VGND.n1624 VGND.t154 135.31
R1574 VGND.n1626 VGND.t153 135.31
R1575 VGND.n1628 VGND.t155 135.31
R1576 VGND.n1630 VGND.t163 135.31
R1577 VGND.n1632 VGND.t294 135.31
R1578 VGND.n1634 VGND.t410 135.31
R1579 VGND.n848 VGND.t224 135.31
R1580 VGND.n849 VGND.t261 135.31
R1581 VGND.n850 VGND.t234 135.31
R1582 VGND.n851 VGND.t233 135.31
R1583 VGND.n852 VGND.t239 135.31
R1584 VGND.n853 VGND.t240 135.31
R1585 VGND.n854 VGND.t281 135.31
R1586 VGND.n857 VGND.t513 135.31
R1587 VGND.n858 VGND.t390 135.31
R1588 VGND.n861 VGND.t411 135.31
R1589 VGND.n862 VGND.t298 135.31
R1590 VGND.n865 VGND.t299 135.31
R1591 VGND.n866 VGND.t450 135.31
R1592 VGND.n869 VGND.t447 135.31
R1593 VGND.n870 VGND.t427 135.31
R1594 VGND.n873 VGND.t425 135.31
R1595 VGND.n874 VGND.t371 135.31
R1596 VGND.n875 VGND.t547 135.31
R1597 VGND.n876 VGND.t280 135.31
R1598 VGND.n877 VGND.t229 135.31
R1599 VGND.n878 VGND.t540 135.31
R1600 VGND.n879 VGND.t377 135.31
R1601 VGND.n1102 VGND.t158 135.31
R1602 VGND.n1103 VGND.t341 135.31
R1603 VGND.n1105 VGND.t216 135.31
R1604 VGND.n1107 VGND.t212 135.31
R1605 VGND.n1109 VGND.t215 135.31
R1606 VGND.n1111 VGND.t293 135.31
R1607 VGND.n1113 VGND.t295 135.31
R1608 VGND.n1115 VGND.t430 135.31
R1609 VGND.n590 VGND.t274 135.31
R1610 VGND.n593 VGND.t178 135.31
R1611 VGND.n594 VGND.t408 135.31
R1612 VGND.n597 VGND.t352 135.31
R1613 VGND.n1045 VGND.t112 131.389
R1614 VGND.n1048 VGND.t111 131.389
R1615 VGND.n587 VGND.t127 131.389
R1616 VGND.n644 VGND.t103 131.389
R1617 VGND.n647 VGND.t104 131.389
R1618 VGND.n608 VGND.t40 131.389
R1619 VGND.n605 VGND.t41 131.389
R1620 VGND.n585 VGND.t128 131.389
R1621 VGND.n2077 VGND.t82 131.389
R1622 VGND.n2238 VGND.t68 131.389
R1623 VGND.n2241 VGND.t69 131.389
R1624 VGND.n2200 VGND.t83 131.389
R1625 VGND.n832 VGND.t145 131.389
R1626 VGND.n827 VGND.t144 131.389
R1627 VGND.n1196 VGND.t61 131.389
R1628 VGND.n1396 VGND.t32 131.389
R1629 VGND.n1399 VGND.t33 131.389
R1630 VGND.n1199 VGND.t62 131.389
R1631 VGND.n712 VGND.t89 131.389
R1632 VGND.n728 VGND.t90 131.389
R1633 VGND.n1540 VGND.t76 131.389
R1634 VGND.n1706 VGND.t100 131.389
R1635 VGND.n1711 VGND.t101 131.389
R1636 VGND.n1620 VGND.t65 131.389
R1637 VGND.n1636 VGND.t66 131.389
R1638 VGND.n1774 VGND.t75 131.389
R1639 VGND.n1024 VGND.t54 131.389
R1640 VGND.n2033 VGND.t79 131.389
R1641 VGND.n2036 VGND.t80 131.389
R1642 VGND.n1027 VGND.t55 131.389
R1643 VGND.n1117 VGND.t50 131.389
R1644 VGND.n1100 VGND.t51 131.389
R1645 VGND.n1062 VGND.t269 131.389
R1646 VGND.n1057 VGND.t173 131.389
R1647 VGND.n1052 VGND.t429 131.389
R1648 VGND.n1971 VGND.n1084 129.032
R1649 VGND.n1922 VGND.n1921 116.118
R1650 VGND.n1043 VGND.t110 115.755
R1651 VGND.t110 VGND.n1041 115.755
R1652 VGND.t268 VGND.n1075 115.755
R1653 VGND.n1076 VGND.t268 115.755
R1654 VGND.n1077 VGND.t172 115.755
R1655 VGND.t172 VGND.n1036 115.755
R1656 VGND.n2725 VGND.t71 115.721
R1657 VGND.n85 VGND.t71 115.721
R1658 VGND.n2719 VGND.t271 115.721
R1659 VGND.t271 VGND.n2718 115.721
R1660 VGND.n2717 VGND.t347 115.721
R1661 VGND.n90 VGND.t347 115.721
R1662 VGND.t151 VGND.n90 115.721
R1663 VGND.n2711 VGND.t151 115.721
R1664 VGND.n2710 VGND.t14 115.721
R1665 VGND.t14 VGND.n2709 115.721
R1666 VGND.t13 VGND.n91 115.721
R1667 VGND.n2703 VGND.t13 115.721
R1668 VGND.n2703 VGND.t206 115.721
R1669 VGND.t206 VGND.n2702 115.721
R1670 VGND.n2701 VGND.t208 115.721
R1671 VGND.n97 VGND.t208 115.721
R1672 VGND.n2695 VGND.t169 115.721
R1673 VGND.t169 VGND.n2694 115.721
R1674 VGND.n2693 VGND.t523 115.721
R1675 VGND.n101 VGND.t523 115.721
R1676 VGND.t521 VGND.n101 115.721
R1677 VGND.n2687 VGND.t521 115.721
R1678 VGND.n2687 VGND.t530 115.721
R1679 VGND.t530 VGND.n2686 115.721
R1680 VGND.n2686 VGND.t528 115.721
R1681 VGND.t528 VGND.n2685 115.721
R1682 VGND.t490 VGND.n102 115.721
R1683 VGND.n2679 VGND.t490 115.721
R1684 VGND.n2679 VGND.t492 115.721
R1685 VGND.t492 VGND.n2678 115.721
R1686 VGND.n2678 VGND.t496 115.721
R1687 VGND.t496 VGND.n2677 115.721
R1688 VGND.n2677 VGND.t494 115.721
R1689 VGND.n109 VGND.t494 115.721
R1690 VGND.n2671 VGND.t456 115.721
R1691 VGND.t456 VGND.n2670 115.721
R1692 VGND.n2670 VGND.t458 115.721
R1693 VGND.t458 VGND.n2669 115.721
R1694 VGND.n2669 VGND.t460 115.721
R1695 VGND.n114 VGND.t460 115.721
R1696 VGND.t454 VGND.n114 115.721
R1697 VGND.n2663 VGND.t454 115.721
R1698 VGND.n2662 VGND.t475 115.721
R1699 VGND.t475 VGND.n2661 115.721
R1700 VGND.n2661 VGND.t481 115.721
R1701 VGND.n117 VGND.t481 115.721
R1702 VGND.t477 VGND.n117 115.721
R1703 VGND.n2655 VGND.t477 115.721
R1704 VGND.n2655 VGND.t483 115.721
R1705 VGND.t483 VGND.n2654 115.721
R1706 VGND.n2653 VGND.t416 115.721
R1707 VGND.n121 VGND.t416 115.721
R1708 VGND.t412 VGND.n121 115.721
R1709 VGND.n2647 VGND.t412 115.721
R1710 VGND.n2647 VGND.t414 115.721
R1711 VGND.t414 VGND.n2646 115.721
R1712 VGND.n2646 VGND.t418 115.721
R1713 VGND.t418 VGND.n2645 115.721
R1714 VGND.t453 VGND.n122 115.721
R1715 VGND.n2639 VGND.t453 115.721
R1716 VGND.n2639 VGND.t197 115.721
R1717 VGND.t197 VGND.n2638 115.721
R1718 VGND.n2638 VGND.t367 115.721
R1719 VGND.t367 VGND.n2637 115.721
R1720 VGND.t452 VGND.n126 115.721
R1721 VGND.n2631 VGND.t452 115.721
R1722 VGND.n2631 VGND.t196 115.721
R1723 VGND.t196 VGND.n2630 115.721
R1724 VGND.n2630 VGND.t536 115.721
R1725 VGND.t536 VGND.n2629 115.721
R1726 VGND.t167 VGND.n130 115.721
R1727 VGND.n2623 VGND.t167 115.721
R1728 VGND.n2622 VGND.t263 115.721
R1729 VGND.t263 VGND.n2621 115.721
R1730 VGND.t538 VGND.n135 115.721
R1731 VGND.n2615 VGND.t538 115.721
R1732 VGND.n2614 VGND.t365 115.721
R1733 VGND.t365 VGND.n2613 115.721
R1734 VGND.t451 VGND.n139 115.721
R1735 VGND.n2607 VGND.t451 115.721
R1736 VGND.n2606 VGND.t106 115.721
R1737 VGND.t106 VGND.n2605 115.721
R1738 VGND.n2332 VGND.t188 115.034
R1739 VGND.n771 VGND.t188 115.034
R1740 VGND.n2327 VGND.t386 115.034
R1741 VGND.t386 VGND.n2326 115.034
R1742 VGND.n2326 VGND.t304 115.034
R1743 VGND.t304 VGND.n2325 115.034
R1744 VGND.t186 VGND.n772 115.034
R1745 VGND.n2319 VGND.t186 115.034
R1746 VGND.n2319 VGND.t227 115.034
R1747 VGND.t227 VGND.n2318 115.034
R1748 VGND.n2317 VGND.t275 115.034
R1749 VGND.n779 VGND.t275 115.034
R1750 VGND.n2311 VGND.t187 115.034
R1751 VGND.t187 VGND.n2310 115.034
R1752 VGND.n2310 VGND.t225 115.034
R1753 VGND.t225 VGND.n2309 115.034
R1754 VGND.t387 VGND.n780 115.034
R1755 VGND.n2303 VGND.t387 115.034
R1756 VGND.n2303 VGND.t479 115.034
R1757 VGND.t479 VGND.n2302 115.034
R1758 VGND.n2301 VGND.t384 115.034
R1759 VGND.n787 VGND.t384 115.034
R1760 VGND.n2295 VGND.t434 115.034
R1761 VGND.t434 VGND.n2294 115.034
R1762 VGND.n2293 VGND.t147 115.034
R1763 VGND.t147 VGND.n82 115.034
R1764 VGND.n1656 VGND.n1655 110.749
R1765 VGND.n1692 VGND.n735 110.749
R1766 VGND.n807 VGND.n736 110.749
R1767 VGND.n2455 VGND.n2454 97.8962
R1768 VGND.n1138 VGND.n1137 97.8962
R1769 VGND.n1213 VGND.n1212 97.8962
R1770 VGND.n1217 VGND.n1216 97.8962
R1771 VGND.n1221 VGND.n1220 97.8962
R1772 VGND.n1225 VGND.n1224 97.8962
R1773 VGND.n1229 VGND.n1228 97.8962
R1774 VGND.n1489 VGND.n1488 97.8962
R1775 VGND.n1496 VGND.n1495 97.8962
R1776 VGND.n1503 VGND.n1502 97.8962
R1777 VGND.n1510 VGND.n1509 97.8962
R1778 VGND.n1517 VGND.n1516 97.8962
R1779 VGND.n2009 VGND.n2008 97.8962
R1780 VGND.n2016 VGND.n2015 97.8962
R1781 VGND.n22 VGND.n21 97.8962
R1782 VGND.n26 VGND.n25 97.8962
R1783 VGND.n30 VGND.n29 97.8962
R1784 VGND.n34 VGND.n33 97.8962
R1785 VGND.n38 VGND.n37 97.8962
R1786 VGND.n2553 VGND.n2552 97.8962
R1787 VGND.n2560 VGND.n2559 97.8962
R1788 VGND.n2567 VGND.n2566 97.8962
R1789 VGND.n2574 VGND.n2573 97.8962
R1790 VGND.n2581 VGND.n2580 97.8962
R1791 VGND.t53 VGND.n1973 97.7783
R1792 VGND.n1975 VGND.t53 97.7783
R1793 VGND.n1974 VGND.t223 97.7783
R1794 VGND.n1982 VGND.t223 97.7783
R1795 VGND.n2211 VGND.n2210 96.4212
R1796 VGND.n2215 VGND.n2214 96.4212
R1797 VGND.n2219 VGND.n2218 96.4212
R1798 VGND.n2223 VGND.n2222 96.4212
R1799 VGND.n2227 VGND.n2226 96.4212
R1800 VGND.n1169 VGND.n1168 96.4212
R1801 VGND.n1173 VGND.n1172 96.4212
R1802 VGND.n1177 VGND.n1176 96.4212
R1803 VGND.n1181 VGND.n1180 96.4212
R1804 VGND.n1185 VGND.n1184 96.4212
R1805 VGND.n1730 VGND.n1729 96.4212
R1806 VGND.n1737 VGND.n1736 96.4212
R1807 VGND.n1744 VGND.n1743 96.4212
R1808 VGND.n1751 VGND.n1750 96.4212
R1809 VGND.n1758 VGND.n1757 96.4212
R1810 VGND.n856 VGND.n855 96.4212
R1811 VGND.n860 VGND.n859 96.4212
R1812 VGND.n864 VGND.n863 96.4212
R1813 VGND.n868 VGND.n867 96.4212
R1814 VGND.n872 VGND.n871 96.4212
R1815 VGND.n596 VGND.n595 96.4212
R1816 VGND.n1084 VGND.n1083 72.3473
R1817 VGND.n602 VGND.n574 70.5775
R1818 VGND.n615 VGND.n575 70.5775
R1819 VGND.n619 VGND.n576 70.5775
R1820 VGND.n623 VGND.n577 70.5775
R1821 VGND.n627 VGND.n578 70.5775
R1822 VGND.n631 VGND.n579 70.5775
R1823 VGND.n635 VGND.n580 70.5775
R1824 VGND.n639 VGND.n581 70.5775
R1825 VGND.n2493 VGND.n532 70.5775
R1826 VGND.n2490 VGND.n533 70.5775
R1827 VGND.n2486 VGND.n534 70.5775
R1828 VGND.n2482 VGND.n535 70.5775
R1829 VGND.n2478 VGND.n536 70.5775
R1830 VGND.n2474 VGND.n537 70.5775
R1831 VGND.n2470 VGND.n538 70.5775
R1832 VGND.n2501 VGND.n531 70.5775
R1833 VGND.n2440 VGND.n2439 70.5775
R1834 VGND.n552 VGND.n545 70.5775
R1835 VGND.n556 VGND.n546 70.5775
R1836 VGND.n560 VGND.n547 70.5775
R1837 VGND.n564 VGND.n548 70.5775
R1838 VGND.n568 VGND.n549 70.5775
R1839 VGND.n573 VGND.n572 70.5775
R1840 VGND.n2194 VGND.n51 70.5775
R1841 VGND.n2190 VGND.n52 70.5775
R1842 VGND.n2186 VGND.n53 70.5775
R1843 VGND.n2182 VGND.n54 70.5775
R1844 VGND.n2178 VGND.n55 70.5775
R1845 VGND.n2174 VGND.n56 70.5775
R1846 VGND.n2170 VGND.n57 70.5775
R1847 VGND.n2166 VGND.n58 70.5775
R1848 VGND.n2162 VGND.n59 70.5775
R1849 VGND.n2158 VGND.n60 70.5775
R1850 VGND.n2154 VGND.n61 70.5775
R1851 VGND.n2150 VGND.n62 70.5775
R1852 VGND.n2146 VGND.n63 70.5775
R1853 VGND.n2142 VGND.n64 70.5775
R1854 VGND.n2138 VGND.n65 70.5775
R1855 VGND.n2134 VGND.n66 70.5775
R1856 VGND.n2130 VGND.n67 70.5775
R1857 VGND.n2126 VGND.n68 70.5775
R1858 VGND.n2122 VGND.n69 70.5775
R1859 VGND.n2118 VGND.n70 70.5775
R1860 VGND.n2114 VGND.n71 70.5775
R1861 VGND.n2110 VGND.n72 70.5775
R1862 VGND.n2106 VGND.n73 70.5775
R1863 VGND.n2102 VGND.n74 70.5775
R1864 VGND.n2098 VGND.n75 70.5775
R1865 VGND.n2094 VGND.n76 70.5775
R1866 VGND.n2090 VGND.n77 70.5775
R1867 VGND.n2086 VGND.n78 70.5775
R1868 VGND.n2082 VGND.n79 70.5775
R1869 VGND.n2431 VGND.n699 70.5775
R1870 VGND.n2428 VGND.n700 70.5775
R1871 VGND.n2424 VGND.n701 70.5775
R1872 VGND.n2420 VGND.n702 70.5775
R1873 VGND.n2416 VGND.n703 70.5775
R1874 VGND.n2412 VGND.n704 70.5775
R1875 VGND.n2408 VGND.n705 70.5775
R1876 VGND.n2404 VGND.n706 70.5775
R1877 VGND.n2400 VGND.n707 70.5775
R1878 VGND.n1612 VGND.n1569 70.5775
R1879 VGND.n1609 VGND.n1570 70.5775
R1880 VGND.n1605 VGND.n1571 70.5775
R1881 VGND.n1601 VGND.n1572 70.5775
R1882 VGND.n1597 VGND.n1573 70.5775
R1883 VGND.n1593 VGND.n1574 70.5775
R1884 VGND.n1589 VGND.n1575 70.5775
R1885 VGND.n1585 VGND.n1576 70.5775
R1886 VGND.n1581 VGND.n1577 70.5775
R1887 VGND.n1097 VGND.n1085 70.5775
R1888 VGND.n1968 VGND.n1967 70.5775
R1889 VGND.n1963 VGND.n1095 70.5775
R1890 VGND.n1960 VGND.n1094 70.5775
R1891 VGND.n1956 VGND.n1093 70.5775
R1892 VGND.n1952 VGND.n1092 70.5775
R1893 VGND.n1948 VGND.n1091 70.5775
R1894 VGND.n1944 VGND.n1090 70.5775
R1895 VGND.n1940 VGND.n1089 70.5775
R1896 VGND.n1936 VGND.n1088 70.5775
R1897 VGND.n1932 VGND.n1087 70.5775
R1898 VGND.n1277 VGND.n669 70.5775
R1899 VGND.n1281 VGND.n670 70.5775
R1900 VGND.n1285 VGND.n671 70.5775
R1901 VGND.n1289 VGND.n672 70.5775
R1902 VGND.n1293 VGND.n673 70.5775
R1903 VGND.n1297 VGND.n674 70.5775
R1904 VGND.n1301 VGND.n675 70.5775
R1905 VGND.n1305 VGND.n676 70.5775
R1906 VGND.n1309 VGND.n677 70.5775
R1907 VGND.n1313 VGND.n678 70.5775
R1908 VGND.n1317 VGND.n679 70.5775
R1909 VGND.n1321 VGND.n680 70.5775
R1910 VGND.n1325 VGND.n681 70.5775
R1911 VGND.n1329 VGND.n682 70.5775
R1912 VGND.n1333 VGND.n683 70.5775
R1913 VGND.n1337 VGND.n684 70.5775
R1914 VGND.n1341 VGND.n685 70.5775
R1915 VGND.n1345 VGND.n686 70.5775
R1916 VGND.n1349 VGND.n687 70.5775
R1917 VGND.n1353 VGND.n688 70.5775
R1918 VGND.n1357 VGND.n689 70.5775
R1919 VGND.n1361 VGND.n690 70.5775
R1920 VGND.n1365 VGND.n691 70.5775
R1921 VGND.n1369 VGND.n692 70.5775
R1922 VGND.n1373 VGND.n693 70.5775
R1923 VGND.n1377 VGND.n694 70.5775
R1924 VGND.n1381 VGND.n695 70.5775
R1925 VGND.n1385 VGND.n696 70.5775
R1926 VGND.n1389 VGND.n697 70.5775
R1927 VGND.n1276 VGND.n668 70.5775
R1928 VGND.n1280 VGND.n669 70.5775
R1929 VGND.n1284 VGND.n670 70.5775
R1930 VGND.n1288 VGND.n671 70.5775
R1931 VGND.n1292 VGND.n672 70.5775
R1932 VGND.n1296 VGND.n673 70.5775
R1933 VGND.n1300 VGND.n674 70.5775
R1934 VGND.n1304 VGND.n675 70.5775
R1935 VGND.n1308 VGND.n676 70.5775
R1936 VGND.n1312 VGND.n677 70.5775
R1937 VGND.n1316 VGND.n678 70.5775
R1938 VGND.n1320 VGND.n679 70.5775
R1939 VGND.n1324 VGND.n680 70.5775
R1940 VGND.n1328 VGND.n681 70.5775
R1941 VGND.n1332 VGND.n682 70.5775
R1942 VGND.n1336 VGND.n683 70.5775
R1943 VGND.n1340 VGND.n684 70.5775
R1944 VGND.n1344 VGND.n685 70.5775
R1945 VGND.n1348 VGND.n686 70.5775
R1946 VGND.n1352 VGND.n687 70.5775
R1947 VGND.n1356 VGND.n688 70.5775
R1948 VGND.n1360 VGND.n689 70.5775
R1949 VGND.n1364 VGND.n690 70.5775
R1950 VGND.n1368 VGND.n691 70.5775
R1951 VGND.n1372 VGND.n692 70.5775
R1952 VGND.n1376 VGND.n693 70.5775
R1953 VGND.n1380 VGND.n694 70.5775
R1954 VGND.n1384 VGND.n695 70.5775
R1955 VGND.n1388 VGND.n696 70.5775
R1956 VGND.n1391 VGND.n697 70.5775
R1957 VGND.n1900 VGND.n1899 70.5775
R1958 VGND.n1893 VGND.n1446 70.5775
R1959 VGND.n1892 VGND.n1447 70.5775
R1960 VGND.n1888 VGND.n1448 70.5775
R1961 VGND.n1884 VGND.n1449 70.5775
R1962 VGND.n1880 VGND.n1879 70.5775
R1963 VGND.n1873 VGND.n1451 70.5775
R1964 VGND.n1872 VGND.n1871 70.5775
R1965 VGND.n1865 VGND.n1453 70.5775
R1966 VGND.n1864 VGND.n1454 70.5775
R1967 VGND.n1860 VGND.n1455 70.5775
R1968 VGND.n1856 VGND.n1456 70.5775
R1969 VGND.n1852 VGND.n1851 70.5775
R1970 VGND.n1845 VGND.n1458 70.5775
R1971 VGND.n1844 VGND.n1459 70.5775
R1972 VGND.n1840 VGND.n1460 70.5775
R1973 VGND.n1836 VGND.n1461 70.5775
R1974 VGND.n1832 VGND.n1831 70.5775
R1975 VGND.n1825 VGND.n1463 70.5775
R1976 VGND.n1824 VGND.n1464 70.5775
R1977 VGND.n1820 VGND.n1465 70.5775
R1978 VGND.n1816 VGND.n1466 70.5775
R1979 VGND.n1812 VGND.n1467 70.5775
R1980 VGND.n1808 VGND.n1468 70.5775
R1981 VGND.n1804 VGND.n1469 70.5775
R1982 VGND.n1800 VGND.n1470 70.5775
R1983 VGND.n1796 VGND.n1471 70.5775
R1984 VGND.n1792 VGND.n1472 70.5775
R1985 VGND.n1788 VGND.n1473 70.5775
R1986 VGND.n1901 VGND.n1444 70.5775
R1987 VGND.n1899 VGND.n1898 70.5775
R1988 VGND.n1894 VGND.n1893 70.5775
R1989 VGND.n1889 VGND.n1447 70.5775
R1990 VGND.n1885 VGND.n1448 70.5775
R1991 VGND.n1881 VGND.n1449 70.5775
R1992 VGND.n1879 VGND.n1878 70.5775
R1993 VGND.n1874 VGND.n1873 70.5775
R1994 VGND.n1871 VGND.n1870 70.5775
R1995 VGND.n1866 VGND.n1865 70.5775
R1996 VGND.n1861 VGND.n1454 70.5775
R1997 VGND.n1857 VGND.n1455 70.5775
R1998 VGND.n1853 VGND.n1456 70.5775
R1999 VGND.n1851 VGND.n1850 70.5775
R2000 VGND.n1846 VGND.n1845 70.5775
R2001 VGND.n1841 VGND.n1459 70.5775
R2002 VGND.n1837 VGND.n1460 70.5775
R2003 VGND.n1833 VGND.n1461 70.5775
R2004 VGND.n1831 VGND.n1830 70.5775
R2005 VGND.n1826 VGND.n1825 70.5775
R2006 VGND.n1821 VGND.n1464 70.5775
R2007 VGND.n1817 VGND.n1465 70.5775
R2008 VGND.n1813 VGND.n1466 70.5775
R2009 VGND.n1809 VGND.n1467 70.5775
R2010 VGND.n1805 VGND.n1468 70.5775
R2011 VGND.n1801 VGND.n1469 70.5775
R2012 VGND.n1797 VGND.n1470 70.5775
R2013 VGND.n1793 VGND.n1471 70.5775
R2014 VGND.n1789 VGND.n1472 70.5775
R2015 VGND.n1785 VGND.n1473 70.5775
R2016 VGND.n1022 VGND.n889 70.5775
R2017 VGND.n1985 VGND.n1984 70.5775
R2018 VGND.n916 VGND.n890 70.5775
R2019 VGND.n920 VGND.n891 70.5775
R2020 VGND.n924 VGND.n892 70.5775
R2021 VGND.n928 VGND.n893 70.5775
R2022 VGND.n932 VGND.n894 70.5775
R2023 VGND.n936 VGND.n895 70.5775
R2024 VGND.n940 VGND.n896 70.5775
R2025 VGND.n944 VGND.n897 70.5775
R2026 VGND.n948 VGND.n898 70.5775
R2027 VGND.n952 VGND.n899 70.5775
R2028 VGND.n956 VGND.n900 70.5775
R2029 VGND.n960 VGND.n901 70.5775
R2030 VGND.n964 VGND.n902 70.5775
R2031 VGND.n968 VGND.n903 70.5775
R2032 VGND.n972 VGND.n904 70.5775
R2033 VGND.n976 VGND.n905 70.5775
R2034 VGND.n980 VGND.n906 70.5775
R2035 VGND.n984 VGND.n907 70.5775
R2036 VGND.n988 VGND.n908 70.5775
R2037 VGND.n992 VGND.n909 70.5775
R2038 VGND.n996 VGND.n910 70.5775
R2039 VGND.n1000 VGND.n911 70.5775
R2040 VGND.n1004 VGND.n912 70.5775
R2041 VGND.n1008 VGND.n913 70.5775
R2042 VGND.n1012 VGND.n914 70.5775
R2043 VGND.n1017 VGND.n1016 70.5775
R2044 VGND.n889 VGND.n887 70.5775
R2045 VGND.n1984 VGND.n888 70.5775
R2046 VGND.n919 VGND.n890 70.5775
R2047 VGND.n923 VGND.n891 70.5775
R2048 VGND.n927 VGND.n892 70.5775
R2049 VGND.n931 VGND.n893 70.5775
R2050 VGND.n935 VGND.n894 70.5775
R2051 VGND.n939 VGND.n895 70.5775
R2052 VGND.n943 VGND.n896 70.5775
R2053 VGND.n947 VGND.n897 70.5775
R2054 VGND.n951 VGND.n898 70.5775
R2055 VGND.n955 VGND.n899 70.5775
R2056 VGND.n959 VGND.n900 70.5775
R2057 VGND.n963 VGND.n901 70.5775
R2058 VGND.n967 VGND.n902 70.5775
R2059 VGND.n971 VGND.n903 70.5775
R2060 VGND.n975 VGND.n904 70.5775
R2061 VGND.n979 VGND.n905 70.5775
R2062 VGND.n983 VGND.n906 70.5775
R2063 VGND.n987 VGND.n907 70.5775
R2064 VGND.n991 VGND.n908 70.5775
R2065 VGND.n995 VGND.n909 70.5775
R2066 VGND.n999 VGND.n910 70.5775
R2067 VGND.n1003 VGND.n911 70.5775
R2068 VGND.n1007 VGND.n912 70.5775
R2069 VGND.n1011 VGND.n913 70.5775
R2070 VGND.n915 VGND.n914 70.5775
R2071 VGND.n1018 VGND.n1017 70.5775
R2072 VGND.n1968 VGND.n1096 70.5775
R2073 VGND.n1961 VGND.n1095 70.5775
R2074 VGND.n1957 VGND.n1094 70.5775
R2075 VGND.n1953 VGND.n1093 70.5775
R2076 VGND.n1949 VGND.n1092 70.5775
R2077 VGND.n1945 VGND.n1091 70.5775
R2078 VGND.n1941 VGND.n1090 70.5775
R2079 VGND.n1937 VGND.n1089 70.5775
R2080 VGND.n1933 VGND.n1088 70.5775
R2081 VGND.n1929 VGND.n1087 70.5775
R2082 VGND.n1616 VGND.n1579 70.5775
R2083 VGND.n1610 VGND.n1569 70.5775
R2084 VGND.n1606 VGND.n1570 70.5775
R2085 VGND.n1602 VGND.n1571 70.5775
R2086 VGND.n1598 VGND.n1572 70.5775
R2087 VGND.n1594 VGND.n1573 70.5775
R2088 VGND.n1590 VGND.n1574 70.5775
R2089 VGND.n1586 VGND.n1575 70.5775
R2090 VGND.n1582 VGND.n1576 70.5775
R2091 VGND.n1577 VGND.n1568 70.5775
R2092 VGND.n2435 VGND.n710 70.5775
R2093 VGND.n2429 VGND.n699 70.5775
R2094 VGND.n2425 VGND.n700 70.5775
R2095 VGND.n2421 VGND.n701 70.5775
R2096 VGND.n2417 VGND.n702 70.5775
R2097 VGND.n2413 VGND.n703 70.5775
R2098 VGND.n2409 VGND.n704 70.5775
R2099 VGND.n2405 VGND.n705 70.5775
R2100 VGND.n2401 VGND.n706 70.5775
R2101 VGND.n2397 VGND.n707 70.5775
R2102 VGND.n2333 VGND.n759 70.5775
R2103 VGND.n2367 VGND.n760 70.5775
R2104 VGND.n2363 VGND.n761 70.5775
R2105 VGND.n2359 VGND.n762 70.5775
R2106 VGND.n2355 VGND.n763 70.5775
R2107 VGND.n2351 VGND.n764 70.5775
R2108 VGND.n2347 VGND.n765 70.5775
R2109 VGND.n2343 VGND.n766 70.5775
R2110 VGND.n2339 VGND.n767 70.5775
R2111 VGND.n2335 VGND.n768 70.5775
R2112 VGND.n2368 VGND.n759 70.5775
R2113 VGND.n2364 VGND.n760 70.5775
R2114 VGND.n2360 VGND.n761 70.5775
R2115 VGND.n2356 VGND.n762 70.5775
R2116 VGND.n2352 VGND.n763 70.5775
R2117 VGND.n2348 VGND.n764 70.5775
R2118 VGND.n2344 VGND.n765 70.5775
R2119 VGND.n2340 VGND.n766 70.5775
R2120 VGND.n2336 VGND.n767 70.5775
R2121 VGND.n768 VGND.n758 70.5775
R2122 VGND.n2195 VGND.n50 70.5775
R2123 VGND.n2191 VGND.n51 70.5775
R2124 VGND.n2187 VGND.n52 70.5775
R2125 VGND.n2183 VGND.n53 70.5775
R2126 VGND.n2179 VGND.n54 70.5775
R2127 VGND.n2175 VGND.n55 70.5775
R2128 VGND.n2171 VGND.n56 70.5775
R2129 VGND.n2167 VGND.n57 70.5775
R2130 VGND.n2163 VGND.n58 70.5775
R2131 VGND.n2159 VGND.n59 70.5775
R2132 VGND.n2155 VGND.n60 70.5775
R2133 VGND.n2151 VGND.n61 70.5775
R2134 VGND.n2147 VGND.n62 70.5775
R2135 VGND.n2143 VGND.n63 70.5775
R2136 VGND.n2139 VGND.n64 70.5775
R2137 VGND.n2135 VGND.n65 70.5775
R2138 VGND.n2131 VGND.n66 70.5775
R2139 VGND.n2127 VGND.n67 70.5775
R2140 VGND.n2123 VGND.n68 70.5775
R2141 VGND.n2119 VGND.n69 70.5775
R2142 VGND.n2115 VGND.n70 70.5775
R2143 VGND.n2111 VGND.n71 70.5775
R2144 VGND.n2107 VGND.n72 70.5775
R2145 VGND.n2103 VGND.n73 70.5775
R2146 VGND.n2099 VGND.n74 70.5775
R2147 VGND.n2095 VGND.n75 70.5775
R2148 VGND.n2091 VGND.n76 70.5775
R2149 VGND.n2087 VGND.n77 70.5775
R2150 VGND.n2083 VGND.n78 70.5775
R2151 VGND.n79 VGND.n49 70.5775
R2152 VGND.n2441 VGND.n542 70.5775
R2153 VGND.n2439 VGND.n544 70.5775
R2154 VGND.n555 VGND.n545 70.5775
R2155 VGND.n559 VGND.n546 70.5775
R2156 VGND.n563 VGND.n547 70.5775
R2157 VGND.n567 VGND.n548 70.5775
R2158 VGND.n550 VGND.n549 70.5775
R2159 VGND.n2499 VGND.n540 70.5775
R2160 VGND.n2491 VGND.n532 70.5775
R2161 VGND.n2487 VGND.n533 70.5775
R2162 VGND.n2483 VGND.n534 70.5775
R2163 VGND.n2479 VGND.n535 70.5775
R2164 VGND.n2475 VGND.n536 70.5775
R2165 VGND.n2471 VGND.n537 70.5775
R2166 VGND.n2467 VGND.n538 70.5775
R2167 VGND.n665 VGND.n583 70.5775
R2168 VGND.n614 VGND.n574 70.5775
R2169 VGND.n618 VGND.n575 70.5775
R2170 VGND.n622 VGND.n576 70.5775
R2171 VGND.n626 VGND.n577 70.5775
R2172 VGND.n630 VGND.n578 70.5775
R2173 VGND.n634 VGND.n579 70.5775
R2174 VGND.n638 VGND.n580 70.5775
R2175 VGND.n642 VGND.n641 60.9887
R2176 VGND.n612 VGND.n611 60.9887
R2177 VGND.n2729 VGND.n47 60.9887
R2178 VGND.n2374 VGND.n756 60.9887
R2179 VGND.n1394 VGND.n1393 60.9887
R2180 VGND.n2396 VGND.n2395 60.9887
R2181 VGND.n1274 VGND.n1202 60.9887
R2182 VGND.n1903 VGND.n1443 60.9887
R2183 VGND.n1646 VGND.n1645 60.9887
R2184 VGND.n1783 VGND 60.9887
R2185 VGND VGND.n1782 60.9887
R2186 VGND.n2031 VGND.n2030 60.9887
R2187 VGND.n1031 VGND.n1030 60.9887
R2188 VGND.n1928 VGND 60.9887
R2189 VGND VGND.n1927 60.9887
R2190 VGND.n2198 VGND.n2197 60.9887
R2191 VGND.n664 VGND.n663 60.9887
R2192 VGND.n2285 VGND 57.4162
R2193 VGND.n1046 VGND 46.7832
R2194 VGND.n1049 VGND 46.7832
R2195 VGND.n1063 VGND 46.7832
R2196 VGND.n1058 VGND 46.7832
R2197 VGND.n1053 VGND 46.7832
R2198 VGND.n1071 VGND 46.0805
R2199 VGND.n1070 VGND.n1069 42.2405
R2200 VGND.n2498 VGND 40.6593
R2201 VGND VGND.n2502 40.6593
R2202 VGND.n2466 VGND 40.6593
R2203 VGND.n1393 VGND 40.6593
R2204 VGND.n2396 VGND 40.6593
R2205 VGND.n1274 VGND 40.6593
R2206 VGND VGND.n1903 40.6593
R2207 VGND VGND.n1646 40.6593
R2208 VGND VGND.n1987 40.6593
R2209 VGND.n2030 VGND 40.6593
R2210 VGND VGND.n2374 40.6593
R2211 VGND VGND.n2729 40.6593
R2212 VGND.n2290 VGND 40.6593
R2213 VGND.n2197 VGND 40.6593
R2214 VGND.n2723 VGND 40.6593
R2215 VGND.n2603 VGND 40.6593
R2216 VGND.n2454 VGND.t301 38.8894
R2217 VGND.n2454 VGND.t303 38.8894
R2218 VGND.n2210 VGND.t510 38.8894
R2219 VGND.n2210 VGND.t515 38.8894
R2220 VGND.n2214 VGND.t26 38.8894
R2221 VGND.n2214 VGND.t29 38.8894
R2222 VGND.n2218 VGND.t401 38.8894
R2223 VGND.n2218 VGND.t445 38.8894
R2224 VGND.n2222 VGND.t468 38.8894
R2225 VGND.n2222 VGND.t470 38.8894
R2226 VGND.n2226 VGND.t498 38.8894
R2227 VGND.n2226 VGND.t500 38.8894
R2228 VGND.n1137 VGND.t10 38.8894
R2229 VGND.n1137 VGND.t464 38.8894
R2230 VGND.n1168 VGND.t524 38.8894
R2231 VGND.n1168 VGND.t525 38.8894
R2232 VGND.n1172 VGND.t344 38.8894
R2233 VGND.n1172 VGND.t342 38.8894
R2234 VGND.n1176 VGND.t338 38.8894
R2235 VGND.n1176 VGND.t340 38.8894
R2236 VGND.n1180 VGND.t473 38.8894
R2237 VGND.n1180 VGND.t472 38.8894
R2238 VGND.n1184 VGND.t321 38.8894
R2239 VGND.n1184 VGND.t320 38.8894
R2240 VGND.n1212 VGND.t511 38.8894
R2241 VGND.n1212 VGND.t518 38.8894
R2242 VGND.n1216 VGND.t532 38.8894
R2243 VGND.n1216 VGND.t534 38.8894
R2244 VGND.n1220 VGND.t489 38.8894
R2245 VGND.n1220 VGND.t486 38.8894
R2246 VGND.n1224 VGND.t326 38.8894
R2247 VGND.n1224 VGND.t327 38.8894
R2248 VGND.n1228 VGND.t312 38.8894
R2249 VGND.n1228 VGND.t309 38.8894
R2250 VGND.n1729 VGND.t502 38.8894
R2251 VGND.n1729 VGND.t503 38.8894
R2252 VGND.n1736 VGND.t286 38.8894
R2253 VGND.n1736 VGND.t287 38.8894
R2254 VGND.n1743 VGND.t289 38.8894
R2255 VGND.n1743 VGND.t291 38.8894
R2256 VGND.n1750 VGND.t441 38.8894
R2257 VGND.n1750 VGND.t438 38.8894
R2258 VGND.n1757 VGND.t351 38.8894
R2259 VGND.n1757 VGND.t442 38.8894
R2260 VGND.n1488 VGND.t517 38.8894
R2261 VGND.n1488 VGND.t505 38.8894
R2262 VGND.n1495 VGND.t403 38.8894
R2263 VGND.n1495 VGND.t402 38.8894
R2264 VGND.n1502 VGND.t335 38.8894
R2265 VGND.n1502 VGND.t333 38.8894
R2266 VGND.n1509 VGND.t420 38.8894
R2267 VGND.n1509 VGND.t421 38.8894
R2268 VGND.n1516 VGND.t162 38.8894
R2269 VGND.n1516 VGND.t159 38.8894
R2270 VGND.n855 VGND.t504 38.8894
R2271 VGND.n855 VGND.t516 38.8894
R2272 VGND.n859 VGND.t389 38.8894
R2273 VGND.n859 VGND.t388 38.8894
R2274 VGND.n863 VGND.t300 38.8894
R2275 VGND.n863 VGND.t297 38.8894
R2276 VGND.n867 VGND.t448 38.8894
R2277 VGND.n867 VGND.t449 38.8894
R2278 VGND.n871 VGND.t424 38.8894
R2279 VGND.n871 VGND.t426 38.8894
R2280 VGND.n2008 VGND.t380 38.8894
R2281 VGND.n2008 VGND.t381 38.8894
R2282 VGND.n2015 VGND.t284 38.8894
R2283 VGND.n2015 VGND.t283 38.8894
R2284 VGND.n21 VGND.t526 38.8894
R2285 VGND.n21 VGND.t519 38.8894
R2286 VGND.n25 VGND.t392 38.8894
R2287 VGND.n25 VGND.t394 38.8894
R2288 VGND.n29 VGND.t397 38.8894
R2289 VGND.n29 VGND.t399 38.8894
R2290 VGND.n33 VGND.t356 38.8894
R2291 VGND.n33 VGND.t354 38.8894
R2292 VGND.n37 VGND.t324 38.8894
R2293 VGND.n37 VGND.t323 38.8894
R2294 VGND.n2552 VGND.t522 38.8894
R2295 VGND.n2552 VGND.t531 38.8894
R2296 VGND.n2559 VGND.t493 38.8894
R2297 VGND.n2559 VGND.t497 38.8894
R2298 VGND.n2566 VGND.t459 38.8894
R2299 VGND.n2566 VGND.t461 38.8894
R2300 VGND.n2573 VGND.t482 38.8894
R2301 VGND.n2573 VGND.t478 38.8894
R2302 VGND.n2580 VGND.t413 38.8894
R2303 VGND.n2580 VGND.t415 38.8894
R2304 VGND.n595 VGND.t407 38.8894
R2305 VGND.n595 VGND.t406 38.8894
R2306 VGND.n2446 VGND.n2445 38.024
R2307 VGND.n2504 VGND.n2503 38.024
R2308 VGND.n2465 VGND.n2464 38.024
R2309 VGND.n1239 VGND.n1238 38.024
R2310 VGND.n1677 VGND.n1676 38.024
R2311 VGND.n1273 VGND.n1272 38.024
R2312 VGND.n1906 VGND.n1904 38.024
R2313 VGND.n1648 VGND.n1647 38.024
R2314 VGND.n1538 VGND.n1537 38.024
R2315 VGND.n1989 VGND.n1988 38.024
R2316 VGND.n2029 VGND.n2028 38.024
R2317 VGND.n1147 VGND.n1146 38.024
R2318 VGND.n2376 VGND.n2375 38.024
R2319 VGND.n2731 VGND.n2730 38.024
R2320 VGND.n2289 VGND.n2288 38.024
R2321 VGND.n2080 VGND.n2079 38.024
R2322 VGND.n2535 VGND.n2534 38.024
R2323 VGND.n2602 VGND.n2601 38.024
R2324 VGND.n2437 VGND.n2436 35.2005
R2325 VGND.n1617 VGND.n667 35.2005
R2326 VGND.n301 VGND 35.171
R2327 VGND.n648 VGND.n646 34.2593
R2328 VGND.n646 VGND.n645 34.2593
R2329 VGND.n610 VGND.n606 34.2593
R2330 VGND.n610 VGND.n609 34.2593
R2331 VGND.n662 VGND.n661 34.2593
R2332 VGND.n2242 VGND.n2240 34.2593
R2333 VGND.n2240 VGND.n2239 34.2593
R2334 VGND.n2201 VGND.n2199 34.2593
R2335 VGND.n833 VGND.n831 34.2593
R2336 VGND.n831 VGND.n830 34.2593
R2337 VGND.n1400 VGND.n1398 34.2593
R2338 VGND.n1398 VGND.n1397 34.2593
R2339 VGND.n1201 VGND.n1200 34.2593
R2340 VGND.n2394 VGND.n711 34.2593
R2341 VGND.n2394 VGND.n2393 34.2593
R2342 VGND.n1201 VGND.n1197 34.2593
R2343 VGND.n1781 VGND.n1780 34.2593
R2344 VGND.n1712 VGND.n1710 34.2593
R2345 VGND.n1710 VGND.n1709 34.2593
R2346 VGND.n1644 VGND.n1619 34.2593
R2347 VGND.n1644 VGND.n1643 34.2593
R2348 VGND.n1781 VGND.n1539 34.2593
R2349 VGND.n2037 VGND.n2035 34.2593
R2350 VGND.n2035 VGND.n2034 34.2593
R2351 VGND.n1029 VGND.n1028 34.2593
R2352 VGND.n1029 VGND.n1025 34.2593
R2353 VGND.n1926 VGND.n1925 34.2593
R2354 VGND.n1926 VGND.n1099 34.2593
R2355 VGND.n2199 VGND.n2078 34.2593
R2356 VGND.n662 VGND.n584 34.2593
R2357 VGND.n1069 VGND 32.8538
R2358 VGND.n1069 VGND 32.8538
R2359 VGND.n2372 VGND.n81 31.26
R2360 VGND.n405 VGND 28.2358
R2361 VGND.n2464 VGND 26.7299
R2362 VGND VGND.n2446 26.7299
R2363 VGND.n2446 VGND 26.7299
R2364 VGND VGND.n2504 26.7299
R2365 VGND.n2504 VGND 26.7299
R2366 VGND.n2464 VGND 26.7299
R2367 VGND.n2601 VGND 26.7299
R2368 VGND.n2376 VGND 26.7299
R2369 VGND VGND.n1147 26.7299
R2370 VGND.n2028 VGND 26.7299
R2371 VGND VGND.n1677 26.7299
R2372 VGND.n1272 VGND 26.7299
R2373 VGND.n1272 VGND 26.7299
R2374 VGND VGND.n1239 26.7299
R2375 VGND.n1239 VGND 26.7299
R2376 VGND.n1677 VGND 26.7299
R2377 VGND VGND.n1648 26.7299
R2378 VGND VGND.n1906 26.7299
R2379 VGND.n1906 VGND 26.7299
R2380 VGND.n1537 VGND 26.7299
R2381 VGND.n1537 VGND 26.7299
R2382 VGND.n1648 VGND 26.7299
R2383 VGND VGND.n1989 26.7299
R2384 VGND.n1989 VGND 26.7299
R2385 VGND.n2028 VGND 26.7299
R2386 VGND.n1147 VGND 26.7299
R2387 VGND VGND.n2376 26.7299
R2388 VGND.n2079 VGND 26.7299
R2389 VGND.n2079 VGND 26.7299
R2390 VGND VGND.n2731 26.7299
R2391 VGND.n2731 VGND 26.7299
R2392 VGND.n2288 VGND 26.7299
R2393 VGND.n2288 VGND 26.7299
R2394 VGND VGND.n2535 26.7299
R2395 VGND.n2535 VGND 26.7299
R2396 VGND.n2601 VGND 26.7299
R2397 VGND VGND.n1070 23.0405
R2398 VGND VGND.n642 20.3299
R2399 VGND.n611 VGND 20.3299
R2400 VGND.n2445 VGND 20.3299
R2401 VGND.n2503 VGND 20.3299
R2402 VGND VGND.n2465 20.3299
R2403 VGND VGND.n47 20.3299
R2404 VGND VGND.n756 20.3299
R2405 VGND VGND.n1394 20.3299
R2406 VGND.n1238 VGND 20.3299
R2407 VGND.n1676 VGND 20.3299
R2408 VGND.n2395 VGND 20.3299
R2409 VGND.n1202 VGND 20.3299
R2410 VGND VGND.n1273 20.3299
R2411 VGND VGND.n1443 20.3299
R2412 VGND.n1904 VGND 20.3299
R2413 VGND.n1647 VGND 20.3299
R2414 VGND.n1645 VGND 20.3299
R2415 VGND VGND.n1538 20.3299
R2416 VGND.n1783 VGND 20.3299
R2417 VGND.n1782 VGND 20.3299
R2418 VGND VGND.n2031 20.3299
R2419 VGND.n1030 VGND 20.3299
R2420 VGND.n1988 VGND 20.3299
R2421 VGND VGND.n2029 20.3299
R2422 VGND.n1146 VGND 20.3299
R2423 VGND.n1928 VGND 20.3299
R2424 VGND.n1927 VGND 20.3299
R2425 VGND.n2375 VGND 20.3299
R2426 VGND.n2730 VGND 20.3299
R2427 VGND VGND.n2289 20.3299
R2428 VGND VGND.n2198 20.3299
R2429 VGND VGND.n2080 20.3299
R2430 VGND.n2534 VGND 20.3299
R2431 VGND VGND.n2602 20.3299
R2432 VGND.n663 VGND 20.3299
R2433 VGND.n2525 VGND 19.0185
R2434 VGND.n646 VGND 17.6946
R2435 VGND VGND.n610 17.6946
R2436 VGND.n2240 VGND 17.6946
R2437 VGND.n831 VGND 17.6946
R2438 VGND.n1398 VGND 17.6946
R2439 VGND VGND.n2394 17.6946
R2440 VGND VGND.n1201 17.6946
R2441 VGND.n1710 VGND 17.6946
R2442 VGND VGND.n1644 17.6946
R2443 VGND VGND.n1781 17.6946
R2444 VGND.n2035 VGND 17.6946
R2445 VGND VGND.n1029 17.6946
R2446 VGND VGND.n1926 17.6946
R2447 VGND.n2199 VGND 17.6946
R2448 VGND VGND.n662 17.6946
R2449 VGND.n2203 VGND 15.2133
R2450 VGND.n2204 VGND 15.2133
R2451 VGND.n2205 VGND 15.2133
R2452 VGND.n2206 VGND 15.2133
R2453 VGND.n2207 VGND 15.2133
R2454 VGND.n2208 VGND 15.2133
R2455 VGND.n2209 VGND 15.2133
R2456 VGND.n2211 VGND 15.2133
R2457 VGND.n2212 VGND 15.2133
R2458 VGND.n2213 VGND 15.2133
R2459 VGND.n2215 VGND 15.2133
R2460 VGND.n2216 VGND 15.2133
R2461 VGND.n2217 VGND 15.2133
R2462 VGND.n2219 VGND 15.2133
R2463 VGND.n2220 VGND 15.2133
R2464 VGND.n2221 VGND 15.2133
R2465 VGND.n2223 VGND 15.2133
R2466 VGND.n2224 VGND 15.2133
R2467 VGND.n2225 VGND 15.2133
R2468 VGND.n2227 VGND 15.2133
R2469 VGND.n2228 VGND 15.2133
R2470 VGND.n2229 VGND 15.2133
R2471 VGND.n2230 VGND 15.2133
R2472 VGND.n2231 VGND 15.2133
R2473 VGND.n2232 VGND 15.2133
R2474 VGND.n2233 VGND 15.2133
R2475 VGND.n2234 VGND 15.2133
R2476 VGND.n810 VGND 15.2133
R2477 VGND.n811 VGND 15.2133
R2478 VGND.n813 VGND 15.2133
R2479 VGND.n815 VGND 15.2133
R2480 VGND.n817 VGND 15.2133
R2481 VGND.n819 VGND 15.2133
R2482 VGND.n821 VGND 15.2133
R2483 VGND.n823 VGND 15.2133
R2484 VGND.n1161 VGND 15.2133
R2485 VGND.n1162 VGND 15.2133
R2486 VGND.n1163 VGND 15.2133
R2487 VGND.n1164 VGND 15.2133
R2488 VGND.n1165 VGND 15.2133
R2489 VGND.n1166 VGND 15.2133
R2490 VGND.n1167 VGND 15.2133
R2491 VGND.n1169 VGND 15.2133
R2492 VGND.n1170 VGND 15.2133
R2493 VGND.n1171 VGND 15.2133
R2494 VGND.n1173 VGND 15.2133
R2495 VGND.n1174 VGND 15.2133
R2496 VGND.n1175 VGND 15.2133
R2497 VGND.n1177 VGND 15.2133
R2498 VGND.n1178 VGND 15.2133
R2499 VGND.n1179 VGND 15.2133
R2500 VGND.n1181 VGND 15.2133
R2501 VGND.n1182 VGND 15.2133
R2502 VGND.n1183 VGND 15.2133
R2503 VGND.n1185 VGND 15.2133
R2504 VGND.n1186 VGND 15.2133
R2505 VGND.n1187 VGND 15.2133
R2506 VGND.n1188 VGND 15.2133
R2507 VGND.n1189 VGND 15.2133
R2508 VGND.n1190 VGND 15.2133
R2509 VGND.n1191 VGND 15.2133
R2510 VGND.n1192 VGND 15.2133
R2511 VGND.n713 VGND 15.2133
R2512 VGND.n714 VGND 15.2133
R2513 VGND.n716 VGND 15.2133
R2514 VGND.n718 VGND 15.2133
R2515 VGND.n720 VGND 15.2133
R2516 VGND.n722 VGND 15.2133
R2517 VGND.n724 VGND 15.2133
R2518 VGND.n726 VGND 15.2133
R2519 VGND.n1715 VGND 15.2133
R2520 VGND.n1717 VGND 15.2133
R2521 VGND.n1719 VGND 15.2133
R2522 VGND.n1721 VGND 15.2133
R2523 VGND.n1723 VGND 15.2133
R2524 VGND.n1725 VGND 15.2133
R2525 VGND.n1727 VGND 15.2133
R2526 VGND.n1730 VGND 15.2133
R2527 VGND.n1732 VGND 15.2133
R2528 VGND.n1734 VGND 15.2133
R2529 VGND.n1737 VGND 15.2133
R2530 VGND.n1739 VGND 15.2133
R2531 VGND.n1741 VGND 15.2133
R2532 VGND.n1744 VGND 15.2133
R2533 VGND.n1746 VGND 15.2133
R2534 VGND.n1748 VGND 15.2133
R2535 VGND.n1751 VGND 15.2133
R2536 VGND.n1753 VGND 15.2133
R2537 VGND.n1755 VGND 15.2133
R2538 VGND.n1758 VGND 15.2133
R2539 VGND.n1760 VGND 15.2133
R2540 VGND.n1762 VGND 15.2133
R2541 VGND.n1764 VGND 15.2133
R2542 VGND.n1766 VGND 15.2133
R2543 VGND.n1768 VGND 15.2133
R2544 VGND.n1770 VGND 15.2133
R2545 VGND.n1772 VGND 15.2133
R2546 VGND.n1621 VGND 15.2133
R2547 VGND.n1622 VGND 15.2133
R2548 VGND.n1624 VGND 15.2133
R2549 VGND.n1626 VGND 15.2133
R2550 VGND.n1628 VGND 15.2133
R2551 VGND.n1630 VGND 15.2133
R2552 VGND.n1632 VGND 15.2133
R2553 VGND.n1634 VGND 15.2133
R2554 VGND.n848 VGND 15.2133
R2555 VGND.n849 VGND 15.2133
R2556 VGND.n850 VGND 15.2133
R2557 VGND.n851 VGND 15.2133
R2558 VGND.n852 VGND 15.2133
R2559 VGND.n853 VGND 15.2133
R2560 VGND.n854 VGND 15.2133
R2561 VGND.n856 VGND 15.2133
R2562 VGND.n857 VGND 15.2133
R2563 VGND.n858 VGND 15.2133
R2564 VGND.n860 VGND 15.2133
R2565 VGND.n861 VGND 15.2133
R2566 VGND.n862 VGND 15.2133
R2567 VGND.n864 VGND 15.2133
R2568 VGND.n865 VGND 15.2133
R2569 VGND.n866 VGND 15.2133
R2570 VGND.n868 VGND 15.2133
R2571 VGND.n869 VGND 15.2133
R2572 VGND.n870 VGND 15.2133
R2573 VGND.n872 VGND 15.2133
R2574 VGND.n873 VGND 15.2133
R2575 VGND.n874 VGND 15.2133
R2576 VGND.n875 VGND 15.2133
R2577 VGND.n876 VGND 15.2133
R2578 VGND.n877 VGND 15.2133
R2579 VGND.n878 VGND 15.2133
R2580 VGND.n879 VGND 15.2133
R2581 VGND.n1102 VGND 15.2133
R2582 VGND.n1103 VGND 15.2133
R2583 VGND.n1105 VGND 15.2133
R2584 VGND.n1107 VGND 15.2133
R2585 VGND.n1109 VGND 15.2133
R2586 VGND.n1111 VGND 15.2133
R2587 VGND.n1113 VGND 15.2133
R2588 VGND.n1115 VGND 15.2133
R2589 VGND.n590 VGND 15.2133
R2590 VGND.n593 VGND 15.2133
R2591 VGND.n594 VGND 15.2133
R2592 VGND.n596 VGND 15.2133
R2593 VGND.n597 VGND 15.2133
R2594 VGND.n599 VGND 13.5534
R2595 VGND.n643 VGND 13.5534
R2596 VGND.n604 VGND 13.5534
R2597 VGND.n607 VGND 13.5534
R2598 VGND.n586 VGND 13.5534
R2599 VGND.n2236 VGND 13.5534
R2600 VGND.n2237 VGND 13.5534
R2601 VGND.n2075 VGND 13.5534
R2602 VGND.n826 VGND 13.5534
R2603 VGND.n828 VGND 13.5534
R2604 VGND.n1194 VGND 13.5534
R2605 VGND.n1395 VGND 13.5534
R2606 VGND.n1198 VGND 13.5534
R2607 VGND.n729 VGND 13.5534
R2608 VGND.n2391 VGND 13.5534
R2609 VGND.n1195 VGND 13.5534
R2610 VGND.n1541 VGND 13.5534
R2611 VGND.n1705 VGND 13.5534
R2612 VGND.n1707 VGND 13.5534
R2613 VGND.n1637 VGND 13.5534
R2614 VGND.n1641 VGND 13.5534
R2615 VGND.n1775 VGND 13.5534
R2616 VGND.n881 VGND 13.5534
R2617 VGND.n2032 VGND 13.5534
R2618 VGND.n1026 VGND 13.5534
R2619 VGND.n1023 VGND 13.5534
R2620 VGND.n1101 VGND 13.5534
R2621 VGND.n1118 VGND 13.5534
R2622 VGND.n2076 VGND 13.5534
R2623 VGND.n588 VGND 13.5534
R2624 VGND.n1048 VGND.n1047 12.8005
R2625 VGND.n648 VGND.n647 12.8005
R2626 VGND.n645 VGND.n644 12.8005
R2627 VGND.n606 VGND.n605 12.8005
R2628 VGND.n609 VGND.n608 12.8005
R2629 VGND.n661 VGND.n585 12.8005
R2630 VGND.n527 VGND 12.8005
R2631 VGND.n2242 VGND.n2241 12.8005
R2632 VGND.n2239 VGND.n2238 12.8005
R2633 VGND.n2201 VGND.n2200 12.8005
R2634 VGND.n833 VGND.n832 12.8005
R2635 VGND.n830 VGND.n827 12.8005
R2636 VGND.n1400 VGND.n1399 12.8005
R2637 VGND.n1397 VGND.n1396 12.8005
R2638 VGND.n1200 VGND.n1199 12.8005
R2639 VGND.n728 VGND.n711 12.8005
R2640 VGND.n2393 VGND.n712 12.8005
R2641 VGND.n1197 VGND.n1196 12.8005
R2642 VGND.n1780 VGND.n1540 12.8005
R2643 VGND.n1712 VGND.n1711 12.8005
R2644 VGND.n1709 VGND.n1706 12.8005
R2645 VGND.n1636 VGND.n1619 12.8005
R2646 VGND.n1643 VGND.n1620 12.8005
R2647 VGND.n1774 VGND.n1539 12.8005
R2648 VGND.n2037 VGND.n2036 12.8005
R2649 VGND.n2034 VGND.n2033 12.8005
R2650 VGND.n1028 VGND.n1027 12.8005
R2651 VGND.n1025 VGND.n1024 12.8005
R2652 VGND.n1925 VGND.n1100 12.8005
R2653 VGND.n1117 VGND.n1099 12.8005
R2654 VGND.n2078 VGND.n2077 12.8005
R2655 VGND.n587 VGND.n584 12.8005
R2656 VGND.n1068 VGND.n1045 12.8005
R2657 VGND.n1062 VGND.n1061 12.8005
R2658 VGND.n1057 VGND.n1056 12.8005
R2659 VGND.n1052 VGND.n1051 12.8005
R2660 VGND.n2451 VGND 10.6647
R2661 VGND.n2447 VGND 10.6647
R2662 VGND VGND.n2444 10.6647
R2663 VGND.n2505 VGND 10.6647
R2664 VGND VGND.n529 10.6647
R2665 VGND VGND.n2463 10.6647
R2666 VGND.n2449 VGND 10.6647
R2667 VGND.n2452 VGND 10.6647
R2668 VGND.n2453 VGND 10.6647
R2669 VGND.n2455 VGND 10.6647
R2670 VGND.n2456 VGND 10.6647
R2671 VGND.n2597 VGND 10.6647
R2672 VGND.n739 VGND 10.6647
R2673 VGND.n740 VGND 10.6647
R2674 VGND.n742 VGND 10.6647
R2675 VGND.n744 VGND 10.6647
R2676 VGND.n746 VGND 10.6647
R2677 VGND.n748 VGND 10.6647
R2678 VGND.n750 VGND 10.6647
R2679 VGND.n752 VGND 10.6647
R2680 VGND VGND.n755 10.6647
R2681 VGND.n1124 VGND 10.6647
R2682 VGND.n1125 VGND 10.6647
R2683 VGND.n1127 VGND 10.6647
R2684 VGND.n1129 VGND 10.6647
R2685 VGND.n1131 VGND 10.6647
R2686 VGND.n1133 VGND 10.6647
R2687 VGND.n1135 VGND 10.6647
R2688 VGND.n1138 VGND 10.6647
R2689 VGND.n1140 VGND 10.6647
R2690 VGND.n1142 VGND 10.6647
R2691 VGND.n1148 VGND 10.6647
R2692 VGND.n2024 VGND 10.6647
R2693 VGND.n1659 VGND 10.6647
R2694 VGND.n1660 VGND 10.6647
R2695 VGND.n1662 VGND 10.6647
R2696 VGND.n1664 VGND 10.6647
R2697 VGND.n1666 VGND 10.6647
R2698 VGND.n1668 VGND 10.6647
R2699 VGND.n1670 VGND 10.6647
R2700 VGND.n1672 VGND 10.6647
R2701 VGND.n1678 VGND 10.6647
R2702 VGND.n1203 VGND 10.6647
R2703 VGND VGND.n1271 10.6647
R2704 VGND.n1240 VGND 10.6647
R2705 VGND VGND.n1237 10.6647
R2706 VGND.n1205 VGND 10.6647
R2707 VGND.n1206 VGND 10.6647
R2708 VGND.n1207 VGND 10.6647
R2709 VGND.n1208 VGND 10.6647
R2710 VGND.n1209 VGND 10.6647
R2711 VGND.n1210 VGND 10.6647
R2712 VGND.n1211 VGND 10.6647
R2713 VGND.n1213 VGND 10.6647
R2714 VGND.n1214 VGND 10.6647
R2715 VGND.n1215 VGND 10.6647
R2716 VGND.n1217 VGND 10.6647
R2717 VGND.n1218 VGND 10.6647
R2718 VGND.n1219 VGND 10.6647
R2719 VGND.n1221 VGND 10.6647
R2720 VGND.n1222 VGND 10.6647
R2721 VGND.n1223 VGND 10.6647
R2722 VGND.n1225 VGND 10.6647
R2723 VGND.n1226 VGND 10.6647
R2724 VGND.n1227 VGND 10.6647
R2725 VGND.n1229 VGND 10.6647
R2726 VGND.n1230 VGND 10.6647
R2727 VGND.n1231 VGND 10.6647
R2728 VGND.n1232 VGND 10.6647
R2729 VGND.n1233 VGND 10.6647
R2730 VGND.n1234 VGND 10.6647
R2731 VGND.n1235 VGND 10.6647
R2732 VGND.n1236 VGND 10.6647
R2733 VGND VGND.n1675 10.6647
R2734 VGND.n1550 VGND 10.6647
R2735 VGND.n1551 VGND 10.6647
R2736 VGND.n1553 VGND 10.6647
R2737 VGND.n1555 VGND 10.6647
R2738 VGND.n1557 VGND 10.6647
R2739 VGND.n1559 VGND 10.6647
R2740 VGND.n1561 VGND 10.6647
R2741 VGND.n1563 VGND 10.6647
R2742 VGND.n1649 VGND 10.6647
R2743 VGND.n1907 VGND 10.6647
R2744 VGND VGND.n1905 10.6647
R2745 VGND.n1533 VGND 10.6647
R2746 VGND VGND.n1536 10.6647
R2747 VGND.n1474 VGND 10.6647
R2748 VGND.n1476 VGND 10.6647
R2749 VGND.n1478 VGND 10.6647
R2750 VGND.n1480 VGND 10.6647
R2751 VGND.n1482 VGND 10.6647
R2752 VGND.n1484 VGND 10.6647
R2753 VGND.n1486 VGND 10.6647
R2754 VGND.n1489 VGND 10.6647
R2755 VGND.n1491 VGND 10.6647
R2756 VGND.n1493 VGND 10.6647
R2757 VGND.n1496 VGND 10.6647
R2758 VGND.n1498 VGND 10.6647
R2759 VGND.n1500 VGND 10.6647
R2760 VGND.n1503 VGND 10.6647
R2761 VGND.n1505 VGND 10.6647
R2762 VGND.n1507 VGND 10.6647
R2763 VGND.n1510 VGND 10.6647
R2764 VGND.n1512 VGND 10.6647
R2765 VGND.n1514 VGND 10.6647
R2766 VGND.n1517 VGND 10.6647
R2767 VGND.n1519 VGND 10.6647
R2768 VGND.n1521 VGND 10.6647
R2769 VGND.n1523 VGND 10.6647
R2770 VGND.n1525 VGND 10.6647
R2771 VGND.n1527 VGND 10.6647
R2772 VGND.n1529 VGND 10.6647
R2773 VGND.n1531 VGND 10.6647
R2774 VGND VGND.n1566 10.6647
R2775 VGND.n1990 VGND 10.6647
R2776 VGND VGND.n884 10.6647
R2777 VGND VGND.n2027 10.6647
R2778 VGND.n1992 VGND 10.6647
R2779 VGND.n1994 VGND 10.6647
R2780 VGND.n1996 VGND 10.6647
R2781 VGND.n1998 VGND 10.6647
R2782 VGND.n2000 VGND 10.6647
R2783 VGND.n2002 VGND 10.6647
R2784 VGND.n2004 VGND 10.6647
R2785 VGND.n2006 VGND 10.6647
R2786 VGND.n2009 VGND 10.6647
R2787 VGND.n2011 VGND 10.6647
R2788 VGND.n2013 VGND 10.6647
R2789 VGND.n2016 VGND 10.6647
R2790 VGND.n2018 VGND 10.6647
R2791 VGND.n2020 VGND 10.6647
R2792 VGND.n2022 VGND 10.6647
R2793 VGND VGND.n1145 10.6647
R2794 VGND.n2377 VGND 10.6647
R2795 VGND VGND.n12 10.6647
R2796 VGND VGND.n13 10.6647
R2797 VGND.n2732 VGND 10.6647
R2798 VGND VGND.n46 10.6647
R2799 VGND.n14 VGND 10.6647
R2800 VGND.n15 VGND 10.6647
R2801 VGND.n16 VGND 10.6647
R2802 VGND.n17 VGND 10.6647
R2803 VGND.n18 VGND 10.6647
R2804 VGND.n19 VGND 10.6647
R2805 VGND.n20 VGND 10.6647
R2806 VGND.n22 VGND 10.6647
R2807 VGND.n23 VGND 10.6647
R2808 VGND.n24 VGND 10.6647
R2809 VGND.n26 VGND 10.6647
R2810 VGND.n27 VGND 10.6647
R2811 VGND.n28 VGND 10.6647
R2812 VGND.n30 VGND 10.6647
R2813 VGND.n31 VGND 10.6647
R2814 VGND.n32 VGND 10.6647
R2815 VGND.n34 VGND 10.6647
R2816 VGND.n35 VGND 10.6647
R2817 VGND.n36 VGND 10.6647
R2818 VGND.n38 VGND 10.6647
R2819 VGND.n39 VGND 10.6647
R2820 VGND.n40 VGND 10.6647
R2821 VGND.n41 VGND 10.6647
R2822 VGND.n42 VGND 10.6647
R2823 VGND.n43 VGND 10.6647
R2824 VGND.n44 VGND 10.6647
R2825 VGND.n45 VGND 10.6647
R2826 VGND.n790 VGND 10.6647
R2827 VGND.n791 VGND 10.6647
R2828 VGND.n793 VGND 10.6647
R2829 VGND.n795 VGND 10.6647
R2830 VGND.n797 VGND 10.6647
R2831 VGND.n799 VGND 10.6647
R2832 VGND.n801 VGND 10.6647
R2833 VGND.n803 VGND 10.6647
R2834 VGND.n805 VGND 10.6647
R2835 VGND VGND.n2287 10.6647
R2836 VGND.n2536 VGND 10.6647
R2837 VGND VGND.n2533 10.6647
R2838 VGND VGND.n2600 10.6647
R2839 VGND.n2538 VGND 10.6647
R2840 VGND.n2540 VGND 10.6647
R2841 VGND.n2542 VGND 10.6647
R2842 VGND.n2544 VGND 10.6647
R2843 VGND.n2546 VGND 10.6647
R2844 VGND.n2548 VGND 10.6647
R2845 VGND.n2550 VGND 10.6647
R2846 VGND.n2553 VGND 10.6647
R2847 VGND.n2555 VGND 10.6647
R2848 VGND.n2557 VGND 10.6647
R2849 VGND.n2560 VGND 10.6647
R2850 VGND.n2562 VGND 10.6647
R2851 VGND.n2564 VGND 10.6647
R2852 VGND.n2567 VGND 10.6647
R2853 VGND.n2569 VGND 10.6647
R2854 VGND.n2571 VGND 10.6647
R2855 VGND.n2574 VGND 10.6647
R2856 VGND.n2576 VGND 10.6647
R2857 VGND.n2578 VGND 10.6647
R2858 VGND.n2581 VGND 10.6647
R2859 VGND.n2583 VGND 10.6647
R2860 VGND.n2585 VGND 10.6647
R2861 VGND.n2587 VGND 10.6647
R2862 VGND.n2589 VGND 10.6647
R2863 VGND.n2591 VGND 10.6647
R2864 VGND.n2593 VGND 10.6647
R2865 VGND.n2595 VGND 10.6647
R2866 VGND.n2496 VGND.n2495 10.4301
R2867 VGND.n2494 VGND.n2492 10.4301
R2868 VGND.n2489 VGND.n2488 10.4301
R2869 VGND.n2485 VGND.n2484 10.4301
R2870 VGND.n2480 VGND.n2477 10.4301
R2871 VGND.n2472 VGND.n2469 10.4301
R2872 VGND.n2468 VGND.n530 10.4301
R2873 VGND.n2434 VGND.n2433 10.4301
R2874 VGND.n2430 VGND.n2427 10.4301
R2875 VGND.n2423 VGND.n2422 10.4301
R2876 VGND.n2419 VGND.n2418 10.4301
R2877 VGND.n2414 VGND.n2411 10.4301
R2878 VGND.n2407 VGND.n2406 10.4301
R2879 VGND.n2403 VGND.n2402 10.4301
R2880 VGND.n2399 VGND.n2398 10.4301
R2881 VGND.n1278 VGND.n1275 10.4301
R2882 VGND.n1282 VGND.n1279 10.4301
R2883 VGND.n1287 VGND.n1286 10.4301
R2884 VGND.n1291 VGND.n1290 10.4301
R2885 VGND.n1298 VGND.n1295 10.4301
R2886 VGND.n1302 VGND.n1299 10.4301
R2887 VGND.n1306 VGND.n1303 10.4301
R2888 VGND.n1315 VGND.n1314 10.4301
R2889 VGND.n1326 VGND.n1323 10.4301
R2890 VGND.n1335 VGND.n1334 10.4301
R2891 VGND.n1346 VGND.n1343 10.4301
R2892 VGND.n1355 VGND.n1354 10.4301
R2893 VGND.n1363 VGND.n1362 10.4301
R2894 VGND.n1371 VGND.n1370 10.4301
R2895 VGND.n1375 VGND.n1374 10.4301
R2896 VGND.n1379 VGND.n1378 10.4301
R2897 VGND.n1383 VGND.n1382 10.4301
R2898 VGND.n1387 VGND.n1386 10.4301
R2899 VGND.n1392 VGND.n1390 10.4301
R2900 VGND.n1615 VGND.n1614 10.4301
R2901 VGND.n1611 VGND.n1608 10.4301
R2902 VGND.n1604 VGND.n1603 10.4301
R2903 VGND.n1600 VGND.n1599 10.4301
R2904 VGND.n1595 VGND.n1592 10.4301
R2905 VGND.n1588 VGND.n1587 10.4301
R2906 VGND.n1584 VGND.n1583 10.4301
R2907 VGND.n1580 VGND.n1567 10.4301
R2908 VGND.n1902 VGND.n1445 10.4301
R2909 VGND.n1897 VGND.n1896 10.4301
R2910 VGND.n1891 VGND.n1890 10.4301
R2911 VGND.n1887 VGND.n1886 10.4301
R2912 VGND.n1882 VGND.n1450 10.4301
R2913 VGND.n1877 VGND.n1876 10.4301
R2914 VGND.n1875 VGND.n1452 10.4301
R2915 VGND.n1863 VGND.n1862 10.4301
R2916 VGND.n1854 VGND.n1457 10.4301
R2917 VGND.n1843 VGND.n1842 10.4301
R2918 VGND.n1834 VGND.n1462 10.4301
R2919 VGND.n1823 VGND.n1822 10.4301
R2920 VGND.n1815 VGND.n1814 10.4301
R2921 VGND.n1807 VGND.n1806 10.4301
R2922 VGND.n1803 VGND.n1802 10.4301
R2923 VGND.n1799 VGND.n1798 10.4301
R2924 VGND.n1795 VGND.n1794 10.4301
R2925 VGND.n1791 VGND.n1790 10.4301
R2926 VGND.n1787 VGND.n1786 10.4301
R2927 VGND.n1978 VGND.n1977 10.4301
R2928 VGND.n1980 VGND.n1979 10.4301
R2929 VGND.n1986 VGND.n886 10.4301
R2930 VGND.n918 VGND.n917 10.4301
R2931 VGND.n925 VGND.n922 10.4301
R2932 VGND.n1002 VGND.n1001 10.4301
R2933 VGND.n1015 VGND.n882 10.4301
R2934 VGND.n1955 VGND.n1954 10.4301
R2935 VGND.n1951 VGND.n1950 10.4301
R2936 VGND.n1946 VGND.n1943 10.4301
R2937 VGND.n1939 VGND.n1938 10.4301
R2938 VGND.n1935 VGND.n1934 10.4301
R2939 VGND.n1931 VGND.n1930 10.4301
R2940 VGND.n2370 VGND.n2369 10.4301
R2941 VGND.n2365 VGND.n2362 10.4301
R2942 VGND.n2358 VGND.n2357 10.4301
R2943 VGND.n2354 VGND.n2353 10.4301
R2944 VGND.n2349 VGND.n2346 10.4301
R2945 VGND.n2342 VGND.n2341 10.4301
R2946 VGND.n2338 VGND.n2337 10.4301
R2947 VGND.n2334 VGND.n757 10.4301
R2948 VGND.n2330 VGND.n2329 10.4301
R2949 VGND.n2323 VGND.n2322 10.4301
R2950 VGND.n2315 VGND.n777 10.4301
R2951 VGND.n2314 VGND.n2313 10.4301
R2952 VGND.n2307 VGND.n2306 10.4301
R2953 VGND.n2299 VGND.n785 10.4301
R2954 VGND.n2298 VGND.n2297 10.4301
R2955 VGND.n2291 VGND.n789 10.4301
R2956 VGND.n2196 VGND.n2193 10.4301
R2957 VGND.n2192 VGND.n2189 10.4301
R2958 VGND.n2185 VGND.n2184 10.4301
R2959 VGND.n2181 VGND.n2180 10.4301
R2960 VGND.n2176 VGND.n2173 10.4301
R2961 VGND.n2172 VGND.n2169 10.4301
R2962 VGND.n2168 VGND.n2165 10.4301
R2963 VGND.n2157 VGND.n2156 10.4301
R2964 VGND.n2148 VGND.n2145 10.4301
R2965 VGND.n2137 VGND.n2136 10.4301
R2966 VGND.n2128 VGND.n2125 10.4301
R2967 VGND.n2117 VGND.n2116 10.4301
R2968 VGND.n2109 VGND.n2108 10.4301
R2969 VGND.n2101 VGND.n2100 10.4301
R2970 VGND.n2097 VGND.n2096 10.4301
R2971 VGND.n2093 VGND.n2092 10.4301
R2972 VGND.n2089 VGND.n2088 10.4301
R2973 VGND.n2085 VGND.n2084 10.4301
R2974 VGND.n2081 VGND.n48 10.4301
R2975 VGND.n2722 VGND.n2721 10.4301
R2976 VGND.n2715 VGND.n87 10.4301
R2977 VGND.n2713 VGND.n88 10.4301
R2978 VGND.n2707 VGND.n2706 10.4301
R2979 VGND.n2699 VGND.n95 10.4301
R2980 VGND.n2698 VGND.n2697 10.4301
R2981 VGND.n2691 VGND.n99 10.4301
R2982 VGND.n2683 VGND.n2682 10.4301
R2983 VGND.n2674 VGND.n2673 10.4301
R2984 VGND.n2665 VGND.n112 10.4301
R2985 VGND.n2651 VGND.n119 10.4301
R2986 VGND.n2643 VGND.n2642 10.4301
R2987 VGND.n2635 VGND.n2634 10.4301
R2988 VGND.n2627 VGND.n2626 10.4301
R2989 VGND.n2625 VGND.n133 10.4301
R2990 VGND.n2619 VGND.n2618 10.4301
R2991 VGND.n2617 VGND.n137 10.4301
R2992 VGND.n2611 VGND.n2610 10.4301
R2993 VGND.n2609 VGND.n141 10.4301
R2994 VGND.n601 VGND.n600 10.4301
R2995 VGND.n613 VGND.n603 10.4301
R2996 VGND.n617 VGND.n616 10.4301
R2997 VGND.n621 VGND.n620 10.4301
R2998 VGND.n628 VGND.n625 10.4301
R2999 VGND.n636 VGND.n633 10.4301
R3000 VGND.n640 VGND.n637 10.4301
R3001 VGND.n2442 VGND.n543 10.4301
R3002 VGND.n553 VGND.n551 10.4301
R3003 VGND.n557 VGND.n554 10.4301
R3004 VGND.n561 VGND.n558 10.4301
R3005 VGND.n565 VGND.n562 10.4301
R3006 VGND.n569 VGND.n566 10.4301
R3007 VGND.n571 VGND.n570 10.4301
R3008 VGND.n1073 VGND.n1072 10.4301
R3009 VGND.n1079 VGND.n1039 10.4301
R3010 VGND.n1081 VGND.n1080 10.4301
R3011 VGND.n1050 VGND.n1047 9.3947
R3012 VGND.n1068 VGND.n1067 9.3947
R3013 VGND.n1064 VGND.n1061 9.3947
R3014 VGND.n1059 VGND.n1056 9.3947
R3015 VGND.n1054 VGND.n1051 9.3947
R3016 VGND.n649 VGND.n599 9.39464
R3017 VGND.n649 VGND.n648 9.39464
R3018 VGND.n643 VGND.n598 9.39464
R3019 VGND.n645 VGND.n598 9.39464
R3020 VGND.n604 VGND.n592 9.39464
R3021 VGND.n606 VGND.n592 9.39464
R3022 VGND.n607 VGND.n591 9.39464
R3023 VGND.n609 VGND.n591 9.39464
R3024 VGND.n660 VGND.n586 9.39464
R3025 VGND.n661 VGND.n660 9.39464
R3026 VGND.n2243 VGND.n2236 9.39464
R3027 VGND.n2243 VGND.n2242 9.39464
R3028 VGND.n2237 VGND.n2235 9.39464
R3029 VGND.n2239 VGND.n2235 9.39464
R3030 VGND.n2202 VGND.n2075 9.39464
R3031 VGND.n2202 VGND.n2201 9.39464
R3032 VGND.n834 VGND.n826 9.39464
R3033 VGND.n834 VGND.n833 9.39464
R3034 VGND.n829 VGND.n828 9.39464
R3035 VGND.n1401 VGND.n1194 9.39464
R3036 VGND.n1401 VGND.n1400 9.39464
R3037 VGND.n1395 VGND.n1193 9.39464
R3038 VGND.n1397 VGND.n1193 9.39464
R3039 VGND.n1198 VGND.n1160 9.39464
R3040 VGND.n1200 VGND.n1160 9.39464
R3041 VGND.n730 VGND.n729 9.39464
R3042 VGND.n730 VGND.n711 9.39464
R3043 VGND.n2392 VGND.n2391 9.39464
R3044 VGND.n2393 VGND.n2392 9.39464
R3045 VGND.n1197 VGND.n1159 9.39464
R3046 VGND.n1195 VGND.n1159 9.39464
R3047 VGND.n1779 VGND.n1541 9.39464
R3048 VGND.n1780 VGND.n1779 9.39464
R3049 VGND.n1713 VGND.n1705 9.39464
R3050 VGND.n1713 VGND.n1712 9.39464
R3051 VGND.n1708 VGND.n1707 9.39464
R3052 VGND.n1709 VGND.n1708 9.39464
R3053 VGND.n1638 VGND.n1637 9.39464
R3054 VGND.n1638 VGND.n1619 9.39464
R3055 VGND.n1642 VGND.n1641 9.39464
R3056 VGND.n1643 VGND.n1642 9.39464
R3057 VGND.n1776 VGND.n1539 9.39464
R3058 VGND.n1776 VGND.n1775 9.39464
R3059 VGND.n2038 VGND.n881 9.39464
R3060 VGND.n2038 VGND.n2037 9.39464
R3061 VGND.n2032 VGND.n880 9.39464
R3062 VGND.n2034 VGND.n880 9.39464
R3063 VGND.n1026 VGND.n847 9.39464
R3064 VGND.n1028 VGND.n847 9.39464
R3065 VGND.n1025 VGND.n846 9.39464
R3066 VGND.n1023 VGND.n846 9.39464
R3067 VGND.n1924 VGND.n1101 9.39464
R3068 VGND.n1925 VGND.n1924 9.39464
R3069 VGND.n1119 VGND.n1099 9.39464
R3070 VGND.n1119 VGND.n1118 9.39464
R3071 VGND.n830 VGND.n829 9.39464
R3072 VGND.n2078 VGND.n2074 9.39464
R3073 VGND.n2076 VGND.n2074 9.39464
R3074 VGND.n589 VGND.n584 9.39464
R3075 VGND.n589 VGND.n588 9.39464
R3076 VGND.n1050 VGND.n1049 9.39457
R3077 VGND.n1067 VGND.n1046 9.39457
R3078 VGND.n1064 VGND.n1063 9.39457
R3079 VGND.n1059 VGND.n1058 9.39457
R3080 VGND.n1054 VGND.n1053 9.39457
R3081 VGND VGND.n810 9.36745
R3082 VGND VGND.n713 9.36745
R3083 VGND VGND.n1621 9.36745
R3084 VGND VGND.n1102 9.36745
R3085 VGND.n2272 VGND.n2203 9.34497
R3086 VGND.n2271 VGND.n2204 9.34497
R3087 VGND.n2270 VGND.n2205 9.34497
R3088 VGND.n2269 VGND.n2206 9.34497
R3089 VGND.n2268 VGND.n2207 9.34497
R3090 VGND.n2267 VGND.n2208 9.34497
R3091 VGND.n2266 VGND.n2209 9.34497
R3092 VGND.n2265 VGND.n2211 9.34497
R3093 VGND.n2264 VGND.n2212 9.34497
R3094 VGND.n2263 VGND.n2213 9.34497
R3095 VGND.n2262 VGND.n2215 9.34497
R3096 VGND.n2261 VGND.n2216 9.34497
R3097 VGND.n2260 VGND.n2217 9.34497
R3098 VGND.n2259 VGND.n2219 9.34497
R3099 VGND.n2258 VGND.n2220 9.34497
R3100 VGND.n2257 VGND.n2221 9.34497
R3101 VGND.n2256 VGND.n2223 9.34497
R3102 VGND.n2255 VGND.n2224 9.34497
R3103 VGND.n2254 VGND.n2225 9.34497
R3104 VGND.n2253 VGND.n2227 9.34497
R3105 VGND.n2252 VGND.n2228 9.34497
R3106 VGND.n2251 VGND.n2229 9.34497
R3107 VGND.n2250 VGND.n2230 9.34497
R3108 VGND.n2249 VGND.n2231 9.34497
R3109 VGND.n2248 VGND.n2232 9.34497
R3110 VGND.n2247 VGND.n2233 9.34497
R3111 VGND.n2246 VGND.n2234 9.34497
R3112 VGND.n812 VGND.n811 9.34497
R3113 VGND.n814 VGND.n813 9.34497
R3114 VGND.n816 VGND.n815 9.34497
R3115 VGND.n818 VGND.n817 9.34497
R3116 VGND.n820 VGND.n819 9.34497
R3117 VGND.n822 VGND.n821 9.34497
R3118 VGND.n824 VGND.n823 9.34497
R3119 VGND.n1430 VGND.n1161 9.34497
R3120 VGND.n1429 VGND.n1162 9.34497
R3121 VGND.n1428 VGND.n1163 9.34497
R3122 VGND.n1427 VGND.n1164 9.34497
R3123 VGND.n1426 VGND.n1165 9.34497
R3124 VGND.n1425 VGND.n1166 9.34497
R3125 VGND.n1424 VGND.n1167 9.34497
R3126 VGND.n1423 VGND.n1169 9.34497
R3127 VGND.n1422 VGND.n1170 9.34497
R3128 VGND.n1421 VGND.n1171 9.34497
R3129 VGND.n1420 VGND.n1173 9.34497
R3130 VGND.n1419 VGND.n1174 9.34497
R3131 VGND.n1418 VGND.n1175 9.34497
R3132 VGND.n1417 VGND.n1177 9.34497
R3133 VGND.n1416 VGND.n1178 9.34497
R3134 VGND.n1415 VGND.n1179 9.34497
R3135 VGND.n1414 VGND.n1181 9.34497
R3136 VGND.n1413 VGND.n1182 9.34497
R3137 VGND.n1412 VGND.n1183 9.34497
R3138 VGND.n1411 VGND.n1185 9.34497
R3139 VGND.n1410 VGND.n1186 9.34497
R3140 VGND.n1409 VGND.n1187 9.34497
R3141 VGND.n1408 VGND.n1188 9.34497
R3142 VGND.n1407 VGND.n1189 9.34497
R3143 VGND.n1406 VGND.n1190 9.34497
R3144 VGND.n1405 VGND.n1191 9.34497
R3145 VGND.n1404 VGND.n1192 9.34497
R3146 VGND.n715 VGND.n714 9.34497
R3147 VGND.n717 VGND.n716 9.34497
R3148 VGND.n719 VGND.n718 9.34497
R3149 VGND.n721 VGND.n720 9.34497
R3150 VGND.n723 VGND.n722 9.34497
R3151 VGND.n725 VGND.n724 9.34497
R3152 VGND.n727 VGND.n726 9.34497
R3153 VGND.n1716 VGND.n1715 9.34497
R3154 VGND.n1718 VGND.n1717 9.34497
R3155 VGND.n1720 VGND.n1719 9.34497
R3156 VGND.n1722 VGND.n1721 9.34497
R3157 VGND.n1724 VGND.n1723 9.34497
R3158 VGND.n1726 VGND.n1725 9.34497
R3159 VGND.n1728 VGND.n1727 9.34497
R3160 VGND.n1731 VGND.n1730 9.34497
R3161 VGND.n1733 VGND.n1732 9.34497
R3162 VGND.n1735 VGND.n1734 9.34497
R3163 VGND.n1738 VGND.n1737 9.34497
R3164 VGND.n1740 VGND.n1739 9.34497
R3165 VGND.n1742 VGND.n1741 9.34497
R3166 VGND.n1745 VGND.n1744 9.34497
R3167 VGND.n1747 VGND.n1746 9.34497
R3168 VGND.n1749 VGND.n1748 9.34497
R3169 VGND.n1752 VGND.n1751 9.34497
R3170 VGND.n1754 VGND.n1753 9.34497
R3171 VGND.n1756 VGND.n1755 9.34497
R3172 VGND.n1759 VGND.n1758 9.34497
R3173 VGND.n1761 VGND.n1760 9.34497
R3174 VGND.n1763 VGND.n1762 9.34497
R3175 VGND.n1765 VGND.n1764 9.34497
R3176 VGND.n1767 VGND.n1766 9.34497
R3177 VGND.n1769 VGND.n1768 9.34497
R3178 VGND.n1771 VGND.n1770 9.34497
R3179 VGND.n1773 VGND.n1772 9.34497
R3180 VGND.n1623 VGND.n1622 9.34497
R3181 VGND.n1625 VGND.n1624 9.34497
R3182 VGND.n1627 VGND.n1626 9.34497
R3183 VGND.n1629 VGND.n1628 9.34497
R3184 VGND.n1631 VGND.n1630 9.34497
R3185 VGND.n1633 VGND.n1632 9.34497
R3186 VGND.n1635 VGND.n1634 9.34497
R3187 VGND.n2067 VGND.n848 9.34497
R3188 VGND.n2066 VGND.n849 9.34497
R3189 VGND.n2065 VGND.n850 9.34497
R3190 VGND.n2064 VGND.n851 9.34497
R3191 VGND.n2063 VGND.n852 9.34497
R3192 VGND.n2062 VGND.n853 9.34497
R3193 VGND.n2061 VGND.n854 9.34497
R3194 VGND.n2060 VGND.n856 9.34497
R3195 VGND.n2059 VGND.n857 9.34497
R3196 VGND.n2058 VGND.n858 9.34497
R3197 VGND.n2057 VGND.n860 9.34497
R3198 VGND.n2056 VGND.n861 9.34497
R3199 VGND.n2055 VGND.n862 9.34497
R3200 VGND.n2054 VGND.n864 9.34497
R3201 VGND.n2053 VGND.n865 9.34497
R3202 VGND.n2052 VGND.n866 9.34497
R3203 VGND.n2051 VGND.n868 9.34497
R3204 VGND.n2050 VGND.n869 9.34497
R3205 VGND.n2049 VGND.n870 9.34497
R3206 VGND.n2048 VGND.n872 9.34497
R3207 VGND.n2047 VGND.n873 9.34497
R3208 VGND.n2046 VGND.n874 9.34497
R3209 VGND.n2045 VGND.n875 9.34497
R3210 VGND.n2044 VGND.n876 9.34497
R3211 VGND.n2043 VGND.n877 9.34497
R3212 VGND.n2042 VGND.n878 9.34497
R3213 VGND.n2041 VGND.n879 9.34497
R3214 VGND.n1104 VGND.n1103 9.34497
R3215 VGND.n1106 VGND.n1105 9.34497
R3216 VGND.n1108 VGND.n1107 9.34497
R3217 VGND.n1110 VGND.n1109 9.34497
R3218 VGND.n1112 VGND.n1111 9.34497
R3219 VGND.n1114 VGND.n1113 9.34497
R3220 VGND.n1116 VGND.n1115 9.34497
R3221 VGND.n658 VGND.n590 9.34497
R3222 VGND.n655 VGND.n593 9.34497
R3223 VGND.n654 VGND.n594 9.34497
R3224 VGND.n653 VGND.n596 9.34497
R3225 VGND.n652 VGND.n597 9.34497
R3226 VGND.n2527 VGND.n146 9.3005
R3227 VGND.n2529 VGND.n146 9.3005
R3228 VGND.n2277 VGND.n146 9.3005
R3229 VGND.n837 VGND.n146 9.3005
R3230 VGND.n157 VGND.n146 9.3005
R3231 VGND.n1435 VGND.n146 9.3005
R3232 VGND.n1157 VGND.n146 9.3005
R3233 VGND.n1685 VGND.n146 9.3005
R3234 VGND.n1681 VGND.n146 9.3005
R3235 VGND.n1543 VGND.n146 9.3005
R3236 VGND.n1545 VGND.n146 9.3005
R3237 VGND.n1911 VGND.n146 9.3005
R3238 VGND.n1440 VGND.n146 9.3005
R3239 VGND.n841 VGND.n146 9.3005
R3240 VGND.n843 VGND.n146 9.3005
R3241 VGND.n1154 VGND.n146 9.3005
R3242 VGND.n1150 VGND.n146 9.3005
R3243 VGND.n2526 VGND.n157 9.3005
R3244 VGND.n2448 VGND.n2444 7.91498
R3245 VGND VGND.n739 7.89251
R3246 VGND VGND.n1124 7.89251
R3247 VGND VGND.n1659 7.89251
R3248 VGND VGND.n1550 7.89251
R3249 VGND VGND.n790 7.89251
R3250 VGND.n529 VGND.n528 7.87003
R3251 VGND.n2506 VGND.n2505 7.87003
R3252 VGND.n2461 VGND.n2451 7.87003
R3253 VGND.n2448 VGND.n2447 7.87003
R3254 VGND.n755 VGND.n754 7.87003
R3255 VGND.n1241 VGND.n1240 7.87003
R3256 VGND.n1675 VGND.n1674 7.87003
R3257 VGND.n1908 VGND.n1907 7.87003
R3258 VGND.n1566 VGND.n1565 7.87003
R3259 VGND.n884 VGND.n883 7.87003
R3260 VGND.n2025 VGND.n2024 7.87003
R3261 VGND.n1991 VGND.n1990 7.87003
R3262 VGND.n1145 VGND.n1144 7.87003
R3263 VGND.n2733 VGND.n2732 7.87003
R3264 VGND.n806 VGND.n805 7.87003
R3265 VGND.n2533 VGND.n2532 7.87003
R3266 VGND.n2598 VGND.n2597 7.87003
R3267 VGND.n2537 VGND.n2536 7.87003
R3268 VGND.n2463 VGND.n2462 7.87003
R3269 VGND.n2450 VGND.n2449 7.87003
R3270 VGND.n2460 VGND.n2452 7.87003
R3271 VGND.n2459 VGND.n2453 7.87003
R3272 VGND.n2458 VGND.n2455 7.87003
R3273 VGND.n2457 VGND.n2456 7.87003
R3274 VGND.n741 VGND.n740 7.87003
R3275 VGND.n743 VGND.n742 7.87003
R3276 VGND.n745 VGND.n744 7.87003
R3277 VGND.n747 VGND.n746 7.87003
R3278 VGND.n749 VGND.n748 7.87003
R3279 VGND.n751 VGND.n750 7.87003
R3280 VGND.n753 VGND.n752 7.87003
R3281 VGND.n1126 VGND.n1125 7.87003
R3282 VGND.n1128 VGND.n1127 7.87003
R3283 VGND.n1130 VGND.n1129 7.87003
R3284 VGND.n1132 VGND.n1131 7.87003
R3285 VGND.n1134 VGND.n1133 7.87003
R3286 VGND.n1136 VGND.n1135 7.87003
R3287 VGND.n1139 VGND.n1138 7.87003
R3288 VGND.n1141 VGND.n1140 7.87003
R3289 VGND.n1143 VGND.n1142 7.87003
R3290 VGND.n1149 VGND.n1148 7.87003
R3291 VGND.n1661 VGND.n1660 7.87003
R3292 VGND.n1663 VGND.n1662 7.87003
R3293 VGND.n1665 VGND.n1664 7.87003
R3294 VGND.n1667 VGND.n1666 7.87003
R3295 VGND.n1669 VGND.n1668 7.87003
R3296 VGND.n1671 VGND.n1670 7.87003
R3297 VGND.n1673 VGND.n1672 7.87003
R3298 VGND.n1679 VGND.n1678 7.87003
R3299 VGND.n1204 VGND.n1203 7.87003
R3300 VGND.n1271 VGND.n1270 7.87003
R3301 VGND.n1242 VGND.n1237 7.87003
R3302 VGND.n1269 VGND.n1205 7.87003
R3303 VGND.n1268 VGND.n1206 7.87003
R3304 VGND.n1267 VGND.n1207 7.87003
R3305 VGND.n1266 VGND.n1208 7.87003
R3306 VGND.n1265 VGND.n1209 7.87003
R3307 VGND.n1264 VGND.n1210 7.87003
R3308 VGND.n1263 VGND.n1211 7.87003
R3309 VGND.n1262 VGND.n1213 7.87003
R3310 VGND.n1261 VGND.n1214 7.87003
R3311 VGND.n1260 VGND.n1215 7.87003
R3312 VGND.n1259 VGND.n1217 7.87003
R3313 VGND.n1258 VGND.n1218 7.87003
R3314 VGND.n1257 VGND.n1219 7.87003
R3315 VGND.n1256 VGND.n1221 7.87003
R3316 VGND.n1255 VGND.n1222 7.87003
R3317 VGND.n1254 VGND.n1223 7.87003
R3318 VGND.n1253 VGND.n1225 7.87003
R3319 VGND.n1252 VGND.n1226 7.87003
R3320 VGND.n1251 VGND.n1227 7.87003
R3321 VGND.n1250 VGND.n1229 7.87003
R3322 VGND.n1249 VGND.n1230 7.87003
R3323 VGND.n1248 VGND.n1231 7.87003
R3324 VGND.n1247 VGND.n1232 7.87003
R3325 VGND.n1246 VGND.n1233 7.87003
R3326 VGND.n1245 VGND.n1234 7.87003
R3327 VGND.n1244 VGND.n1235 7.87003
R3328 VGND.n1243 VGND.n1236 7.87003
R3329 VGND.n1552 VGND.n1551 7.87003
R3330 VGND.n1554 VGND.n1553 7.87003
R3331 VGND.n1556 VGND.n1555 7.87003
R3332 VGND.n1558 VGND.n1557 7.87003
R3333 VGND.n1560 VGND.n1559 7.87003
R3334 VGND.n1562 VGND.n1561 7.87003
R3335 VGND.n1564 VGND.n1563 7.87003
R3336 VGND.n1650 VGND.n1649 7.87003
R3337 VGND.n1905 VGND.n1442 7.87003
R3338 VGND.n1534 VGND.n1533 7.87003
R3339 VGND.n1536 VGND.n1535 7.87003
R3340 VGND.n1475 VGND.n1474 7.87003
R3341 VGND.n1477 VGND.n1476 7.87003
R3342 VGND.n1479 VGND.n1478 7.87003
R3343 VGND.n1481 VGND.n1480 7.87003
R3344 VGND.n1483 VGND.n1482 7.87003
R3345 VGND.n1485 VGND.n1484 7.87003
R3346 VGND.n1487 VGND.n1486 7.87003
R3347 VGND.n1490 VGND.n1489 7.87003
R3348 VGND.n1492 VGND.n1491 7.87003
R3349 VGND.n1494 VGND.n1493 7.87003
R3350 VGND.n1497 VGND.n1496 7.87003
R3351 VGND.n1499 VGND.n1498 7.87003
R3352 VGND.n1501 VGND.n1500 7.87003
R3353 VGND.n1504 VGND.n1503 7.87003
R3354 VGND.n1506 VGND.n1505 7.87003
R3355 VGND.n1508 VGND.n1507 7.87003
R3356 VGND.n1511 VGND.n1510 7.87003
R3357 VGND.n1513 VGND.n1512 7.87003
R3358 VGND.n1515 VGND.n1514 7.87003
R3359 VGND.n1518 VGND.n1517 7.87003
R3360 VGND.n1520 VGND.n1519 7.87003
R3361 VGND.n1522 VGND.n1521 7.87003
R3362 VGND.n1524 VGND.n1523 7.87003
R3363 VGND.n1526 VGND.n1525 7.87003
R3364 VGND.n1528 VGND.n1527 7.87003
R3365 VGND.n1530 VGND.n1529 7.87003
R3366 VGND.n1532 VGND.n1531 7.87003
R3367 VGND.n2027 VGND.n2026 7.87003
R3368 VGND.n1993 VGND.n1992 7.87003
R3369 VGND.n1995 VGND.n1994 7.87003
R3370 VGND.n1997 VGND.n1996 7.87003
R3371 VGND.n1999 VGND.n1998 7.87003
R3372 VGND.n2001 VGND.n2000 7.87003
R3373 VGND.n2003 VGND.n2002 7.87003
R3374 VGND.n2005 VGND.n2004 7.87003
R3375 VGND.n2007 VGND.n2006 7.87003
R3376 VGND.n2010 VGND.n2009 7.87003
R3377 VGND.n2012 VGND.n2011 7.87003
R3378 VGND.n2014 VGND.n2013 7.87003
R3379 VGND.n2017 VGND.n2016 7.87003
R3380 VGND.n2019 VGND.n2018 7.87003
R3381 VGND.n2021 VGND.n2020 7.87003
R3382 VGND.n2023 VGND.n2022 7.87003
R3383 VGND.n2378 VGND.n2377 7.87003
R3384 VGND.n2763 VGND.n12 7.87003
R3385 VGND.n2762 VGND.n13 7.87003
R3386 VGND.n2734 VGND.n46 7.87003
R3387 VGND.n2761 VGND.n14 7.87003
R3388 VGND.n2760 VGND.n15 7.87003
R3389 VGND.n2759 VGND.n16 7.87003
R3390 VGND.n2758 VGND.n17 7.87003
R3391 VGND.n2757 VGND.n18 7.87003
R3392 VGND.n2756 VGND.n19 7.87003
R3393 VGND.n2755 VGND.n20 7.87003
R3394 VGND.n2754 VGND.n22 7.87003
R3395 VGND.n2753 VGND.n23 7.87003
R3396 VGND.n2752 VGND.n24 7.87003
R3397 VGND.n2751 VGND.n26 7.87003
R3398 VGND.n2750 VGND.n27 7.87003
R3399 VGND.n2749 VGND.n28 7.87003
R3400 VGND.n2748 VGND.n30 7.87003
R3401 VGND.n2747 VGND.n31 7.87003
R3402 VGND.n2746 VGND.n32 7.87003
R3403 VGND.n2745 VGND.n34 7.87003
R3404 VGND.n2744 VGND.n35 7.87003
R3405 VGND.n2743 VGND.n36 7.87003
R3406 VGND.n2742 VGND.n38 7.87003
R3407 VGND.n2741 VGND.n39 7.87003
R3408 VGND.n2740 VGND.n40 7.87003
R3409 VGND.n2739 VGND.n41 7.87003
R3410 VGND.n2738 VGND.n42 7.87003
R3411 VGND.n2737 VGND.n43 7.87003
R3412 VGND.n2736 VGND.n44 7.87003
R3413 VGND.n2735 VGND.n45 7.87003
R3414 VGND.n792 VGND.n791 7.87003
R3415 VGND.n794 VGND.n793 7.87003
R3416 VGND.n796 VGND.n795 7.87003
R3417 VGND.n798 VGND.n797 7.87003
R3418 VGND.n800 VGND.n799 7.87003
R3419 VGND.n802 VGND.n801 7.87003
R3420 VGND.n804 VGND.n803 7.87003
R3421 VGND.n2287 VGND.n2286 7.87003
R3422 VGND.n2600 VGND.n2599 7.87003
R3423 VGND.n2539 VGND.n2538 7.87003
R3424 VGND.n2541 VGND.n2540 7.87003
R3425 VGND.n2543 VGND.n2542 7.87003
R3426 VGND.n2545 VGND.n2544 7.87003
R3427 VGND.n2547 VGND.n2546 7.87003
R3428 VGND.n2549 VGND.n2548 7.87003
R3429 VGND.n2551 VGND.n2550 7.87003
R3430 VGND.n2554 VGND.n2553 7.87003
R3431 VGND.n2556 VGND.n2555 7.87003
R3432 VGND.n2558 VGND.n2557 7.87003
R3433 VGND.n2561 VGND.n2560 7.87003
R3434 VGND.n2563 VGND.n2562 7.87003
R3435 VGND.n2565 VGND.n2564 7.87003
R3436 VGND.n2568 VGND.n2567 7.87003
R3437 VGND.n2570 VGND.n2569 7.87003
R3438 VGND.n2572 VGND.n2571 7.87003
R3439 VGND.n2575 VGND.n2574 7.87003
R3440 VGND.n2577 VGND.n2576 7.87003
R3441 VGND.n2579 VGND.n2578 7.87003
R3442 VGND.n2582 VGND.n2581 7.87003
R3443 VGND.n2584 VGND.n2583 7.87003
R3444 VGND.n2586 VGND.n2585 7.87003
R3445 VGND.n2588 VGND.n2587 7.87003
R3446 VGND.n2590 VGND.n2589 7.87003
R3447 VGND.n2592 VGND.n2591 7.87003
R3448 VGND.n2594 VGND.n2593 7.87003
R3449 VGND.n2596 VGND.n2595 7.87003
R3450 VGND.n2495 VGND 7.82272
R3451 VGND.n2488 VGND 7.82272
R3452 VGND.n2484 VGND 7.82272
R3453 VGND.n2481 VGND 7.82272
R3454 VGND.n2477 VGND 7.82272
R3455 VGND.n2476 VGND 7.82272
R3456 VGND.n2473 VGND 7.82272
R3457 VGND.n2469 VGND 7.82272
R3458 VGND.n2433 VGND 7.82272
R3459 VGND.n2432 VGND 7.82272
R3460 VGND.n2427 VGND 7.82272
R3461 VGND.n2426 VGND 7.82272
R3462 VGND.n2422 VGND 7.82272
R3463 VGND.n2418 VGND 7.82272
R3464 VGND.n2415 VGND 7.82272
R3465 VGND.n2411 VGND 7.82272
R3466 VGND.n2410 VGND 7.82272
R3467 VGND.n2406 VGND 7.82272
R3468 VGND.n2402 VGND 7.82272
R3469 VGND VGND.n1278 7.82272
R3470 VGND VGND.n1282 7.82272
R3471 VGND.n1283 VGND 7.82272
R3472 VGND.n1287 VGND 7.82272
R3473 VGND.n1291 VGND 7.82272
R3474 VGND VGND.n1294 7.82272
R3475 VGND VGND.n1298 7.82272
R3476 VGND VGND.n1302 7.82272
R3477 VGND VGND.n1306 7.82272
R3478 VGND.n1307 VGND 7.82272
R3479 VGND VGND.n1310 7.82272
R3480 VGND.n1311 VGND 7.82272
R3481 VGND.n1315 VGND 7.82272
R3482 VGND VGND.n1318 7.82272
R3483 VGND.n1319 VGND 7.82272
R3484 VGND VGND.n1322 7.82272
R3485 VGND VGND.n1326 7.82272
R3486 VGND.n1327 VGND 7.82272
R3487 VGND VGND.n1330 7.82272
R3488 VGND.n1331 VGND 7.82272
R3489 VGND.n1335 VGND 7.82272
R3490 VGND VGND.n1338 7.82272
R3491 VGND.n1339 VGND 7.82272
R3492 VGND VGND.n1342 7.82272
R3493 VGND VGND.n1346 7.82272
R3494 VGND.n1347 VGND 7.82272
R3495 VGND VGND.n1350 7.82272
R3496 VGND.n1351 VGND 7.82272
R3497 VGND.n1355 VGND 7.82272
R3498 VGND VGND.n1358 7.82272
R3499 VGND.n1359 VGND 7.82272
R3500 VGND.n1363 VGND 7.82272
R3501 VGND VGND.n1366 7.82272
R3502 VGND.n1367 VGND 7.82272
R3503 VGND.n1371 VGND 7.82272
R3504 VGND.n1375 VGND 7.82272
R3505 VGND.n1379 VGND 7.82272
R3506 VGND.n1383 VGND 7.82272
R3507 VGND.n1387 VGND 7.82272
R3508 VGND.n1614 VGND 7.82272
R3509 VGND.n1613 VGND 7.82272
R3510 VGND.n1608 VGND 7.82272
R3511 VGND.n1607 VGND 7.82272
R3512 VGND.n1603 VGND 7.82272
R3513 VGND.n1599 VGND 7.82272
R3514 VGND.n1596 VGND 7.82272
R3515 VGND.n1592 VGND 7.82272
R3516 VGND.n1591 VGND 7.82272
R3517 VGND.n1587 VGND 7.82272
R3518 VGND.n1583 VGND 7.82272
R3519 VGND VGND.n1445 7.82272
R3520 VGND.n1896 VGND 7.82272
R3521 VGND.n1895 VGND 7.82272
R3522 VGND.n1890 VGND 7.82272
R3523 VGND.n1886 VGND 7.82272
R3524 VGND.n1883 VGND 7.82272
R3525 VGND VGND.n1450 7.82272
R3526 VGND.n1876 VGND 7.82272
R3527 VGND VGND.n1452 7.82272
R3528 VGND.n1869 VGND 7.82272
R3529 VGND.n1868 VGND 7.82272
R3530 VGND.n1867 VGND 7.82272
R3531 VGND.n1862 VGND 7.82272
R3532 VGND.n1859 VGND 7.82272
R3533 VGND.n1858 VGND 7.82272
R3534 VGND.n1855 VGND 7.82272
R3535 VGND VGND.n1457 7.82272
R3536 VGND.n1849 VGND 7.82272
R3537 VGND.n1848 VGND 7.82272
R3538 VGND.n1847 VGND 7.82272
R3539 VGND.n1842 VGND 7.82272
R3540 VGND.n1839 VGND 7.82272
R3541 VGND.n1838 VGND 7.82272
R3542 VGND.n1835 VGND 7.82272
R3543 VGND VGND.n1462 7.82272
R3544 VGND.n1829 VGND 7.82272
R3545 VGND.n1828 VGND 7.82272
R3546 VGND.n1827 VGND 7.82272
R3547 VGND.n1822 VGND 7.82272
R3548 VGND.n1819 VGND 7.82272
R3549 VGND.n1818 VGND 7.82272
R3550 VGND.n1814 VGND 7.82272
R3551 VGND.n1811 VGND 7.82272
R3552 VGND.n1810 VGND 7.82272
R3553 VGND.n1806 VGND 7.82272
R3554 VGND.n1802 VGND 7.82272
R3555 VGND.n1798 VGND 7.82272
R3556 VGND.n1794 VGND 7.82272
R3557 VGND.n1790 VGND 7.82272
R3558 VGND VGND.n1978 7.82272
R3559 VGND.n1979 VGND 7.82272
R3560 VGND VGND.n886 7.82272
R3561 VGND.n918 VGND 7.82272
R3562 VGND VGND.n921 7.82272
R3563 VGND VGND.n925 7.82272
R3564 VGND.n926 VGND 7.82272
R3565 VGND VGND.n929 7.82272
R3566 VGND.n930 VGND 7.82272
R3567 VGND VGND.n933 7.82272
R3568 VGND.n934 VGND 7.82272
R3569 VGND VGND.n937 7.82272
R3570 VGND.n938 VGND 7.82272
R3571 VGND VGND.n941 7.82272
R3572 VGND.n942 VGND 7.82272
R3573 VGND VGND.n945 7.82272
R3574 VGND.n946 VGND 7.82272
R3575 VGND VGND.n949 7.82272
R3576 VGND.n950 VGND 7.82272
R3577 VGND VGND.n953 7.82272
R3578 VGND.n954 VGND 7.82272
R3579 VGND VGND.n957 7.82272
R3580 VGND.n958 VGND 7.82272
R3581 VGND VGND.n961 7.82272
R3582 VGND.n962 VGND 7.82272
R3583 VGND VGND.n965 7.82272
R3584 VGND.n966 VGND 7.82272
R3585 VGND VGND.n969 7.82272
R3586 VGND.n970 VGND 7.82272
R3587 VGND VGND.n973 7.82272
R3588 VGND.n974 VGND 7.82272
R3589 VGND VGND.n977 7.82272
R3590 VGND.n978 VGND 7.82272
R3591 VGND VGND.n981 7.82272
R3592 VGND.n982 VGND 7.82272
R3593 VGND VGND.n985 7.82272
R3594 VGND.n986 VGND 7.82272
R3595 VGND VGND.n989 7.82272
R3596 VGND.n990 VGND 7.82272
R3597 VGND VGND.n993 7.82272
R3598 VGND.n994 VGND 7.82272
R3599 VGND VGND.n997 7.82272
R3600 VGND.n998 VGND 7.82272
R3601 VGND.n1002 VGND 7.82272
R3602 VGND VGND.n1005 7.82272
R3603 VGND.n1006 VGND 7.82272
R3604 VGND VGND.n1009 7.82272
R3605 VGND.n1010 VGND 7.82272
R3606 VGND VGND.n1013 7.82272
R3607 VGND VGND.n1014 7.82272
R3608 VGND VGND.n1098 7.82272
R3609 VGND.n1966 VGND 7.82272
R3610 VGND.n1965 VGND 7.82272
R3611 VGND.n1964 VGND 7.82272
R3612 VGND.n1962 VGND 7.82272
R3613 VGND.n1959 VGND 7.82272
R3614 VGND.n1958 VGND 7.82272
R3615 VGND.n1954 VGND 7.82272
R3616 VGND.n1950 VGND 7.82272
R3617 VGND.n1947 VGND 7.82272
R3618 VGND.n1943 VGND 7.82272
R3619 VGND.n1942 VGND 7.82272
R3620 VGND.n1938 VGND 7.82272
R3621 VGND.n1934 VGND 7.82272
R3622 VGND.n2369 VGND 7.82272
R3623 VGND.n2366 VGND 7.82272
R3624 VGND.n2362 VGND 7.82272
R3625 VGND.n2361 VGND 7.82272
R3626 VGND.n2357 VGND 7.82272
R3627 VGND.n2353 VGND 7.82272
R3628 VGND.n2350 VGND 7.82272
R3629 VGND.n2346 VGND 7.82272
R3630 VGND.n2345 VGND 7.82272
R3631 VGND.n2341 VGND 7.82272
R3632 VGND.n2337 VGND 7.82272
R3633 VGND.n2329 VGND 7.82272
R3634 VGND VGND.n774 7.82272
R3635 VGND.n2322 VGND 7.82272
R3636 VGND.n2321 VGND 7.82272
R3637 VGND.n2315 VGND 7.82272
R3638 VGND.n2313 VGND 7.82272
R3639 VGND VGND.n782 7.82272
R3640 VGND.n2306 VGND 7.82272
R3641 VGND.n2305 VGND 7.82272
R3642 VGND.n2299 VGND 7.82272
R3643 VGND.n2297 VGND 7.82272
R3644 VGND.n2193 VGND 7.82272
R3645 VGND.n2189 VGND 7.82272
R3646 VGND.n2188 VGND 7.82272
R3647 VGND.n2184 VGND 7.82272
R3648 VGND.n2180 VGND 7.82272
R3649 VGND.n2177 VGND 7.82272
R3650 VGND.n2173 VGND 7.82272
R3651 VGND.n2169 VGND 7.82272
R3652 VGND.n2165 VGND 7.82272
R3653 VGND.n2164 VGND 7.82272
R3654 VGND.n2161 VGND 7.82272
R3655 VGND.n2160 VGND 7.82272
R3656 VGND.n2156 VGND 7.82272
R3657 VGND.n2153 VGND 7.82272
R3658 VGND.n2152 VGND 7.82272
R3659 VGND.n2149 VGND 7.82272
R3660 VGND.n2145 VGND 7.82272
R3661 VGND.n2144 VGND 7.82272
R3662 VGND.n2141 VGND 7.82272
R3663 VGND.n2140 VGND 7.82272
R3664 VGND.n2136 VGND 7.82272
R3665 VGND.n2133 VGND 7.82272
R3666 VGND.n2132 VGND 7.82272
R3667 VGND.n2129 VGND 7.82272
R3668 VGND.n2125 VGND 7.82272
R3669 VGND.n2124 VGND 7.82272
R3670 VGND.n2121 VGND 7.82272
R3671 VGND.n2120 VGND 7.82272
R3672 VGND.n2116 VGND 7.82272
R3673 VGND.n2113 VGND 7.82272
R3674 VGND.n2112 VGND 7.82272
R3675 VGND.n2108 VGND 7.82272
R3676 VGND.n2105 VGND 7.82272
R3677 VGND.n2104 VGND 7.82272
R3678 VGND.n2100 VGND 7.82272
R3679 VGND.n2096 VGND 7.82272
R3680 VGND.n2092 VGND 7.82272
R3681 VGND.n2088 VGND 7.82272
R3682 VGND.n2084 VGND 7.82272
R3683 VGND.n2721 VGND 7.82272
R3684 VGND.n2715 VGND 7.82272
R3685 VGND.n2714 VGND 7.82272
R3686 VGND VGND.n88 7.82272
R3687 VGND.n2706 VGND 7.82272
R3688 VGND.n2705 VGND 7.82272
R3689 VGND.n2699 VGND 7.82272
R3690 VGND.n2697 VGND 7.82272
R3691 VGND.n2691 VGND 7.82272
R3692 VGND.n2690 VGND 7.82272
R3693 VGND.n2689 VGND 7.82272
R3694 VGND VGND.n104 7.82272
R3695 VGND.n2682 VGND 7.82272
R3696 VGND.n2681 VGND 7.82272
R3697 VGND VGND.n107 7.82272
R3698 VGND.n2675 VGND 7.82272
R3699 VGND.n2673 VGND 7.82272
R3700 VGND VGND.n111 7.82272
R3701 VGND.n2667 VGND 7.82272
R3702 VGND.n2666 VGND 7.82272
R3703 VGND VGND.n112 7.82272
R3704 VGND.n2659 VGND 7.82272
R3705 VGND.n2658 VGND 7.82272
R3706 VGND.n2657 VGND 7.82272
R3707 VGND.n2651 VGND 7.82272
R3708 VGND.n2650 VGND 7.82272
R3709 VGND.n2649 VGND 7.82272
R3710 VGND VGND.n124 7.82272
R3711 VGND.n2642 VGND 7.82272
R3712 VGND.n2641 VGND 7.82272
R3713 VGND VGND.n128 7.82272
R3714 VGND.n2634 VGND 7.82272
R3715 VGND.n2633 VGND 7.82272
R3716 VGND VGND.n132 7.82272
R3717 VGND.n2626 VGND 7.82272
R3718 VGND VGND.n133 7.82272
R3719 VGND.n2618 VGND 7.82272
R3720 VGND VGND.n137 7.82272
R3721 VGND.n2610 VGND 7.82272
R3722 VGND VGND.n601 7.82272
R3723 VGND.n617 VGND 7.82272
R3724 VGND.n621 VGND 7.82272
R3725 VGND VGND.n624 7.82272
R3726 VGND VGND.n628 7.82272
R3727 VGND.n629 VGND 7.82272
R3728 VGND VGND.n632 7.82272
R3729 VGND VGND.n636 7.82272
R3730 VGND VGND.n543 7.82272
R3731 VGND VGND.n553 7.82272
R3732 VGND VGND.n557 7.82272
R3733 VGND VGND.n561 7.82272
R3734 VGND VGND.n565 7.82272
R3735 VGND VGND.n569 7.82272
R3736 VGND.n571 VGND 7.82272
R3737 VGND.n1073 VGND 7.82272
R3738 VGND VGND.n1079 7.82272
R3739 VGND.n1081 VGND 7.82272
R3740 VGND.n1047 VGND 7.52991
R3741 VGND VGND.n1068 7.52991
R3742 VGND.n1061 VGND 7.52991
R3743 VGND.n1056 VGND 7.52991
R3744 VGND.n1051 VGND 7.52991
R3745 VGND.n1928 VGND 7.43276
R3746 VGND.n1783 VGND 7.43276
R3747 VGND.n1655 VGND.n1121 7.23528
R3748 VGND.n1694 VGND.n1656 7.23528
R3749 VGND.n1693 VGND.n1692 7.23528
R3750 VGND.n2385 VGND.n735 7.23528
R3751 VGND.n2384 VGND.n736 7.23528
R3752 VGND.n2284 VGND.n807 7.23528
R3753 VGND.n471 VGND.n405 6.93569
R3754 VGND.n1049 VGND.n1048 6.77697
R3755 VGND.n647 VGND.n599 6.77697
R3756 VGND.n644 VGND.n643 6.77697
R3757 VGND.n605 VGND.n604 6.77697
R3758 VGND.n608 VGND.n607 6.77697
R3759 VGND.n586 VGND.n585 6.77697
R3760 VGND.n2241 VGND.n2236 6.77697
R3761 VGND.n2238 VGND.n2237 6.77697
R3762 VGND.n2200 VGND.n2075 6.77697
R3763 VGND.n832 VGND.n826 6.77697
R3764 VGND.n828 VGND.n827 6.77697
R3765 VGND.n1399 VGND.n1194 6.77697
R3766 VGND.n1396 VGND.n1395 6.77697
R3767 VGND.n1199 VGND.n1198 6.77697
R3768 VGND.n729 VGND.n728 6.77697
R3769 VGND.n2391 VGND.n712 6.77697
R3770 VGND.n1196 VGND.n1195 6.77697
R3771 VGND.n1541 VGND.n1540 6.77697
R3772 VGND.n1711 VGND.n1705 6.77697
R3773 VGND.n1707 VGND.n1706 6.77697
R3774 VGND.n1637 VGND.n1636 6.77697
R3775 VGND.n1641 VGND.n1620 6.77697
R3776 VGND.n1775 VGND.n1774 6.77697
R3777 VGND.n2036 VGND.n881 6.77697
R3778 VGND.n2033 VGND.n2032 6.77697
R3779 VGND.n1027 VGND.n1026 6.77697
R3780 VGND.n1024 VGND.n1023 6.77697
R3781 VGND.n1101 VGND.n1100 6.77697
R3782 VGND.n1118 VGND.n1117 6.77697
R3783 VGND.n2077 VGND.n2076 6.77697
R3784 VGND.n588 VGND.n587 6.77697
R3785 VGND.n1046 VGND.n1045 6.77697
R3786 VGND.n1063 VGND.n1062 6.77697
R3787 VGND.n1058 VGND.n1057 6.77697
R3788 VGND.n1053 VGND.n1052 6.77697
R3789 VGND.n405 VGND 6.4005
R3790 VGND VGND.n527 6.4005
R3791 VGND.n300 VGND.n202 6.36865
R3792 VGND.n303 VGND.n200 6.1255
R3793 VGND.n304 VGND.n199 6.1255
R3794 VGND.n305 VGND.n198 6.1255
R3795 VGND.n306 VGND.n197 6.1255
R3796 VGND.n307 VGND.n196 6.1255
R3797 VGND.n308 VGND.n195 6.1255
R3798 VGND.n309 VGND.n194 6.1255
R3799 VGND.n310 VGND.n193 6.1255
R3800 VGND.n311 VGND.n192 6.1255
R3801 VGND.n312 VGND.n191 6.1255
R3802 VGND.n313 VGND.n190 6.1255
R3803 VGND.n314 VGND.n189 6.1255
R3804 VGND.n315 VGND.n188 6.1255
R3805 VGND.n316 VGND.n187 6.1255
R3806 VGND.n317 VGND.n186 6.1255
R3807 VGND.n318 VGND.n185 6.1255
R3808 VGND.n319 VGND.n184 6.1255
R3809 VGND.n320 VGND.n183 6.1255
R3810 VGND.n321 VGND.n182 6.1255
R3811 VGND.n322 VGND.n181 6.1255
R3812 VGND.n323 VGND.n180 6.1255
R3813 VGND.n324 VGND.n179 6.1255
R3814 VGND.n325 VGND.n178 6.1255
R3815 VGND.n326 VGND.n177 6.1255
R3816 VGND.n327 VGND.n176 6.1255
R3817 VGND.n328 VGND.n175 6.1255
R3818 VGND.n329 VGND.n174 6.1255
R3819 VGND.n330 VGND.n173 6.1255
R3820 VGND.n331 VGND.n172 6.1255
R3821 VGND.n332 VGND.n171 6.1255
R3822 VGND.n299 VGND.n201 6.1255
R3823 VGND.n298 VGND.n200 6.1255
R3824 VGND.n297 VGND.n199 6.1255
R3825 VGND.n296 VGND.n198 6.1255
R3826 VGND.n295 VGND.n197 6.1255
R3827 VGND.n294 VGND.n196 6.1255
R3828 VGND.n293 VGND.n195 6.1255
R3829 VGND.n292 VGND.n194 6.1255
R3830 VGND.n291 VGND.n193 6.1255
R3831 VGND.n290 VGND.n192 6.1255
R3832 VGND.n289 VGND.n191 6.1255
R3833 VGND.n288 VGND.n190 6.1255
R3834 VGND.n287 VGND.n189 6.1255
R3835 VGND.n286 VGND.n188 6.1255
R3836 VGND.n285 VGND.n187 6.1255
R3837 VGND.n284 VGND.n186 6.1255
R3838 VGND.n283 VGND.n185 6.1255
R3839 VGND.n282 VGND.n184 6.1255
R3840 VGND.n281 VGND.n183 6.1255
R3841 VGND.n280 VGND.n182 6.1255
R3842 VGND.n279 VGND.n181 6.1255
R3843 VGND.n278 VGND.n180 6.1255
R3844 VGND.n277 VGND.n179 6.1255
R3845 VGND.n276 VGND.n178 6.1255
R3846 VGND.n275 VGND.n177 6.1255
R3847 VGND.n274 VGND.n176 6.1255
R3848 VGND.n273 VGND.n175 6.1255
R3849 VGND.n272 VGND.n174 6.1255
R3850 VGND.n271 VGND.n173 6.1255
R3851 VGND.n270 VGND.n172 6.1255
R3852 VGND.n269 VGND.n171 6.1255
R3853 VGND.n299 VGND.n203 6.1255
R3854 VGND.n298 VGND.n204 6.1255
R3855 VGND.n297 VGND.n205 6.1255
R3856 VGND.n296 VGND.n206 6.1255
R3857 VGND.n295 VGND.n207 6.1255
R3858 VGND.n294 VGND.n208 6.1255
R3859 VGND.n293 VGND.n209 6.1255
R3860 VGND.n292 VGND.n210 6.1255
R3861 VGND.n291 VGND.n211 6.1255
R3862 VGND.n290 VGND.n212 6.1255
R3863 VGND.n289 VGND.n213 6.1255
R3864 VGND.n288 VGND.n214 6.1255
R3865 VGND.n287 VGND.n215 6.1255
R3866 VGND.n286 VGND.n216 6.1255
R3867 VGND.n285 VGND.n217 6.1255
R3868 VGND.n284 VGND.n218 6.1255
R3869 VGND.n283 VGND.n219 6.1255
R3870 VGND.n282 VGND.n220 6.1255
R3871 VGND.n281 VGND.n221 6.1255
R3872 VGND.n280 VGND.n222 6.1255
R3873 VGND.n279 VGND.n223 6.1255
R3874 VGND.n278 VGND.n224 6.1255
R3875 VGND.n277 VGND.n225 6.1255
R3876 VGND.n276 VGND.n226 6.1255
R3877 VGND.n275 VGND.n227 6.1255
R3878 VGND.n274 VGND.n228 6.1255
R3879 VGND.n273 VGND.n229 6.1255
R3880 VGND.n272 VGND.n230 6.1255
R3881 VGND.n271 VGND.n231 6.1255
R3882 VGND.n270 VGND.n232 6.1255
R3883 VGND.n269 VGND.n233 6.1255
R3884 VGND.n263 VGND.n233 6.1255
R3885 VGND.n262 VGND.n232 6.1255
R3886 VGND.n261 VGND.n231 6.1255
R3887 VGND.n260 VGND.n230 6.1255
R3888 VGND.n259 VGND.n229 6.1255
R3889 VGND.n258 VGND.n228 6.1255
R3890 VGND.n257 VGND.n227 6.1255
R3891 VGND.n256 VGND.n226 6.1255
R3892 VGND.n255 VGND.n225 6.1255
R3893 VGND.n254 VGND.n224 6.1255
R3894 VGND.n253 VGND.n223 6.1255
R3895 VGND.n252 VGND.n222 6.1255
R3896 VGND.n251 VGND.n221 6.1255
R3897 VGND.n250 VGND.n220 6.1255
R3898 VGND.n249 VGND.n219 6.1255
R3899 VGND.n248 VGND.n218 6.1255
R3900 VGND.n247 VGND.n217 6.1255
R3901 VGND.n246 VGND.n216 6.1255
R3902 VGND.n245 VGND.n215 6.1255
R3903 VGND.n244 VGND.n214 6.1255
R3904 VGND.n243 VGND.n213 6.1255
R3905 VGND.n242 VGND.n212 6.1255
R3906 VGND.n241 VGND.n211 6.1255
R3907 VGND.n240 VGND.n210 6.1255
R3908 VGND.n239 VGND.n209 6.1255
R3909 VGND.n238 VGND.n208 6.1255
R3910 VGND.n237 VGND.n207 6.1255
R3911 VGND.n236 VGND.n206 6.1255
R3912 VGND.n235 VGND.n205 6.1255
R3913 VGND.n234 VGND.n204 6.1255
R3914 VGND.n267 VGND.n266 6.1255
R3915 VGND.n268 VGND.n267 6.1255
R3916 VGND.n268 VGND.n170 6.1255
R3917 VGND.n333 VGND.n170 6.1255
R3918 VGND.n476 VGND.n401 6.1255
R3919 VGND.n477 VGND.n399 6.1255
R3920 VGND.n478 VGND.n397 6.1255
R3921 VGND.n479 VGND.n395 6.1255
R3922 VGND.n480 VGND.n393 6.1255
R3923 VGND.n481 VGND.n391 6.1255
R3924 VGND.n482 VGND.n389 6.1255
R3925 VGND.n483 VGND.n387 6.1255
R3926 VGND.n484 VGND.n385 6.1255
R3927 VGND.n485 VGND.n383 6.1255
R3928 VGND.n486 VGND.n381 6.1255
R3929 VGND.n487 VGND.n379 6.1255
R3930 VGND.n488 VGND.n377 6.1255
R3931 VGND.n489 VGND.n375 6.1255
R3932 VGND.n490 VGND.n373 6.1255
R3933 VGND.n491 VGND.n371 6.1255
R3934 VGND.n492 VGND.n369 6.1255
R3935 VGND.n493 VGND.n367 6.1255
R3936 VGND.n494 VGND.n365 6.1255
R3937 VGND.n495 VGND.n363 6.1255
R3938 VGND.n496 VGND.n361 6.1255
R3939 VGND.n497 VGND.n359 6.1255
R3940 VGND.n498 VGND.n357 6.1255
R3941 VGND.n499 VGND.n355 6.1255
R3942 VGND.n500 VGND.n353 6.1255
R3943 VGND.n501 VGND.n351 6.1255
R3944 VGND.n502 VGND.n349 6.1255
R3945 VGND.n503 VGND.n347 6.1255
R3946 VGND.n504 VGND.n345 6.1255
R3947 VGND.n505 VGND.n343 6.1255
R3948 VGND.n506 VGND.n342 6.1255
R3949 VGND.n506 VGND.n337 6.1255
R3950 VGND.n505 VGND.n344 6.1255
R3951 VGND.n504 VGND.n346 6.1255
R3952 VGND.n503 VGND.n348 6.1255
R3953 VGND.n502 VGND.n350 6.1255
R3954 VGND.n501 VGND.n352 6.1255
R3955 VGND.n500 VGND.n354 6.1255
R3956 VGND.n499 VGND.n356 6.1255
R3957 VGND.n498 VGND.n358 6.1255
R3958 VGND.n497 VGND.n360 6.1255
R3959 VGND.n496 VGND.n362 6.1255
R3960 VGND.n495 VGND.n364 6.1255
R3961 VGND.n494 VGND.n366 6.1255
R3962 VGND.n493 VGND.n368 6.1255
R3963 VGND.n492 VGND.n370 6.1255
R3964 VGND.n491 VGND.n372 6.1255
R3965 VGND.n490 VGND.n374 6.1255
R3966 VGND.n489 VGND.n376 6.1255
R3967 VGND.n488 VGND.n378 6.1255
R3968 VGND.n487 VGND.n380 6.1255
R3969 VGND.n486 VGND.n382 6.1255
R3970 VGND.n485 VGND.n384 6.1255
R3971 VGND.n484 VGND.n386 6.1255
R3972 VGND.n483 VGND.n388 6.1255
R3973 VGND.n482 VGND.n390 6.1255
R3974 VGND.n481 VGND.n392 6.1255
R3975 VGND.n480 VGND.n394 6.1255
R3976 VGND.n479 VGND.n396 6.1255
R3977 VGND.n478 VGND.n398 6.1255
R3978 VGND.n477 VGND.n400 6.1255
R3979 VGND.n476 VGND.n402 6.1255
R3980 VGND.n436 VGND.n337 6.1255
R3981 VGND.n435 VGND.n344 6.1255
R3982 VGND.n434 VGND.n346 6.1255
R3983 VGND.n433 VGND.n348 6.1255
R3984 VGND.n432 VGND.n350 6.1255
R3985 VGND.n431 VGND.n352 6.1255
R3986 VGND.n430 VGND.n354 6.1255
R3987 VGND.n429 VGND.n356 6.1255
R3988 VGND.n428 VGND.n358 6.1255
R3989 VGND.n427 VGND.n360 6.1255
R3990 VGND.n426 VGND.n362 6.1255
R3991 VGND.n425 VGND.n364 6.1255
R3992 VGND.n424 VGND.n366 6.1255
R3993 VGND.n423 VGND.n368 6.1255
R3994 VGND.n422 VGND.n370 6.1255
R3995 VGND.n421 VGND.n372 6.1255
R3996 VGND.n420 VGND.n374 6.1255
R3997 VGND.n419 VGND.n376 6.1255
R3998 VGND.n418 VGND.n378 6.1255
R3999 VGND.n417 VGND.n380 6.1255
R4000 VGND.n416 VGND.n382 6.1255
R4001 VGND.n415 VGND.n384 6.1255
R4002 VGND.n414 VGND.n386 6.1255
R4003 VGND.n413 VGND.n388 6.1255
R4004 VGND.n412 VGND.n390 6.1255
R4005 VGND.n411 VGND.n392 6.1255
R4006 VGND.n410 VGND.n394 6.1255
R4007 VGND.n409 VGND.n396 6.1255
R4008 VGND.n408 VGND.n398 6.1255
R4009 VGND.n407 VGND.n400 6.1255
R4010 VGND.n406 VGND.n402 6.1255
R4011 VGND.n437 VGND.n436 6.1255
R4012 VGND.n438 VGND.n435 6.1255
R4013 VGND.n439 VGND.n434 6.1255
R4014 VGND.n440 VGND.n433 6.1255
R4015 VGND.n441 VGND.n432 6.1255
R4016 VGND.n442 VGND.n431 6.1255
R4017 VGND.n443 VGND.n430 6.1255
R4018 VGND.n444 VGND.n429 6.1255
R4019 VGND.n445 VGND.n428 6.1255
R4020 VGND.n446 VGND.n427 6.1255
R4021 VGND.n447 VGND.n426 6.1255
R4022 VGND.n448 VGND.n425 6.1255
R4023 VGND.n449 VGND.n424 6.1255
R4024 VGND.n450 VGND.n423 6.1255
R4025 VGND.n451 VGND.n422 6.1255
R4026 VGND.n452 VGND.n421 6.1255
R4027 VGND.n453 VGND.n420 6.1255
R4028 VGND.n454 VGND.n419 6.1255
R4029 VGND.n455 VGND.n418 6.1255
R4030 VGND.n456 VGND.n417 6.1255
R4031 VGND.n457 VGND.n416 6.1255
R4032 VGND.n458 VGND.n415 6.1255
R4033 VGND.n459 VGND.n414 6.1255
R4034 VGND.n460 VGND.n413 6.1255
R4035 VGND.n461 VGND.n412 6.1255
R4036 VGND.n462 VGND.n411 6.1255
R4037 VGND.n463 VGND.n410 6.1255
R4038 VGND.n464 VGND.n409 6.1255
R4039 VGND.n465 VGND.n408 6.1255
R4040 VGND.n466 VGND.n407 6.1255
R4041 VGND.n467 VGND.n406 6.1255
R4042 VGND.n468 VGND.n404 6.1255
R4043 VGND.n470 VGND.n469 6.1255
R4044 VGND.n475 VGND.n474 6.1255
R4045 VGND.n474 VGND.n404 6.1255
R4046 VGND.n473 VGND.n472 6.1255
R4047 VGND.n2521 VGND.n163 6.05932
R4048 VGND.n2520 VGND.n2519 6.05932
R4049 VGND.n2514 VGND.n167 6.05932
R4050 VGND.n509 VGND.n339 6.05932
R4051 VGND.n521 VGND.n340 6.05932
R4052 VGND.n517 VGND.n516 6.05932
R4053 VGND.n1916 VGND 5.8572
R4054 VGND.n2767 VGND 5.81001
R4055 VGND.n301 VGND.n300 5.77624
R4056 VGND.n473 VGND.n471 5.77624
R4057 VGND.n2492 VGND.n2466 5.21532
R4058 VGND.n2502 VGND.n530 5.21532
R4059 VGND.n2398 VGND.n2396 5.21532
R4060 VGND.n1393 VGND.n1392 5.21532
R4061 VGND.n1646 VGND.n1567 5.21532
R4062 VGND.n1987 VGND.n885 5.21532
R4063 VGND.n2030 VGND.n882 5.21532
R4064 VGND.n2374 VGND.n757 5.21532
R4065 VGND.n2291 VGND.n2290 5.21532
R4066 VGND.n2729 VGND.n48 5.21532
R4067 VGND.n2603 VGND.n141 5.21532
R4068 VGND.n613 VGND.n612 5.21532
R4069 VGND.n641 VGND.n640 5.21532
R4070 VGND.n526 VGND.n334 5.20068
R4071 VGND.n525 VGND.n335 5.20068
R4072 VGND.n524 VGND.n523 5.20068
R4073 VGND.n507 VGND.n159 5.20068
R4074 VGND.n2382 VGND.n736 4.6505
R4075 VGND.n735 VGND.n734 4.6505
R4076 VGND.n1693 VGND.n1657 4.6505
R4077 VGND.n1696 VGND.n1656 4.6505
R4078 VGND.n1548 VGND.n1121 4.6505
R4079 VGND.n2384 VGND.n2383 4.6505
R4080 VGND.n2386 VGND.n2385 4.6505
R4081 VGND.n1692 VGND.n1691 4.6505
R4082 VGND.n1695 VGND.n1694 4.6505
R4083 VGND.n1655 VGND.n1654 4.6505
R4084 VGND.n2284 VGND.n2283 4.6505
R4085 VGND.n808 VGND.n807 4.6505
R4086 VGND.n155 VGND.n147 4.63736
R4087 VGND.n2528 VGND.n2526 4.6334
R4088 VGND.n2526 VGND.n158 4.6334
R4089 VGND.n2526 VGND.n153 4.6334
R4090 VGND.n2526 VGND.n152 4.6334
R4091 VGND.n2526 VGND.n151 4.6334
R4092 VGND.n2526 VGND.n150 4.6334
R4093 VGND.n2526 VGND.n149 4.6334
R4094 VGND.n2526 VGND.n148 4.6334
R4095 VGND.n1783 VGND 4.62272
R4096 VGND.n1928 VGND 4.62272
R4097 VGND.n265 VGND.n264 4.59498
R4098 VGND.n2513 VGND.n2511 4.59498
R4099 VGND.n510 VGND.n341 4.59498
R4100 VGND.n514 VGND.n512 4.59498
R4101 VGND.n163 VGND.n161 4.5005
R4102 VGND.n2520 VGND.n162 4.5005
R4103 VGND.n2522 VGND.n2521 4.5005
R4104 VGND.n2517 VGND.n167 4.5005
R4105 VGND.n2519 VGND.n2518 4.5005
R4106 VGND.n2515 VGND.n2514 4.5005
R4107 VGND.n339 VGND.n338 4.5005
R4108 VGND.n522 VGND.n521 4.5005
R4109 VGND.n340 VGND.n336 4.5005
R4110 VGND.n517 VGND.n513 4.5005
R4111 VGND.n516 VGND.n515 4.5005
R4112 VGND.n509 VGND.n508 4.5005
R4113 VGND.n1066 VGND.n1050 3.95786
R4114 VGND.n264 VGND.n164 3.9554
R4115 VGND.n2513 VGND.n2512 3.9554
R4116 VGND.n511 VGND.n510 3.9554
R4117 VGND.n518 VGND.n512 3.9554
R4118 VGND.n659 VGND.n589 3.95489
R4119 VGND.n1055 VGND.n1054 3.9165
R4120 VGND.n1060 VGND.n1059 3.9165
R4121 VGND.n1065 VGND.n1064 3.9165
R4122 VGND.n1067 VGND.n1066 3.9165
R4123 VGND.n651 VGND.n598 3.90993
R4124 VGND.n657 VGND.n591 3.90993
R4125 VGND.n660 VGND.n659 3.90993
R4126 VGND.n2245 VGND.n2235 3.90993
R4127 VGND.n2273 VGND.n2202 3.90993
R4128 VGND.n1403 VGND.n1193 3.90993
R4129 VGND.n1431 VGND.n1160 3.90993
R4130 VGND.n2392 VGND.n2390 3.90993
R4131 VGND.n2389 VGND.n730 3.90993
R4132 VGND.n1402 VGND.n1401 3.90993
R4133 VGND.n1432 VGND.n1159 3.90993
R4134 VGND.n1779 VGND.n1778 3.90993
R4135 VGND.n1708 VGND.n1704 3.90993
R4136 VGND.n1642 VGND.n1640 3.90993
R4137 VGND.n1639 VGND.n1638 3.90993
R4138 VGND.n1714 VGND.n1713 3.90993
R4139 VGND.n1777 VGND.n1776 3.90993
R4140 VGND.n2040 VGND.n880 3.90993
R4141 VGND.n2068 VGND.n847 3.90993
R4142 VGND.n2039 VGND.n2038 3.90993
R4143 VGND.n2069 VGND.n846 3.90993
R4144 VGND.n1924 VGND.n1923 3.90993
R4145 VGND.n1120 VGND.n1119 3.90993
R4146 VGND.n829 VGND.n825 3.90993
R4147 VGND.n835 VGND.n834 3.90993
R4148 VGND.n2244 VGND.n2243 3.90993
R4149 VGND.n2274 VGND.n2074 3.90993
R4150 VGND.n656 VGND.n592 3.90993
R4151 VGND.n650 VGND.n649 3.90993
R4152 VGND.n2727 VGND.n81 3.81746
R4153 VGND.n303 VGND.n302 3.54879
R4154 VGND.n234 VGND.n202 3.54879
R4155 VGND.n403 VGND.n401 3.54879
R4156 VGND.n2507 VGND 3.43893
R4157 VGND.n2508 VGND 3.43867
R4158 VGND.n2512 VGND.n167 3.4105
R4159 VGND.n2519 VGND.n166 3.4105
R4160 VGND.n2520 VGND.n165 3.4105
R4161 VGND.n2521 VGND.n164 3.4105
R4162 VGND.n518 VGND.n517 3.4105
R4163 VGND.n519 VGND.n340 3.4105
R4164 VGND.n521 VGND.n520 3.4105
R4165 VGND.n511 VGND.n339 3.4105
R4166 VGND.n1687 VGND.n1682 3.4105
R4167 VGND.n1687 VGND.n1686 3.4105
R4168 VGND.n1689 VGND.n1680 3.4105
R4169 VGND.n1690 VGND.n1689 3.4105
R4170 VGND.n2388 VGND.n731 3.4105
R4171 VGND.n2388 VGND.n2387 3.4105
R4172 VGND.n1437 VGND.n1158 3.4105
R4173 VGND.n1437 VGND.n1436 3.4105
R4174 VGND.n1913 VGND.n1441 3.4105
R4175 VGND.n1913 VGND.n1912 3.4105
R4176 VGND.n1652 VGND.n1651 3.4105
R4177 VGND.n1653 VGND.n1652 3.4105
R4178 VGND.n1697 VGND.n1546 3.4105
R4179 VGND.n1547 VGND.n1546 3.4105
R4180 VGND.n1701 VGND.n1700 3.4105
R4181 VGND.n1700 VGND.n1544 3.4105
R4182 VGND.n844 VGND.n840 3.4105
R4183 VGND.n842 VGND.n840 3.4105
R4184 VGND.n1156 VGND.n1151 3.4105
R4185 VGND.n1156 VGND.n1155 3.4105
R4186 VGND.n1920 VGND.n1919 3.4105
R4187 VGND.n1919 VGND.n1122 3.4105
R4188 VGND.n154 VGND.n10 3.4105
R4189 VGND.n156 VGND.n10 3.4105
R4190 VGND.n2379 VGND.n737 3.4105
R4191 VGND.n738 VGND.n737 3.4105
R4192 VGND.n2281 VGND.n836 3.4105
R4193 VGND.n2282 VGND.n2281 3.4105
R4194 VGND.n2279 VGND.n838 3.4105
R4195 VGND.n2279 VGND.n2278 3.4105
R4196 VGND.n2531 VGND.n144 3.4105
R4197 VGND.n2531 VGND.n2530 3.4105
R4198 VGND VGND.n2285 3.38273
R4199 VGND VGND.n1922 3.38248
R4200 VGND.n266 VGND.n265 3.37918
R4201 VGND.n342 VGND.n341 3.37918
R4202 VGND.n1786 VGND.n1783 3.2005
R4203 VGND.n1930 VGND.n1928 3.2005
R4204 VGND.n2523 VGND.n2522 3.13653
R4205 VGND.n2518 VGND.n168 3.13653
R4206 VGND.n2516 VGND.n2515 3.13653
R4207 VGND.n523 VGND.n336 3.13653
R4208 VGND.n515 VGND.n335 3.13653
R4209 VGND.n507 VGND.n338 3.13653
R4210 VGND.n2516 VGND.n169 2.91731
R4211 VGND.n168 VGND.n160 2.91731
R4212 VGND.n2524 VGND.n2523 2.91731
R4213 VGND.n2510 VGND.n2509 2.91731
R4214 VGND.n2523 VGND.n161 2.79829
R4215 VGND.n168 VGND.n162 2.79829
R4216 VGND.n2517 VGND.n2516 2.79829
R4217 VGND.n2511 VGND.n2510 2.79829
R4218 VGND.n513 VGND.n335 2.79829
R4219 VGND.n514 VGND.n334 2.79829
R4220 VGND.n523 VGND.n522 2.79829
R4221 VGND.n508 VGND.n507 2.79829
R4222 VGND VGND.n2496 2.60791
R4223 VGND VGND.n2494 2.60791
R4224 VGND VGND.n2466 2.60791
R4225 VGND.n2489 VGND 2.60791
R4226 VGND.n2485 VGND 2.60791
R4227 VGND.n2481 VGND 2.60791
R4228 VGND VGND.n2480 2.60791
R4229 VGND VGND.n2476 2.60791
R4230 VGND.n2473 VGND 2.60791
R4231 VGND VGND.n2472 2.60791
R4232 VGND VGND.n2468 2.60791
R4233 VGND.n2502 VGND 2.60791
R4234 VGND VGND.n2434 2.60791
R4235 VGND VGND.n2432 2.60791
R4236 VGND VGND.n2430 2.60791
R4237 VGND VGND.n2426 2.60791
R4238 VGND.n2423 VGND 2.60791
R4239 VGND.n2419 VGND 2.60791
R4240 VGND.n2415 VGND 2.60791
R4241 VGND VGND.n2414 2.60791
R4242 VGND VGND.n2410 2.60791
R4243 VGND.n2407 VGND 2.60791
R4244 VGND.n2403 VGND 2.60791
R4245 VGND.n2399 VGND 2.60791
R4246 VGND.n2396 VGND 2.60791
R4247 VGND VGND.n1274 2.60791
R4248 VGND.n1275 VGND 2.60791
R4249 VGND.n1279 VGND 2.60791
R4250 VGND.n1283 VGND 2.60791
R4251 VGND.n1286 VGND 2.60791
R4252 VGND.n1290 VGND 2.60791
R4253 VGND.n1294 VGND 2.60791
R4254 VGND.n1295 VGND 2.60791
R4255 VGND.n1299 VGND 2.60791
R4256 VGND.n1303 VGND 2.60791
R4257 VGND.n1307 VGND 2.60791
R4258 VGND.n1310 VGND 2.60791
R4259 VGND.n1311 VGND 2.60791
R4260 VGND.n1314 VGND 2.60791
R4261 VGND.n1318 VGND 2.60791
R4262 VGND.n1319 VGND 2.60791
R4263 VGND.n1322 VGND 2.60791
R4264 VGND.n1323 VGND 2.60791
R4265 VGND.n1327 VGND 2.60791
R4266 VGND.n1330 VGND 2.60791
R4267 VGND.n1331 VGND 2.60791
R4268 VGND.n1334 VGND 2.60791
R4269 VGND.n1338 VGND 2.60791
R4270 VGND.n1339 VGND 2.60791
R4271 VGND.n1342 VGND 2.60791
R4272 VGND.n1343 VGND 2.60791
R4273 VGND.n1347 VGND 2.60791
R4274 VGND.n1350 VGND 2.60791
R4275 VGND.n1351 VGND 2.60791
R4276 VGND.n1354 VGND 2.60791
R4277 VGND.n1358 VGND 2.60791
R4278 VGND.n1359 VGND 2.60791
R4279 VGND.n1362 VGND 2.60791
R4280 VGND.n1366 VGND 2.60791
R4281 VGND.n1367 VGND 2.60791
R4282 VGND.n1370 VGND 2.60791
R4283 VGND.n1374 VGND 2.60791
R4284 VGND.n1378 VGND 2.60791
R4285 VGND.n1382 VGND 2.60791
R4286 VGND.n1386 VGND 2.60791
R4287 VGND.n1390 VGND 2.60791
R4288 VGND.n1393 VGND 2.60791
R4289 VGND VGND.n1615 2.60791
R4290 VGND VGND.n1613 2.60791
R4291 VGND VGND.n1611 2.60791
R4292 VGND VGND.n1607 2.60791
R4293 VGND.n1604 VGND 2.60791
R4294 VGND.n1600 VGND 2.60791
R4295 VGND.n1596 VGND 2.60791
R4296 VGND VGND.n1595 2.60791
R4297 VGND VGND.n1591 2.60791
R4298 VGND.n1588 VGND 2.60791
R4299 VGND.n1584 VGND 2.60791
R4300 VGND.n1580 VGND 2.60791
R4301 VGND.n1646 VGND 2.60791
R4302 VGND.n1903 VGND 2.60791
R4303 VGND VGND.n1902 2.60791
R4304 VGND.n1897 VGND 2.60791
R4305 VGND VGND.n1895 2.60791
R4306 VGND.n1891 VGND 2.60791
R4307 VGND.n1887 VGND 2.60791
R4308 VGND.n1883 VGND 2.60791
R4309 VGND VGND.n1882 2.60791
R4310 VGND.n1877 VGND 2.60791
R4311 VGND VGND.n1875 2.60791
R4312 VGND.n1869 VGND 2.60791
R4313 VGND VGND.n1868 2.60791
R4314 VGND VGND.n1867 2.60791
R4315 VGND.n1863 VGND 2.60791
R4316 VGND.n1859 VGND 2.60791
R4317 VGND VGND.n1858 2.60791
R4318 VGND.n1855 VGND 2.60791
R4319 VGND VGND.n1854 2.60791
R4320 VGND.n1849 VGND 2.60791
R4321 VGND VGND.n1848 2.60791
R4322 VGND VGND.n1847 2.60791
R4323 VGND.n1843 VGND 2.60791
R4324 VGND.n1839 VGND 2.60791
R4325 VGND VGND.n1838 2.60791
R4326 VGND.n1835 VGND 2.60791
R4327 VGND VGND.n1834 2.60791
R4328 VGND.n1829 VGND 2.60791
R4329 VGND VGND.n1828 2.60791
R4330 VGND VGND.n1827 2.60791
R4331 VGND.n1823 VGND 2.60791
R4332 VGND.n1819 VGND 2.60791
R4333 VGND VGND.n1818 2.60791
R4334 VGND.n1815 VGND 2.60791
R4335 VGND.n1811 VGND 2.60791
R4336 VGND VGND.n1810 2.60791
R4337 VGND.n1807 VGND 2.60791
R4338 VGND.n1803 VGND 2.60791
R4339 VGND.n1799 VGND 2.60791
R4340 VGND.n1795 VGND 2.60791
R4341 VGND.n1791 VGND 2.60791
R4342 VGND.n1787 VGND 2.60791
R4343 VGND.n1031 VGND 2.60791
R4344 VGND.n1977 VGND 2.60791
R4345 VGND.n1980 VGND 2.60791
R4346 VGND VGND.n885 2.60791
R4347 VGND.n1987 VGND 2.60791
R4348 VGND VGND.n1986 2.60791
R4349 VGND.n917 VGND 2.60791
R4350 VGND.n921 VGND 2.60791
R4351 VGND.n922 VGND 2.60791
R4352 VGND.n926 VGND 2.60791
R4353 VGND.n929 VGND 2.60791
R4354 VGND.n930 VGND 2.60791
R4355 VGND.n933 VGND 2.60791
R4356 VGND.n934 VGND 2.60791
R4357 VGND.n937 VGND 2.60791
R4358 VGND.n938 VGND 2.60791
R4359 VGND.n941 VGND 2.60791
R4360 VGND.n942 VGND 2.60791
R4361 VGND.n945 VGND 2.60791
R4362 VGND.n946 VGND 2.60791
R4363 VGND.n949 VGND 2.60791
R4364 VGND.n950 VGND 2.60791
R4365 VGND.n953 VGND 2.60791
R4366 VGND.n954 VGND 2.60791
R4367 VGND.n957 VGND 2.60791
R4368 VGND.n958 VGND 2.60791
R4369 VGND.n961 VGND 2.60791
R4370 VGND.n962 VGND 2.60791
R4371 VGND.n965 VGND 2.60791
R4372 VGND.n966 VGND 2.60791
R4373 VGND.n969 VGND 2.60791
R4374 VGND.n970 VGND 2.60791
R4375 VGND.n973 VGND 2.60791
R4376 VGND.n974 VGND 2.60791
R4377 VGND.n977 VGND 2.60791
R4378 VGND.n978 VGND 2.60791
R4379 VGND.n981 VGND 2.60791
R4380 VGND.n982 VGND 2.60791
R4381 VGND.n985 VGND 2.60791
R4382 VGND.n986 VGND 2.60791
R4383 VGND.n989 VGND 2.60791
R4384 VGND.n990 VGND 2.60791
R4385 VGND.n993 VGND 2.60791
R4386 VGND.n994 VGND 2.60791
R4387 VGND.n997 VGND 2.60791
R4388 VGND.n998 VGND 2.60791
R4389 VGND.n1001 VGND 2.60791
R4390 VGND.n1005 VGND 2.60791
R4391 VGND.n1006 VGND 2.60791
R4392 VGND.n1009 VGND 2.60791
R4393 VGND.n1010 VGND 2.60791
R4394 VGND.n1013 VGND 2.60791
R4395 VGND.n1014 VGND 2.60791
R4396 VGND.n1015 VGND 2.60791
R4397 VGND.n2030 VGND 2.60791
R4398 VGND.n1098 VGND 2.60791
R4399 VGND.n1966 VGND 2.60791
R4400 VGND VGND.n1965 2.60791
R4401 VGND VGND.n1964 2.60791
R4402 VGND VGND.n1962 2.60791
R4403 VGND.n1959 VGND 2.60791
R4404 VGND VGND.n1958 2.60791
R4405 VGND.n1955 VGND 2.60791
R4406 VGND.n1951 VGND 2.60791
R4407 VGND.n1947 VGND 2.60791
R4408 VGND VGND.n1946 2.60791
R4409 VGND VGND.n1942 2.60791
R4410 VGND.n1939 VGND 2.60791
R4411 VGND.n1935 VGND 2.60791
R4412 VGND.n1931 VGND 2.60791
R4413 VGND VGND.n2370 2.60791
R4414 VGND.n2366 VGND 2.60791
R4415 VGND VGND.n2365 2.60791
R4416 VGND VGND.n2361 2.60791
R4417 VGND.n2358 VGND 2.60791
R4418 VGND.n2354 VGND 2.60791
R4419 VGND.n2350 VGND 2.60791
R4420 VGND VGND.n2349 2.60791
R4421 VGND VGND.n2345 2.60791
R4422 VGND.n2342 VGND 2.60791
R4423 VGND.n2338 VGND 2.60791
R4424 VGND.n2334 VGND 2.60791
R4425 VGND.n2374 VGND 2.60791
R4426 VGND VGND.n2330 2.60791
R4427 VGND.n774 VGND 2.60791
R4428 VGND.n2323 VGND 2.60791
R4429 VGND VGND.n2321 2.60791
R4430 VGND.n777 VGND 2.60791
R4431 VGND VGND.n2314 2.60791
R4432 VGND.n782 VGND 2.60791
R4433 VGND.n2307 VGND 2.60791
R4434 VGND VGND.n2305 2.60791
R4435 VGND.n785 VGND 2.60791
R4436 VGND VGND.n2298 2.60791
R4437 VGND.n789 VGND 2.60791
R4438 VGND.n2290 VGND 2.60791
R4439 VGND.n2197 VGND 2.60791
R4440 VGND VGND.n2196 2.60791
R4441 VGND VGND.n2192 2.60791
R4442 VGND VGND.n2188 2.60791
R4443 VGND.n2185 VGND 2.60791
R4444 VGND.n2181 VGND 2.60791
R4445 VGND.n2177 VGND 2.60791
R4446 VGND VGND.n2176 2.60791
R4447 VGND VGND.n2172 2.60791
R4448 VGND VGND.n2168 2.60791
R4449 VGND VGND.n2164 2.60791
R4450 VGND.n2161 VGND 2.60791
R4451 VGND VGND.n2160 2.60791
R4452 VGND.n2157 VGND 2.60791
R4453 VGND.n2153 VGND 2.60791
R4454 VGND VGND.n2152 2.60791
R4455 VGND.n2149 VGND 2.60791
R4456 VGND VGND.n2148 2.60791
R4457 VGND VGND.n2144 2.60791
R4458 VGND.n2141 VGND 2.60791
R4459 VGND VGND.n2140 2.60791
R4460 VGND.n2137 VGND 2.60791
R4461 VGND.n2133 VGND 2.60791
R4462 VGND VGND.n2132 2.60791
R4463 VGND.n2129 VGND 2.60791
R4464 VGND VGND.n2128 2.60791
R4465 VGND VGND.n2124 2.60791
R4466 VGND.n2121 VGND 2.60791
R4467 VGND VGND.n2120 2.60791
R4468 VGND.n2117 VGND 2.60791
R4469 VGND.n2113 VGND 2.60791
R4470 VGND VGND.n2112 2.60791
R4471 VGND.n2109 VGND 2.60791
R4472 VGND.n2105 VGND 2.60791
R4473 VGND VGND.n2104 2.60791
R4474 VGND.n2101 VGND 2.60791
R4475 VGND.n2097 VGND 2.60791
R4476 VGND.n2093 VGND 2.60791
R4477 VGND.n2089 VGND 2.60791
R4478 VGND.n2085 VGND 2.60791
R4479 VGND.n2081 VGND 2.60791
R4480 VGND.n2729 VGND 2.60791
R4481 VGND.n2723 VGND 2.60791
R4482 VGND VGND.n2722 2.60791
R4483 VGND.n87 VGND 2.60791
R4484 VGND VGND.n2714 2.60791
R4485 VGND VGND.n2713 2.60791
R4486 VGND.n2707 VGND 2.60791
R4487 VGND VGND.n2705 2.60791
R4488 VGND.n95 VGND 2.60791
R4489 VGND VGND.n2698 2.60791
R4490 VGND.n99 VGND 2.60791
R4491 VGND VGND.n2690 2.60791
R4492 VGND VGND.n2689 2.60791
R4493 VGND.n104 VGND 2.60791
R4494 VGND.n2683 VGND 2.60791
R4495 VGND VGND.n2681 2.60791
R4496 VGND.n107 VGND 2.60791
R4497 VGND.n2675 VGND 2.60791
R4498 VGND VGND.n2674 2.60791
R4499 VGND.n111 VGND 2.60791
R4500 VGND.n2667 VGND 2.60791
R4501 VGND VGND.n2666 2.60791
R4502 VGND VGND.n2665 2.60791
R4503 VGND.n2659 VGND 2.60791
R4504 VGND VGND.n2658 2.60791
R4505 VGND VGND.n2657 2.60791
R4506 VGND.n119 VGND 2.60791
R4507 VGND VGND.n2650 2.60791
R4508 VGND VGND.n2649 2.60791
R4509 VGND.n124 VGND 2.60791
R4510 VGND.n2643 VGND 2.60791
R4511 VGND VGND.n2641 2.60791
R4512 VGND.n128 VGND 2.60791
R4513 VGND.n2635 VGND 2.60791
R4514 VGND VGND.n2633 2.60791
R4515 VGND.n132 VGND 2.60791
R4516 VGND.n2627 VGND 2.60791
R4517 VGND VGND.n2625 2.60791
R4518 VGND.n2619 VGND 2.60791
R4519 VGND VGND.n2617 2.60791
R4520 VGND.n2611 VGND 2.60791
R4521 VGND VGND.n2609 2.60791
R4522 VGND VGND.n2603 2.60791
R4523 VGND.n600 VGND 2.60791
R4524 VGND.n603 VGND 2.60791
R4525 VGND.n612 VGND 2.60791
R4526 VGND.n616 VGND 2.60791
R4527 VGND.n620 VGND 2.60791
R4528 VGND.n624 VGND 2.60791
R4529 VGND.n625 VGND 2.60791
R4530 VGND.n629 VGND 2.60791
R4531 VGND.n632 VGND 2.60791
R4532 VGND.n633 VGND 2.60791
R4533 VGND.n637 VGND 2.60791
R4534 VGND.n641 VGND 2.60791
R4535 VGND VGND.n2442 2.60791
R4536 VGND.n551 VGND 2.60791
R4537 VGND.n554 VGND 2.60791
R4538 VGND.n558 VGND 2.60791
R4539 VGND.n562 VGND 2.60791
R4540 VGND.n566 VGND 2.60791
R4541 VGND.n570 VGND 2.60791
R4542 VGND VGND.n1071 2.60791
R4543 VGND.n1072 VGND 2.60791
R4544 VGND VGND.n1039 2.60791
R4545 VGND.n1080 VGND 2.60791
R4546 VGND.n1921 VGND.n1920 2.30157
R4547 VGND.n166 VGND.n165 2.27862
R4548 VGND.n520 VGND.n519 2.27862
R4549 VGND.n1921 VGND.n1122 2.27078
R4550 VGND.n838 VGND.n837 2.2505
R4551 VGND.n2278 VGND.n2277 2.2505
R4552 VGND.n1158 VGND.n1157 2.2505
R4553 VGND.n1436 VGND.n1435 2.2505
R4554 VGND.n1680 VGND.n1657 2.2505
R4555 VGND.n1691 VGND.n1690 2.2505
R4556 VGND.n1682 VGND.n1681 2.2505
R4557 VGND.n1686 VGND.n1685 2.2505
R4558 VGND.n734 VGND.n731 2.2505
R4559 VGND.n2387 VGND.n2386 2.2505
R4560 VGND.n1701 VGND.n1545 2.2505
R4561 VGND.n1544 VGND.n1543 2.2505
R4562 VGND.n1651 VGND.n1548 2.2505
R4563 VGND.n1654 VGND.n1653 2.2505
R4564 VGND.n1441 VGND.n1440 2.2505
R4565 VGND.n1912 VGND.n1911 2.2505
R4566 VGND.n1697 VGND.n1696 2.2505
R4567 VGND.n1695 VGND.n1547 2.2505
R4568 VGND.n844 VGND.n843 2.2505
R4569 VGND.n842 VGND.n841 2.2505
R4570 VGND.n1151 VGND.n1150 2.2505
R4571 VGND.n1155 VGND.n1154 2.2505
R4572 VGND.n155 VGND.n154 2.2505
R4573 VGND.n157 VGND.n156 2.2505
R4574 VGND.n2383 VGND.n737 2.2505
R4575 VGND.n2382 VGND.n2381 2.2505
R4576 VGND.n836 VGND.n808 2.2505
R4577 VGND.n2283 VGND.n2282 2.2505
R4578 VGND.n2530 VGND.n2529 2.2505
R4579 VGND.n2527 VGND.n144 2.2505
R4580 VGND.n2497 VGND 2.01531
R4581 VGND VGND.n541 2.01531
R4582 VGND.n2443 VGND 2.01531
R4583 VGND.n0 VGND.t2 1.87438
R4584 VGND.n7 VGND.n6 1.77204
R4585 VGND.n6 VGND.n5 1.77204
R4586 VGND.n5 VGND.n4 1.77204
R4587 VGND.n4 VGND.n3 1.77204
R4588 VGND.n3 VGND.n2 1.77204
R4589 VGND.n2 VGND.n1 1.77204
R4590 VGND.n1 VGND.n0 1.77204
R4591 VGND.n2381 VGND.n2380 1.69938
R4592 VGND.n145 VGND.n143 1.69107
R4593 VGND.n1684 VGND.n1683 1.68852
R4594 VGND.n1688 VGND.n1658 1.68852
R4595 VGND.n733 VGND.n732 1.68852
R4596 VGND.n1434 VGND.n1433 1.68852
R4597 VGND.n1910 VGND.n1909 1.68852
R4598 VGND.n1549 VGND.n1439 1.68852
R4599 VGND.n1699 VGND.n1698 1.68852
R4600 VGND.n1703 VGND.n1702 1.68852
R4601 VGND.n2070 VGND.n845 1.68852
R4602 VGND.n1153 VGND.n1152 1.68852
R4603 VGND.n1918 VGND.n1123 1.68852
R4604 VGND.n2764 VGND.n11 1.68852
R4605 VGND.n2280 VGND.n809 1.68852
R4606 VGND.n2276 VGND.n2275 1.68852
R4607 VGND.n2767 VGND.n7 1.63737
R4608 VGND VGND.n839 1.2612
R4609 VGND.n2767 VGND.n8 0.894125
R4610 VGND.n2072 VGND.n143 0.853
R4611 VGND.n2073 VGND.n2072 0.853
R4612 VGND.n2766 VGND.n2765 0.853
R4613 VGND.n1915 VGND.n1438 0.853
R4614 VGND.n1542 VGND.n9 0.853
R4615 VGND.n1915 VGND.n1914 0.853
R4616 VGND.n2072 VGND.n2071 0.853
R4617 VGND.n1917 VGND.n1916 0.853
R4618 VGND.n2498 VGND.n2497 0.593093
R4619 VGND.n664 VGND.n541 0.593093
R4620 VGND.n235 VGND.n234 0.485794
R4621 VGND.n236 VGND.n235 0.485794
R4622 VGND.n237 VGND.n236 0.485794
R4623 VGND.n238 VGND.n237 0.485794
R4624 VGND.n239 VGND.n238 0.485794
R4625 VGND.n240 VGND.n239 0.485794
R4626 VGND.n241 VGND.n240 0.485794
R4627 VGND.n242 VGND.n241 0.485794
R4628 VGND.n243 VGND.n242 0.485794
R4629 VGND.n244 VGND.n243 0.485794
R4630 VGND.n245 VGND.n244 0.485794
R4631 VGND.n246 VGND.n245 0.485794
R4632 VGND.n247 VGND.n246 0.485794
R4633 VGND.n248 VGND.n247 0.485794
R4634 VGND.n249 VGND.n248 0.485794
R4635 VGND.n250 VGND.n249 0.485794
R4636 VGND.n251 VGND.n250 0.485794
R4637 VGND.n252 VGND.n251 0.485794
R4638 VGND.n253 VGND.n252 0.485794
R4639 VGND.n254 VGND.n253 0.485794
R4640 VGND.n255 VGND.n254 0.485794
R4641 VGND.n256 VGND.n255 0.485794
R4642 VGND.n257 VGND.n256 0.485794
R4643 VGND.n258 VGND.n257 0.485794
R4644 VGND.n259 VGND.n258 0.485794
R4645 VGND.n260 VGND.n259 0.485794
R4646 VGND.n261 VGND.n260 0.485794
R4647 VGND.n262 VGND.n261 0.485794
R4648 VGND.n263 VGND.n262 0.485794
R4649 VGND.n266 VGND.n263 0.485794
R4650 VGND.n204 VGND.n203 0.485794
R4651 VGND.n205 VGND.n204 0.485794
R4652 VGND.n206 VGND.n205 0.485794
R4653 VGND.n207 VGND.n206 0.485794
R4654 VGND.n208 VGND.n207 0.485794
R4655 VGND.n209 VGND.n208 0.485794
R4656 VGND.n210 VGND.n209 0.485794
R4657 VGND.n211 VGND.n210 0.485794
R4658 VGND.n212 VGND.n211 0.485794
R4659 VGND.n213 VGND.n212 0.485794
R4660 VGND.n214 VGND.n213 0.485794
R4661 VGND.n215 VGND.n214 0.485794
R4662 VGND.n216 VGND.n215 0.485794
R4663 VGND.n217 VGND.n216 0.485794
R4664 VGND.n218 VGND.n217 0.485794
R4665 VGND.n219 VGND.n218 0.485794
R4666 VGND.n220 VGND.n219 0.485794
R4667 VGND.n221 VGND.n220 0.485794
R4668 VGND.n222 VGND.n221 0.485794
R4669 VGND.n223 VGND.n222 0.485794
R4670 VGND.n224 VGND.n223 0.485794
R4671 VGND.n225 VGND.n224 0.485794
R4672 VGND.n226 VGND.n225 0.485794
R4673 VGND.n227 VGND.n226 0.485794
R4674 VGND.n228 VGND.n227 0.485794
R4675 VGND.n229 VGND.n228 0.485794
R4676 VGND.n230 VGND.n229 0.485794
R4677 VGND.n231 VGND.n230 0.485794
R4678 VGND.n232 VGND.n231 0.485794
R4679 VGND.n233 VGND.n232 0.485794
R4680 VGND.n267 VGND.n233 0.485794
R4681 VGND.n300 VGND.n299 0.485794
R4682 VGND.n299 VGND.n298 0.485794
R4683 VGND.n298 VGND.n297 0.485794
R4684 VGND.n297 VGND.n296 0.485794
R4685 VGND.n296 VGND.n295 0.485794
R4686 VGND.n295 VGND.n294 0.485794
R4687 VGND.n294 VGND.n293 0.485794
R4688 VGND.n293 VGND.n292 0.485794
R4689 VGND.n292 VGND.n291 0.485794
R4690 VGND.n291 VGND.n290 0.485794
R4691 VGND.n290 VGND.n289 0.485794
R4692 VGND.n289 VGND.n288 0.485794
R4693 VGND.n288 VGND.n287 0.485794
R4694 VGND.n287 VGND.n286 0.485794
R4695 VGND.n286 VGND.n285 0.485794
R4696 VGND.n285 VGND.n284 0.485794
R4697 VGND.n284 VGND.n283 0.485794
R4698 VGND.n283 VGND.n282 0.485794
R4699 VGND.n282 VGND.n281 0.485794
R4700 VGND.n281 VGND.n280 0.485794
R4701 VGND.n280 VGND.n279 0.485794
R4702 VGND.n279 VGND.n278 0.485794
R4703 VGND.n278 VGND.n277 0.485794
R4704 VGND.n277 VGND.n276 0.485794
R4705 VGND.n276 VGND.n275 0.485794
R4706 VGND.n275 VGND.n274 0.485794
R4707 VGND.n274 VGND.n273 0.485794
R4708 VGND.n273 VGND.n272 0.485794
R4709 VGND.n272 VGND.n271 0.485794
R4710 VGND.n271 VGND.n270 0.485794
R4711 VGND.n270 VGND.n269 0.485794
R4712 VGND.n269 VGND.n268 0.485794
R4713 VGND.n201 VGND.n200 0.485794
R4714 VGND.n200 VGND.n199 0.485794
R4715 VGND.n199 VGND.n198 0.485794
R4716 VGND.n198 VGND.n197 0.485794
R4717 VGND.n197 VGND.n196 0.485794
R4718 VGND.n196 VGND.n195 0.485794
R4719 VGND.n195 VGND.n194 0.485794
R4720 VGND.n194 VGND.n193 0.485794
R4721 VGND.n193 VGND.n192 0.485794
R4722 VGND.n192 VGND.n191 0.485794
R4723 VGND.n191 VGND.n190 0.485794
R4724 VGND.n190 VGND.n189 0.485794
R4725 VGND.n189 VGND.n188 0.485794
R4726 VGND.n188 VGND.n187 0.485794
R4727 VGND.n187 VGND.n186 0.485794
R4728 VGND.n186 VGND.n185 0.485794
R4729 VGND.n185 VGND.n184 0.485794
R4730 VGND.n184 VGND.n183 0.485794
R4731 VGND.n183 VGND.n182 0.485794
R4732 VGND.n182 VGND.n181 0.485794
R4733 VGND.n181 VGND.n180 0.485794
R4734 VGND.n180 VGND.n179 0.485794
R4735 VGND.n179 VGND.n178 0.485794
R4736 VGND.n178 VGND.n177 0.485794
R4737 VGND.n177 VGND.n176 0.485794
R4738 VGND.n176 VGND.n175 0.485794
R4739 VGND.n175 VGND.n174 0.485794
R4740 VGND.n174 VGND.n173 0.485794
R4741 VGND.n173 VGND.n172 0.485794
R4742 VGND.n172 VGND.n171 0.485794
R4743 VGND.n171 VGND.n170 0.485794
R4744 VGND.n304 VGND.n303 0.485794
R4745 VGND.n305 VGND.n304 0.485794
R4746 VGND.n306 VGND.n305 0.485794
R4747 VGND.n307 VGND.n306 0.485794
R4748 VGND.n308 VGND.n307 0.485794
R4749 VGND.n309 VGND.n308 0.485794
R4750 VGND.n310 VGND.n309 0.485794
R4751 VGND.n311 VGND.n310 0.485794
R4752 VGND.n312 VGND.n311 0.485794
R4753 VGND.n313 VGND.n312 0.485794
R4754 VGND.n314 VGND.n313 0.485794
R4755 VGND.n315 VGND.n314 0.485794
R4756 VGND.n316 VGND.n315 0.485794
R4757 VGND.n317 VGND.n316 0.485794
R4758 VGND.n318 VGND.n317 0.485794
R4759 VGND.n319 VGND.n318 0.485794
R4760 VGND.n320 VGND.n319 0.485794
R4761 VGND.n321 VGND.n320 0.485794
R4762 VGND.n322 VGND.n321 0.485794
R4763 VGND.n323 VGND.n322 0.485794
R4764 VGND.n324 VGND.n323 0.485794
R4765 VGND.n325 VGND.n324 0.485794
R4766 VGND.n326 VGND.n325 0.485794
R4767 VGND.n327 VGND.n326 0.485794
R4768 VGND.n328 VGND.n327 0.485794
R4769 VGND.n329 VGND.n328 0.485794
R4770 VGND.n330 VGND.n329 0.485794
R4771 VGND.n331 VGND.n330 0.485794
R4772 VGND.n332 VGND.n331 0.485794
R4773 VGND.n333 VGND.n332 0.485794
R4774 VGND.n438 VGND.n437 0.485794
R4775 VGND.n439 VGND.n438 0.485794
R4776 VGND.n440 VGND.n439 0.485794
R4777 VGND.n441 VGND.n440 0.485794
R4778 VGND.n442 VGND.n441 0.485794
R4779 VGND.n443 VGND.n442 0.485794
R4780 VGND.n444 VGND.n443 0.485794
R4781 VGND.n445 VGND.n444 0.485794
R4782 VGND.n446 VGND.n445 0.485794
R4783 VGND.n447 VGND.n446 0.485794
R4784 VGND.n448 VGND.n447 0.485794
R4785 VGND.n449 VGND.n448 0.485794
R4786 VGND.n450 VGND.n449 0.485794
R4787 VGND.n451 VGND.n450 0.485794
R4788 VGND.n452 VGND.n451 0.485794
R4789 VGND.n453 VGND.n452 0.485794
R4790 VGND.n454 VGND.n453 0.485794
R4791 VGND.n455 VGND.n454 0.485794
R4792 VGND.n456 VGND.n455 0.485794
R4793 VGND.n457 VGND.n456 0.485794
R4794 VGND.n458 VGND.n457 0.485794
R4795 VGND.n459 VGND.n458 0.485794
R4796 VGND.n460 VGND.n459 0.485794
R4797 VGND.n461 VGND.n460 0.485794
R4798 VGND.n462 VGND.n461 0.485794
R4799 VGND.n463 VGND.n462 0.485794
R4800 VGND.n464 VGND.n463 0.485794
R4801 VGND.n465 VGND.n464 0.485794
R4802 VGND.n466 VGND.n465 0.485794
R4803 VGND.n467 VGND.n466 0.485794
R4804 VGND.n468 VGND.n467 0.485794
R4805 VGND.n469 VGND.n468 0.485794
R4806 VGND.n436 VGND.n435 0.485794
R4807 VGND.n435 VGND.n434 0.485794
R4808 VGND.n434 VGND.n433 0.485794
R4809 VGND.n433 VGND.n432 0.485794
R4810 VGND.n432 VGND.n431 0.485794
R4811 VGND.n431 VGND.n430 0.485794
R4812 VGND.n430 VGND.n429 0.485794
R4813 VGND.n429 VGND.n428 0.485794
R4814 VGND.n428 VGND.n427 0.485794
R4815 VGND.n427 VGND.n426 0.485794
R4816 VGND.n426 VGND.n425 0.485794
R4817 VGND.n425 VGND.n424 0.485794
R4818 VGND.n424 VGND.n423 0.485794
R4819 VGND.n423 VGND.n422 0.485794
R4820 VGND.n422 VGND.n421 0.485794
R4821 VGND.n421 VGND.n420 0.485794
R4822 VGND.n420 VGND.n419 0.485794
R4823 VGND.n419 VGND.n418 0.485794
R4824 VGND.n418 VGND.n417 0.485794
R4825 VGND.n417 VGND.n416 0.485794
R4826 VGND.n416 VGND.n415 0.485794
R4827 VGND.n415 VGND.n414 0.485794
R4828 VGND.n414 VGND.n413 0.485794
R4829 VGND.n413 VGND.n412 0.485794
R4830 VGND.n412 VGND.n411 0.485794
R4831 VGND.n411 VGND.n410 0.485794
R4832 VGND.n410 VGND.n409 0.485794
R4833 VGND.n409 VGND.n408 0.485794
R4834 VGND.n408 VGND.n407 0.485794
R4835 VGND.n407 VGND.n406 0.485794
R4836 VGND.n406 VGND.n404 0.485794
R4837 VGND.n470 VGND.n404 0.485794
R4838 VGND.n344 VGND.n337 0.485794
R4839 VGND.n346 VGND.n344 0.485794
R4840 VGND.n348 VGND.n346 0.485794
R4841 VGND.n350 VGND.n348 0.485794
R4842 VGND.n352 VGND.n350 0.485794
R4843 VGND.n354 VGND.n352 0.485794
R4844 VGND.n356 VGND.n354 0.485794
R4845 VGND.n358 VGND.n356 0.485794
R4846 VGND.n360 VGND.n358 0.485794
R4847 VGND.n362 VGND.n360 0.485794
R4848 VGND.n364 VGND.n362 0.485794
R4849 VGND.n366 VGND.n364 0.485794
R4850 VGND.n368 VGND.n366 0.485794
R4851 VGND.n370 VGND.n368 0.485794
R4852 VGND.n372 VGND.n370 0.485794
R4853 VGND.n374 VGND.n372 0.485794
R4854 VGND.n376 VGND.n374 0.485794
R4855 VGND.n378 VGND.n376 0.485794
R4856 VGND.n380 VGND.n378 0.485794
R4857 VGND.n382 VGND.n380 0.485794
R4858 VGND.n384 VGND.n382 0.485794
R4859 VGND.n386 VGND.n384 0.485794
R4860 VGND.n388 VGND.n386 0.485794
R4861 VGND.n390 VGND.n388 0.485794
R4862 VGND.n392 VGND.n390 0.485794
R4863 VGND.n394 VGND.n392 0.485794
R4864 VGND.n396 VGND.n394 0.485794
R4865 VGND.n398 VGND.n396 0.485794
R4866 VGND.n400 VGND.n398 0.485794
R4867 VGND.n402 VGND.n400 0.485794
R4868 VGND.n474 VGND.n402 0.485794
R4869 VGND.n474 VGND.n473 0.485794
R4870 VGND.n343 VGND.n342 0.485794
R4871 VGND.n345 VGND.n343 0.485794
R4872 VGND.n347 VGND.n345 0.485794
R4873 VGND.n349 VGND.n347 0.485794
R4874 VGND.n351 VGND.n349 0.485794
R4875 VGND.n353 VGND.n351 0.485794
R4876 VGND.n355 VGND.n353 0.485794
R4877 VGND.n357 VGND.n355 0.485794
R4878 VGND.n359 VGND.n357 0.485794
R4879 VGND.n361 VGND.n359 0.485794
R4880 VGND.n363 VGND.n361 0.485794
R4881 VGND.n365 VGND.n363 0.485794
R4882 VGND.n367 VGND.n365 0.485794
R4883 VGND.n369 VGND.n367 0.485794
R4884 VGND.n371 VGND.n369 0.485794
R4885 VGND.n373 VGND.n371 0.485794
R4886 VGND.n375 VGND.n373 0.485794
R4887 VGND.n377 VGND.n375 0.485794
R4888 VGND.n379 VGND.n377 0.485794
R4889 VGND.n381 VGND.n379 0.485794
R4890 VGND.n383 VGND.n381 0.485794
R4891 VGND.n385 VGND.n383 0.485794
R4892 VGND.n387 VGND.n385 0.485794
R4893 VGND.n389 VGND.n387 0.485794
R4894 VGND.n391 VGND.n389 0.485794
R4895 VGND.n393 VGND.n391 0.485794
R4896 VGND.n395 VGND.n393 0.485794
R4897 VGND.n397 VGND.n395 0.485794
R4898 VGND.n399 VGND.n397 0.485794
R4899 VGND.n401 VGND.n399 0.485794
R4900 VGND.n506 VGND.n505 0.485794
R4901 VGND.n505 VGND.n504 0.485794
R4902 VGND.n504 VGND.n503 0.485794
R4903 VGND.n503 VGND.n502 0.485794
R4904 VGND.n502 VGND.n501 0.485794
R4905 VGND.n501 VGND.n500 0.485794
R4906 VGND.n500 VGND.n499 0.485794
R4907 VGND.n499 VGND.n498 0.485794
R4908 VGND.n498 VGND.n497 0.485794
R4909 VGND.n497 VGND.n496 0.485794
R4910 VGND.n496 VGND.n495 0.485794
R4911 VGND.n495 VGND.n494 0.485794
R4912 VGND.n494 VGND.n493 0.485794
R4913 VGND.n493 VGND.n492 0.485794
R4914 VGND.n492 VGND.n491 0.485794
R4915 VGND.n491 VGND.n490 0.485794
R4916 VGND.n490 VGND.n489 0.485794
R4917 VGND.n489 VGND.n488 0.485794
R4918 VGND.n488 VGND.n487 0.485794
R4919 VGND.n487 VGND.n486 0.485794
R4920 VGND.n486 VGND.n485 0.485794
R4921 VGND.n485 VGND.n484 0.485794
R4922 VGND.n484 VGND.n483 0.485794
R4923 VGND.n483 VGND.n482 0.485794
R4924 VGND.n482 VGND.n481 0.485794
R4925 VGND.n481 VGND.n480 0.485794
R4926 VGND.n480 VGND.n479 0.485794
R4927 VGND.n479 VGND.n478 0.485794
R4928 VGND.n478 VGND.n477 0.485794
R4929 VGND.n477 VGND.n476 0.485794
R4930 VGND.n476 VGND.n475 0.485794
R4931 VGND.n302 VGND.n301 0.467912
R4932 VGND.n1688 VGND.n1687 0.414324
R4933 VGND.n738 VGND.n10 0.414124
R4934 VGND.n1700 VGND.n1699 0.413623
R4935 VGND.n2280 VGND.n2279 0.413122
R4936 VGND.n1438 VGND.n732 0.410318
R4937 VGND.n1914 VGND.n1439 0.410318
R4938 VGND.n1918 VGND.n1917 0.406661
R4939 VGND.n1152 VGND.n883 0.394891
R4940 VGND.n2003 VGND 0.337674
R4941 VGND.n2005 VGND 0.337674
R4942 VGND.n2021 VGND 0.337674
R4943 VGND.n2023 VGND 0.337674
R4944 VGND.n472 VGND.n403 0.243647
R4945 VGND.n437 VGND.n334 0.243147
R4946 VGND.n436 VGND.n335 0.243147
R4947 VGND.n523 VGND.n337 0.243147
R4948 VGND.n507 VGND.n506 0.243147
R4949 VGND.n203 VGND.n202 0.225833
R4950 VGND.n302 VGND.n201 0.225833
R4951 VGND.n475 VGND.n403 0.225833
R4952 VGND.n471 VGND.n470 0.224765
R4953 VGND.n2521 VGND.n2520 0.191676
R4954 VGND.n2519 VGND.n167 0.191676
R4955 VGND.n265 VGND.n161 0.191676
R4956 VGND.n2522 VGND.n162 0.191676
R4957 VGND.n2518 VGND.n2517 0.191676
R4958 VGND.n2515 VGND.n2511 0.191676
R4959 VGND.n513 VGND.n336 0.191676
R4960 VGND.n515 VGND.n514 0.191676
R4961 VGND.n522 VGND.n338 0.191676
R4962 VGND.n521 VGND.n339 0.191676
R4963 VGND.n517 VGND.n340 0.191676
R4964 VGND.n508 VGND.n341 0.191676
R4965 VGND.n267 VGND 0.180647
R4966 VGND.n268 VGND 0.180647
R4967 VGND.n170 VGND 0.180647
R4968 VGND VGND.n333 0.180647
R4969 VGND.n2070 VGND.n2069 0.170109
R4970 VGND.n2532 VGND.n2531 0.170109
R4971 VGND.n1433 VGND.n1432 0.169658
R4972 VGND.n1704 VGND.n1703 0.169157
R4973 VGND.n2275 VGND.n2274 0.169157
R4974 VGND.n2764 VGND.n2763 0.166653
R4975 VGND.n1909 VGND.n1908 0.163147
R4976 VGND VGND.n1248 0.157848
R4977 VGND VGND.n1247 0.157848
R4978 VGND VGND.n1409 0.157848
R4979 VGND VGND.n1408 0.157848
R4980 VGND.n1522 VGND 0.157848
R4981 VGND.n1524 VGND 0.157848
R4982 VGND.n1763 VGND 0.157848
R4983 VGND.n1765 VGND 0.157848
R4984 VGND VGND.n2046 0.157848
R4985 VGND VGND.n2045 0.157848
R4986 VGND VGND.n2740 0.157848
R4987 VGND VGND.n2739 0.157848
R4988 VGND VGND.n2251 0.157848
R4989 VGND VGND.n2250 0.157848
R4990 VGND.n2586 VGND 0.157848
R4991 VGND.n2588 VGND 0.157848
R4992 VGND.n1244 VGND.n1243 0.13537
R4993 VGND.n1405 VGND.n1404 0.13537
R4994 VGND.n1532 VGND.n1530 0.13537
R4995 VGND.n1773 VGND.n1771 0.13537
R4996 VGND.n2042 VGND.n2041 0.13537
R4997 VGND.n2736 VGND.n2735 0.13537
R4998 VGND.n2247 VGND.n2246 0.13537
R4999 VGND.n2596 VGND.n2594 0.13537
R5000 VGND.n1204 VGND.n8 0.117489
R5001 VGND VGND.n2459 0.112891
R5002 VGND VGND.n2458 0.112891
R5003 VGND VGND.n1265 0.112891
R5004 VGND VGND.n1262 0.112891
R5005 VGND.n1243 VGND 0.112891
R5006 VGND.n1661 VGND 0.112891
R5007 VGND.n1663 VGND 0.112891
R5008 VGND.n1667 VGND 0.112891
R5009 VGND.n1669 VGND 0.112891
R5010 VGND.n715 VGND 0.112891
R5011 VGND.n717 VGND 0.112891
R5012 VGND.n721 VGND 0.112891
R5013 VGND.n723 VGND 0.112891
R5014 VGND VGND.n1426 0.112891
R5015 VGND VGND.n1423 0.112891
R5016 VGND.n1404 VGND 0.112891
R5017 VGND.n1483 VGND 0.112891
R5018 VGND.n1490 VGND 0.112891
R5019 VGND VGND.n1532 0.112891
R5020 VGND.n1552 VGND 0.112891
R5021 VGND.n1554 VGND 0.112891
R5022 VGND.n1558 VGND 0.112891
R5023 VGND.n1560 VGND 0.112891
R5024 VGND.n1623 VGND 0.112891
R5025 VGND.n1625 VGND 0.112891
R5026 VGND.n1629 VGND 0.112891
R5027 VGND.n1631 VGND 0.112891
R5028 VGND.n1724 VGND 0.112891
R5029 VGND.n1731 VGND 0.112891
R5030 VGND VGND.n1773 0.112891
R5031 VGND VGND.n2063 0.112891
R5032 VGND VGND.n2060 0.112891
R5033 VGND.n2041 VGND 0.112891
R5034 VGND.n1999 VGND 0.112891
R5035 VGND.n1128 VGND 0.112891
R5036 VGND.n1104 VGND 0.112891
R5037 VGND.n1106 VGND 0.112891
R5038 VGND.n1110 VGND 0.112891
R5039 VGND.n1112 VGND 0.112891
R5040 VGND VGND.n2757 0.112891
R5041 VGND VGND.n2754 0.112891
R5042 VGND.n2735 VGND 0.112891
R5043 VGND.n741 VGND 0.112891
R5044 VGND.n743 VGND 0.112891
R5045 VGND.n747 VGND 0.112891
R5046 VGND.n749 VGND 0.112891
R5047 VGND.n792 VGND 0.112891
R5048 VGND.n794 VGND 0.112891
R5049 VGND.n798 VGND 0.112891
R5050 VGND.n800 VGND 0.112891
R5051 VGND.n812 VGND 0.112891
R5052 VGND.n814 VGND 0.112891
R5053 VGND.n818 VGND 0.112891
R5054 VGND.n820 VGND 0.112891
R5055 VGND VGND.n2268 0.112891
R5056 VGND VGND.n2265 0.112891
R5057 VGND.n2246 VGND 0.112891
R5058 VGND.n2547 VGND 0.112891
R5059 VGND.n2554 VGND 0.112891
R5060 VGND VGND.n2596 0.112891
R5061 VGND VGND.n654 0.112891
R5062 VGND VGND.n653 0.112891
R5063 VGND.n7 VGND.t7 0.102843
R5064 VGND.n6 VGND.t8 0.102843
R5065 VGND.n5 VGND.t3 0.102843
R5066 VGND.n4 VGND.t1 0.102843
R5067 VGND.n3 VGND.t4 0.102843
R5068 VGND.n2 VGND.t6 0.102843
R5069 VGND.n1 VGND.t5 0.102843
R5070 VGND.n0 VGND.t0 0.102843
R5071 VGND.n264 VGND.n163 0.0930382
R5072 VGND.n2514 VGND.n2513 0.0930382
R5073 VGND.n516 VGND.n512 0.0930382
R5074 VGND.n510 VGND.n509 0.0930382
R5075 VGND.n1689 VGND 0.0914348
R5076 VGND VGND.n2388 0.0914348
R5077 VGND.n1652 VGND 0.0914348
R5078 VGND VGND.n1546 0.0914348
R5079 VGND.n2379 VGND 0.0914348
R5080 VGND.n2281 VGND 0.0914348
R5081 VGND.n1268 VGND.n1267 0.090413
R5082 VGND.n1262 VGND.n1261 0.090413
R5083 VGND.n1260 VGND.n1259 0.090413
R5084 VGND.n1259 VGND.n1258 0.090413
R5085 VGND.n1257 VGND.n1256 0.090413
R5086 VGND.n1256 VGND.n1255 0.090413
R5087 VGND.n1254 VGND.n1253 0.090413
R5088 VGND.n1253 VGND.n1252 0.090413
R5089 VGND.n1251 VGND.n1250 0.090413
R5090 VGND.n1250 VGND.n1249 0.090413
R5091 VGND.n1429 VGND.n1428 0.090413
R5092 VGND.n1423 VGND.n1422 0.090413
R5093 VGND.n1421 VGND.n1420 0.090413
R5094 VGND.n1420 VGND.n1419 0.090413
R5095 VGND.n1418 VGND.n1417 0.090413
R5096 VGND.n1417 VGND.n1416 0.090413
R5097 VGND.n1415 VGND.n1414 0.090413
R5098 VGND.n1414 VGND.n1413 0.090413
R5099 VGND.n1412 VGND.n1411 0.090413
R5100 VGND.n1411 VGND.n1410 0.090413
R5101 VGND.n1479 VGND.n1477 0.090413
R5102 VGND.n1492 VGND.n1490 0.090413
R5103 VGND.n1497 VGND.n1494 0.090413
R5104 VGND.n1499 VGND.n1497 0.090413
R5105 VGND.n1504 VGND.n1501 0.090413
R5106 VGND.n1506 VGND.n1504 0.090413
R5107 VGND.n1511 VGND.n1508 0.090413
R5108 VGND.n1513 VGND.n1511 0.090413
R5109 VGND.n1518 VGND.n1515 0.090413
R5110 VGND.n1520 VGND.n1518 0.090413
R5111 VGND.n1720 VGND.n1718 0.090413
R5112 VGND.n1733 VGND.n1731 0.090413
R5113 VGND.n1738 VGND.n1735 0.090413
R5114 VGND.n1740 VGND.n1738 0.090413
R5115 VGND.n1745 VGND.n1742 0.090413
R5116 VGND.n1747 VGND.n1745 0.090413
R5117 VGND.n1752 VGND.n1749 0.090413
R5118 VGND.n1754 VGND.n1752 0.090413
R5119 VGND.n1759 VGND.n1756 0.090413
R5120 VGND.n1761 VGND.n1759 0.090413
R5121 VGND.n2066 VGND.n2065 0.090413
R5122 VGND.n2060 VGND.n2059 0.090413
R5123 VGND.n2058 VGND.n2057 0.090413
R5124 VGND.n2057 VGND.n2056 0.090413
R5125 VGND.n2055 VGND.n2054 0.090413
R5126 VGND.n2054 VGND.n2053 0.090413
R5127 VGND.n2052 VGND.n2051 0.090413
R5128 VGND.n2051 VGND.n2050 0.090413
R5129 VGND.n2049 VGND.n2048 0.090413
R5130 VGND.n2048 VGND.n2047 0.090413
R5131 VGND.n1997 VGND.n1995 0.090413
R5132 VGND.n2010 VGND.n2007 0.090413
R5133 VGND.n2012 VGND.n2010 0.090413
R5134 VGND.n2017 VGND.n2014 0.090413
R5135 VGND.n2019 VGND.n2017 0.090413
R5136 VGND.n1136 VGND.n1134 0.090413
R5137 VGND.n2760 VGND.n2759 0.090413
R5138 VGND.n2754 VGND.n2753 0.090413
R5139 VGND.n2752 VGND.n2751 0.090413
R5140 VGND.n2751 VGND.n2750 0.090413
R5141 VGND.n2749 VGND.n2748 0.090413
R5142 VGND.n2748 VGND.n2747 0.090413
R5143 VGND.n2746 VGND.n2745 0.090413
R5144 VGND.n2745 VGND.n2744 0.090413
R5145 VGND.n2743 VGND.n2742 0.090413
R5146 VGND.n2742 VGND.n2741 0.090413
R5147 VGND.n2271 VGND.n2270 0.090413
R5148 VGND.n2265 VGND.n2264 0.090413
R5149 VGND.n2263 VGND.n2262 0.090413
R5150 VGND.n2262 VGND.n2261 0.090413
R5151 VGND.n2260 VGND.n2259 0.090413
R5152 VGND.n2259 VGND.n2258 0.090413
R5153 VGND.n2257 VGND.n2256 0.090413
R5154 VGND.n2256 VGND.n2255 0.090413
R5155 VGND.n2254 VGND.n2253 0.090413
R5156 VGND.n2253 VGND.n2252 0.090413
R5157 VGND.n2543 VGND.n2541 0.090413
R5158 VGND.n2556 VGND.n2554 0.090413
R5159 VGND.n2561 VGND.n2558 0.090413
R5160 VGND.n2563 VGND.n2561 0.090413
R5161 VGND.n2568 VGND.n2565 0.090413
R5162 VGND.n2570 VGND.n2568 0.090413
R5163 VGND.n2575 VGND.n2572 0.090413
R5164 VGND.n2577 VGND.n2575 0.090413
R5165 VGND.n2582 VGND.n2579 0.090413
R5166 VGND.n2584 VGND.n2582 0.090413
R5167 VGND.n1919 VGND 0.0860757
R5168 VGND.n165 VGND.n164 0.0723824
R5169 VGND.n2512 VGND.n166 0.0723824
R5170 VGND.n520 VGND.n511 0.0723824
R5171 VGND.n519 VGND.n518 0.0723824
R5172 VGND.n1691 VGND.n1657 0.0711522
R5173 VGND.n2386 VGND.n734 0.0711522
R5174 VGND.n1654 VGND.n1548 0.0711522
R5175 VGND.n1696 VGND.n1695 0.0711522
R5176 VGND.n157 VGND.n155 0.0711522
R5177 VGND.n2381 VGND.n737 0.0711522
R5178 VGND.n2383 VGND.n2382 0.0711522
R5179 VGND.n2283 VGND.n808 0.0711522
R5180 VGND.n2450 VGND 0.0679348
R5181 VGND VGND.n2460 0.0679348
R5182 VGND.n2458 VGND 0.0679348
R5183 VGND VGND.n2457 0.0679348
R5184 VGND VGND.n1269 0.0679348
R5185 VGND VGND.n1266 0.0679348
R5186 VGND VGND.n1264 0.0679348
R5187 VGND VGND.n1263 0.0679348
R5188 VGND VGND.n1246 0.0679348
R5189 VGND VGND.n1245 0.0679348
R5190 VGND.n1665 VGND 0.0679348
R5191 VGND.n1671 VGND 0.0679348
R5192 VGND.n1673 VGND 0.0679348
R5193 VGND.n719 VGND 0.0679348
R5194 VGND.n725 VGND 0.0679348
R5195 VGND.n727 VGND 0.0679348
R5196 VGND VGND.n1430 0.0679348
R5197 VGND VGND.n1427 0.0679348
R5198 VGND VGND.n1425 0.0679348
R5199 VGND VGND.n1424 0.0679348
R5200 VGND VGND.n1407 0.0679348
R5201 VGND VGND.n1406 0.0679348
R5202 VGND.n1475 VGND 0.0679348
R5203 VGND.n1481 VGND 0.0679348
R5204 VGND.n1485 VGND 0.0679348
R5205 VGND.n1487 VGND 0.0679348
R5206 VGND.n1526 VGND 0.0679348
R5207 VGND.n1528 VGND 0.0679348
R5208 VGND.n1556 VGND 0.0679348
R5209 VGND.n1562 VGND 0.0679348
R5210 VGND.n1564 VGND 0.0679348
R5211 VGND.n1627 VGND 0.0679348
R5212 VGND.n1633 VGND 0.0679348
R5213 VGND.n1635 VGND 0.0679348
R5214 VGND.n1716 VGND 0.0679348
R5215 VGND.n1722 VGND 0.0679348
R5216 VGND.n1726 VGND 0.0679348
R5217 VGND.n1728 VGND 0.0679348
R5218 VGND.n1767 VGND 0.0679348
R5219 VGND.n1769 VGND 0.0679348
R5220 VGND VGND.n2067 0.0679348
R5221 VGND VGND.n2064 0.0679348
R5222 VGND VGND.n2062 0.0679348
R5223 VGND VGND.n2061 0.0679348
R5224 VGND VGND.n2044 0.0679348
R5225 VGND VGND.n2043 0.0679348
R5226 VGND.n1993 VGND 0.0679348
R5227 VGND.n2001 VGND 0.0679348
R5228 VGND.n1126 VGND 0.0679348
R5229 VGND.n1130 VGND 0.0679348
R5230 VGND.n1132 VGND 0.0679348
R5231 VGND.n1139 VGND 0.0679348
R5232 VGND VGND.n1139 0.0679348
R5233 VGND.n1141 VGND 0.0679348
R5234 VGND.n1143 VGND 0.0679348
R5235 VGND.n1108 VGND 0.0679348
R5236 VGND.n1114 VGND 0.0679348
R5237 VGND.n1116 VGND 0.0679348
R5238 VGND VGND.n2761 0.0679348
R5239 VGND VGND.n2758 0.0679348
R5240 VGND VGND.n2756 0.0679348
R5241 VGND VGND.n2755 0.0679348
R5242 VGND VGND.n2738 0.0679348
R5243 VGND VGND.n2737 0.0679348
R5244 VGND.n745 VGND 0.0679348
R5245 VGND.n751 VGND 0.0679348
R5246 VGND.n753 VGND 0.0679348
R5247 VGND.n796 VGND 0.0679348
R5248 VGND.n802 VGND 0.0679348
R5249 VGND.n804 VGND 0.0679348
R5250 VGND.n816 VGND 0.0679348
R5251 VGND.n822 VGND 0.0679348
R5252 VGND.n824 VGND 0.0679348
R5253 VGND VGND.n2272 0.0679348
R5254 VGND VGND.n2269 0.0679348
R5255 VGND VGND.n2267 0.0679348
R5256 VGND VGND.n2266 0.0679348
R5257 VGND VGND.n2249 0.0679348
R5258 VGND VGND.n2248 0.0679348
R5259 VGND.n2539 VGND 0.0679348
R5260 VGND.n2545 VGND 0.0679348
R5261 VGND.n2549 VGND 0.0679348
R5262 VGND.n2551 VGND 0.0679348
R5263 VGND.n2590 VGND 0.0679348
R5264 VGND.n2592 VGND 0.0679348
R5265 VGND VGND.n658 0.0679348
R5266 VGND VGND.n655 0.0679348
R5267 VGND.n653 VGND 0.0679348
R5268 VGND VGND.n652 0.0679348
R5269 VGND.n1055 VGND 0.06442
R5270 VGND.n2523 VGND 0.063
R5271 VGND VGND.n168 0.063
R5272 VGND.n2516 VGND 0.063
R5273 VGND.n2510 VGND 0.063
R5274 VGND.n469 VGND 0.063
R5275 VGND.n470 VGND 0.063
R5276 VGND.n473 VGND 0.063
R5277 VGND.n472 VGND 0.063
R5278 VGND VGND.n1065 0.06066
R5279 VGND VGND.n1060 0.06066
R5280 VGND VGND.n2767 0.0585758
R5281 VGND.n1683 VGND.n8 0.0511662
R5282 VGND.n2462 VGND.n2461 0.0454565
R5283 VGND.n2506 VGND.n528 0.0454565
R5284 VGND.n1270 VGND.n1204 0.0454565
R5285 VGND.n1245 VGND.n1244 0.0454565
R5286 VGND.n1242 VGND.n1241 0.0454565
R5287 VGND.n1679 VGND.n1674 0.0454565
R5288 VGND.n2390 VGND.n2389 0.0454565
R5289 VGND.n1432 VGND.n1431 0.0454565
R5290 VGND.n1406 VGND.n1405 0.0454565
R5291 VGND.n1403 VGND.n1402 0.0454565
R5292 VGND.n1908 VGND.n1442 0.0454565
R5293 VGND.n1530 VGND.n1528 0.0454565
R5294 VGND.n1535 VGND.n1534 0.0454565
R5295 VGND.n1650 VGND.n1565 0.0454565
R5296 VGND.n1640 VGND.n1639 0.0454565
R5297 VGND.n1714 VGND.n1704 0.0454565
R5298 VGND.n1771 VGND.n1769 0.0454565
R5299 VGND.n1778 VGND.n1777 0.0454565
R5300 VGND.n2069 VGND.n2068 0.0454565
R5301 VGND.n2043 VGND.n2042 0.0454565
R5302 VGND.n2040 VGND.n2039 0.0454565
R5303 VGND.n1991 VGND.n883 0.0454565
R5304 VGND.n2026 VGND.n2025 0.0454565
R5305 VGND.n1149 VGND.n1144 0.0454565
R5306 VGND.n1923 VGND.n1120 0.0454565
R5307 VGND.n2763 VGND.n2762 0.0454565
R5308 VGND.n2737 VGND.n2736 0.0454565
R5309 VGND.n2734 VGND.n2733 0.0454565
R5310 VGND.n2378 VGND.n754 0.0454565
R5311 VGND.n2286 VGND.n806 0.0454565
R5312 VGND.n835 VGND.n825 0.0454565
R5313 VGND.n2274 VGND.n2273 0.0454565
R5314 VGND.n2248 VGND.n2247 0.0454565
R5315 VGND.n2245 VGND.n2244 0.0454565
R5316 VGND.n2537 VGND.n2532 0.0454565
R5317 VGND.n2594 VGND.n2592 0.0454565
R5318 VGND.n2599 VGND.n2598 0.0454565
R5319 VGND.n657 VGND.n656 0.0454565
R5320 VGND.n651 VGND.n650 0.0454565
R5321 VGND.n1060 VGND.n1055 0.04186
R5322 VGND.n2277 VGND.n158 0.0361924
R5323 VGND.n1435 VGND.n153 0.0361924
R5324 VGND.n1685 VGND.n152 0.0361924
R5325 VGND.n1543 VGND.n151 0.0361924
R5326 VGND.n1911 VGND.n150 0.0361924
R5327 VGND.n841 VGND.n149 0.0361924
R5328 VGND.n1154 VGND.n148 0.0361924
R5329 VGND.n2528 VGND.n2527 0.0361924
R5330 VGND.n2529 VGND.n2528 0.0361924
R5331 VGND.n837 VGND.n158 0.0361924
R5332 VGND.n1157 VGND.n153 0.0361924
R5333 VGND.n1681 VGND.n152 0.0361924
R5334 VGND.n1545 VGND.n151 0.0361924
R5335 VGND.n1440 VGND.n150 0.0361924
R5336 VGND.n843 VGND.n149 0.0361924
R5337 VGND.n1150 VGND.n148 0.0361924
R5338 VGND.n2278 VGND.n2276 0.0359639
R5339 VGND.n1123 VGND.n1122 0.0359639
R5340 VGND.n1436 VGND.n1434 0.0359639
R5341 VGND.n1690 VGND.n1658 0.0359639
R5342 VGND.n1686 VGND.n1684 0.0359639
R5343 VGND.n1684 VGND.n1682 0.0359639
R5344 VGND.n1680 VGND.n1658 0.0359639
R5345 VGND.n2387 VGND.n733 0.0359639
R5346 VGND.n733 VGND.n731 0.0359639
R5347 VGND.n1434 VGND.n1158 0.0359639
R5348 VGND.n1702 VGND.n1544 0.0359639
R5349 VGND.n1653 VGND.n1549 0.0359639
R5350 VGND.n1912 VGND.n1910 0.0359639
R5351 VGND.n1910 VGND.n1441 0.0359639
R5352 VGND.n1651 VGND.n1549 0.0359639
R5353 VGND.n1698 VGND.n1547 0.0359639
R5354 VGND.n1698 VGND.n1697 0.0359639
R5355 VGND.n1702 VGND.n1701 0.0359639
R5356 VGND.n845 VGND.n842 0.0359639
R5357 VGND.n845 VGND.n844 0.0359639
R5358 VGND.n1155 VGND.n1153 0.0359639
R5359 VGND.n1153 VGND.n1151 0.0359639
R5360 VGND.n1920 VGND.n1123 0.0359639
R5361 VGND.n156 VGND.n11 0.0359639
R5362 VGND.n154 VGND.n11 0.0359639
R5363 VGND.n2282 VGND.n809 0.0359639
R5364 VGND.n836 VGND.n809 0.0359639
R5365 VGND.n2276 VGND.n838 0.0359639
R5366 VGND.n145 VGND.n144 0.0359639
R5367 VGND.n2530 VGND.n145 0.0359639
R5368 VGND.n2526 VGND.n147 0.0282702
R5369 VGND.n147 VGND.n146 0.0282702
R5370 VGND.n1689 VGND.n1688 0.0270652
R5371 VGND.n2388 VGND.n732 0.0270652
R5372 VGND.n1652 VGND.n1439 0.0270652
R5373 VGND.n1699 VGND.n1546 0.0270652
R5374 VGND.n1156 VGND.n1152 0.0270652
R5375 VGND.n2281 VGND.n2280 0.0270652
R5376 VGND.n2071 VGND.n2070 0.0245109
R5377 VGND.n2531 VGND.n143 0.0245109
R5378 VGND.n1687 VGND.n1683 0.0244608
R5379 VGND.n1437 VGND.n1433 0.0244608
R5380 VGND.n1913 VGND.n1909 0.0244608
R5381 VGND.n1919 VGND.n1918 0.0244608
R5382 VGND.n1066 VGND 0.02306
R5383 VGND.n1065 VGND 0.02306
R5384 VGND VGND.n2448 0.0229783
R5385 VGND VGND.n2450 0.0229783
R5386 VGND.n2462 VGND 0.0229783
R5387 VGND.n2461 VGND 0.0229783
R5388 VGND.n2460 VGND 0.0229783
R5389 VGND.n2459 VGND 0.0229783
R5390 VGND.n2457 VGND 0.0229783
R5391 VGND VGND.n528 0.0229783
R5392 VGND VGND.n2506 0.0229783
R5393 VGND.n1270 VGND 0.0229783
R5394 VGND.n1269 VGND 0.0229783
R5395 VGND VGND.n1268 0.0229783
R5396 VGND.n1267 VGND 0.0229783
R5397 VGND.n1266 VGND 0.0229783
R5398 VGND.n1265 VGND 0.0229783
R5399 VGND.n1264 VGND 0.0229783
R5400 VGND.n1263 VGND 0.0229783
R5401 VGND.n1261 VGND 0.0229783
R5402 VGND VGND.n1260 0.0229783
R5403 VGND.n1258 VGND 0.0229783
R5404 VGND VGND.n1257 0.0229783
R5405 VGND.n1255 VGND 0.0229783
R5406 VGND VGND.n1254 0.0229783
R5407 VGND.n1252 VGND 0.0229783
R5408 VGND VGND.n1251 0.0229783
R5409 VGND.n1249 VGND 0.0229783
R5410 VGND.n1248 VGND 0.0229783
R5411 VGND.n1247 VGND 0.0229783
R5412 VGND.n1246 VGND 0.0229783
R5413 VGND VGND.n1242 0.0229783
R5414 VGND.n1241 VGND 0.0229783
R5415 VGND VGND.n1661 0.0229783
R5416 VGND VGND.n1663 0.0229783
R5417 VGND VGND.n1665 0.0229783
R5418 VGND VGND.n1667 0.0229783
R5419 VGND VGND.n1669 0.0229783
R5420 VGND VGND.n1671 0.0229783
R5421 VGND VGND.n1673 0.0229783
R5422 VGND.n1674 VGND 0.0229783
R5423 VGND VGND.n1679 0.0229783
R5424 VGND VGND.n715 0.0229783
R5425 VGND VGND.n717 0.0229783
R5426 VGND VGND.n719 0.0229783
R5427 VGND VGND.n721 0.0229783
R5428 VGND VGND.n723 0.0229783
R5429 VGND VGND.n725 0.0229783
R5430 VGND VGND.n727 0.0229783
R5431 VGND.n2390 VGND 0.0229783
R5432 VGND.n2389 VGND 0.0229783
R5433 VGND.n1431 VGND 0.0229783
R5434 VGND.n1430 VGND 0.0229783
R5435 VGND VGND.n1429 0.0229783
R5436 VGND.n1428 VGND 0.0229783
R5437 VGND.n1427 VGND 0.0229783
R5438 VGND.n1426 VGND 0.0229783
R5439 VGND.n1425 VGND 0.0229783
R5440 VGND.n1424 VGND 0.0229783
R5441 VGND.n1422 VGND 0.0229783
R5442 VGND VGND.n1421 0.0229783
R5443 VGND.n1419 VGND 0.0229783
R5444 VGND VGND.n1418 0.0229783
R5445 VGND.n1416 VGND 0.0229783
R5446 VGND VGND.n1415 0.0229783
R5447 VGND.n1413 VGND 0.0229783
R5448 VGND VGND.n1412 0.0229783
R5449 VGND.n1410 VGND 0.0229783
R5450 VGND.n1409 VGND 0.0229783
R5451 VGND.n1408 VGND 0.0229783
R5452 VGND.n1407 VGND 0.0229783
R5453 VGND VGND.n1403 0.0229783
R5454 VGND.n1402 VGND 0.0229783
R5455 VGND VGND.n1442 0.0229783
R5456 VGND VGND.n1475 0.0229783
R5457 VGND.n1477 VGND 0.0229783
R5458 VGND VGND.n1479 0.0229783
R5459 VGND VGND.n1481 0.0229783
R5460 VGND VGND.n1483 0.0229783
R5461 VGND VGND.n1485 0.0229783
R5462 VGND VGND.n1487 0.0229783
R5463 VGND VGND.n1492 0.0229783
R5464 VGND.n1494 VGND 0.0229783
R5465 VGND VGND.n1499 0.0229783
R5466 VGND.n1501 VGND 0.0229783
R5467 VGND VGND.n1506 0.0229783
R5468 VGND.n1508 VGND 0.0229783
R5469 VGND VGND.n1513 0.0229783
R5470 VGND.n1515 VGND 0.0229783
R5471 VGND VGND.n1520 0.0229783
R5472 VGND VGND.n1522 0.0229783
R5473 VGND VGND.n1524 0.0229783
R5474 VGND VGND.n1526 0.0229783
R5475 VGND.n1535 VGND 0.0229783
R5476 VGND.n1534 VGND 0.0229783
R5477 VGND VGND.n1552 0.0229783
R5478 VGND VGND.n1554 0.0229783
R5479 VGND VGND.n1556 0.0229783
R5480 VGND VGND.n1558 0.0229783
R5481 VGND VGND.n1560 0.0229783
R5482 VGND VGND.n1562 0.0229783
R5483 VGND VGND.n1564 0.0229783
R5484 VGND.n1565 VGND 0.0229783
R5485 VGND VGND.n1650 0.0229783
R5486 VGND VGND.n1623 0.0229783
R5487 VGND VGND.n1625 0.0229783
R5488 VGND VGND.n1627 0.0229783
R5489 VGND VGND.n1629 0.0229783
R5490 VGND VGND.n1631 0.0229783
R5491 VGND VGND.n1633 0.0229783
R5492 VGND VGND.n1635 0.0229783
R5493 VGND.n1640 VGND 0.0229783
R5494 VGND.n1639 VGND 0.0229783
R5495 VGND VGND.n1714 0.0229783
R5496 VGND VGND.n1716 0.0229783
R5497 VGND.n1718 VGND 0.0229783
R5498 VGND VGND.n1720 0.0229783
R5499 VGND VGND.n1722 0.0229783
R5500 VGND VGND.n1724 0.0229783
R5501 VGND VGND.n1726 0.0229783
R5502 VGND VGND.n1728 0.0229783
R5503 VGND VGND.n1733 0.0229783
R5504 VGND.n1735 VGND 0.0229783
R5505 VGND VGND.n1740 0.0229783
R5506 VGND.n1742 VGND 0.0229783
R5507 VGND VGND.n1747 0.0229783
R5508 VGND.n1749 VGND 0.0229783
R5509 VGND VGND.n1754 0.0229783
R5510 VGND.n1756 VGND 0.0229783
R5511 VGND VGND.n1761 0.0229783
R5512 VGND VGND.n1763 0.0229783
R5513 VGND VGND.n1765 0.0229783
R5514 VGND VGND.n1767 0.0229783
R5515 VGND.n1777 VGND 0.0229783
R5516 VGND.n1778 VGND 0.0229783
R5517 VGND.n2068 VGND 0.0229783
R5518 VGND.n2067 VGND 0.0229783
R5519 VGND VGND.n2066 0.0229783
R5520 VGND.n2065 VGND 0.0229783
R5521 VGND.n2064 VGND 0.0229783
R5522 VGND.n2063 VGND 0.0229783
R5523 VGND.n2062 VGND 0.0229783
R5524 VGND.n2061 VGND 0.0229783
R5525 VGND.n2059 VGND 0.0229783
R5526 VGND VGND.n2058 0.0229783
R5527 VGND.n2056 VGND 0.0229783
R5528 VGND VGND.n2055 0.0229783
R5529 VGND.n2053 VGND 0.0229783
R5530 VGND VGND.n2052 0.0229783
R5531 VGND.n2050 VGND 0.0229783
R5532 VGND VGND.n2049 0.0229783
R5533 VGND.n2047 VGND 0.0229783
R5534 VGND.n2046 VGND 0.0229783
R5535 VGND.n2045 VGND 0.0229783
R5536 VGND.n2044 VGND 0.0229783
R5537 VGND VGND.n2040 0.0229783
R5538 VGND.n2039 VGND 0.0229783
R5539 VGND VGND.n1991 0.0229783
R5540 VGND VGND.n1993 0.0229783
R5541 VGND.n1995 VGND 0.0229783
R5542 VGND VGND.n1997 0.0229783
R5543 VGND VGND.n1999 0.0229783
R5544 VGND VGND.n2001 0.0229783
R5545 VGND VGND.n2003 0.0229783
R5546 VGND VGND.n2005 0.0229783
R5547 VGND.n2007 VGND 0.0229783
R5548 VGND VGND.n2012 0.0229783
R5549 VGND.n2014 VGND 0.0229783
R5550 VGND VGND.n2019 0.0229783
R5551 VGND VGND.n2021 0.0229783
R5552 VGND VGND.n2023 0.0229783
R5553 VGND.n2026 VGND 0.0229783
R5554 VGND.n2025 VGND 0.0229783
R5555 VGND VGND.n1126 0.0229783
R5556 VGND VGND.n1128 0.0229783
R5557 VGND VGND.n1130 0.0229783
R5558 VGND VGND.n1132 0.0229783
R5559 VGND.n1134 VGND 0.0229783
R5560 VGND VGND.n1136 0.0229783
R5561 VGND VGND.n1141 0.0229783
R5562 VGND VGND.n1143 0.0229783
R5563 VGND.n1144 VGND 0.0229783
R5564 VGND VGND.n1149 0.0229783
R5565 VGND VGND.n1104 0.0229783
R5566 VGND VGND.n1106 0.0229783
R5567 VGND VGND.n1108 0.0229783
R5568 VGND VGND.n1110 0.0229783
R5569 VGND VGND.n1112 0.0229783
R5570 VGND VGND.n1114 0.0229783
R5571 VGND VGND.n1116 0.0229783
R5572 VGND.n1120 VGND 0.0229783
R5573 VGND.n1923 VGND 0.0229783
R5574 VGND.n2762 VGND 0.0229783
R5575 VGND.n2761 VGND 0.0229783
R5576 VGND VGND.n2760 0.0229783
R5577 VGND.n2759 VGND 0.0229783
R5578 VGND.n2758 VGND 0.0229783
R5579 VGND.n2757 VGND 0.0229783
R5580 VGND.n2756 VGND 0.0229783
R5581 VGND.n2755 VGND 0.0229783
R5582 VGND.n2753 VGND 0.0229783
R5583 VGND VGND.n2752 0.0229783
R5584 VGND.n2750 VGND 0.0229783
R5585 VGND VGND.n2749 0.0229783
R5586 VGND.n2747 VGND 0.0229783
R5587 VGND VGND.n2746 0.0229783
R5588 VGND.n2744 VGND 0.0229783
R5589 VGND VGND.n2743 0.0229783
R5590 VGND.n2741 VGND 0.0229783
R5591 VGND.n2740 VGND 0.0229783
R5592 VGND.n2739 VGND 0.0229783
R5593 VGND.n2738 VGND 0.0229783
R5594 VGND VGND.n2734 0.0229783
R5595 VGND.n2733 VGND 0.0229783
R5596 VGND VGND.n741 0.0229783
R5597 VGND VGND.n743 0.0229783
R5598 VGND VGND.n745 0.0229783
R5599 VGND VGND.n747 0.0229783
R5600 VGND VGND.n749 0.0229783
R5601 VGND VGND.n751 0.0229783
R5602 VGND VGND.n753 0.0229783
R5603 VGND.n754 VGND 0.0229783
R5604 VGND VGND.n2378 0.0229783
R5605 VGND VGND.n792 0.0229783
R5606 VGND VGND.n794 0.0229783
R5607 VGND VGND.n796 0.0229783
R5608 VGND VGND.n798 0.0229783
R5609 VGND VGND.n800 0.0229783
R5610 VGND VGND.n802 0.0229783
R5611 VGND VGND.n804 0.0229783
R5612 VGND.n806 VGND 0.0229783
R5613 VGND.n2286 VGND 0.0229783
R5614 VGND VGND.n812 0.0229783
R5615 VGND VGND.n814 0.0229783
R5616 VGND VGND.n816 0.0229783
R5617 VGND VGND.n818 0.0229783
R5618 VGND VGND.n820 0.0229783
R5619 VGND VGND.n822 0.0229783
R5620 VGND VGND.n824 0.0229783
R5621 VGND.n825 VGND 0.0229783
R5622 VGND VGND.n835 0.0229783
R5623 VGND.n2273 VGND 0.0229783
R5624 VGND.n2272 VGND 0.0229783
R5625 VGND VGND.n2271 0.0229783
R5626 VGND.n2270 VGND 0.0229783
R5627 VGND.n2269 VGND 0.0229783
R5628 VGND.n2268 VGND 0.0229783
R5629 VGND.n2267 VGND 0.0229783
R5630 VGND.n2266 VGND 0.0229783
R5631 VGND.n2264 VGND 0.0229783
R5632 VGND VGND.n2263 0.0229783
R5633 VGND.n2261 VGND 0.0229783
R5634 VGND VGND.n2260 0.0229783
R5635 VGND.n2258 VGND 0.0229783
R5636 VGND VGND.n2257 0.0229783
R5637 VGND.n2255 VGND 0.0229783
R5638 VGND VGND.n2254 0.0229783
R5639 VGND.n2252 VGND 0.0229783
R5640 VGND.n2251 VGND 0.0229783
R5641 VGND.n2250 VGND 0.0229783
R5642 VGND.n2249 VGND 0.0229783
R5643 VGND VGND.n2245 0.0229783
R5644 VGND.n2244 VGND 0.0229783
R5645 VGND VGND.n2537 0.0229783
R5646 VGND VGND.n2539 0.0229783
R5647 VGND.n2541 VGND 0.0229783
R5648 VGND VGND.n2543 0.0229783
R5649 VGND VGND.n2545 0.0229783
R5650 VGND VGND.n2547 0.0229783
R5651 VGND VGND.n2549 0.0229783
R5652 VGND VGND.n2551 0.0229783
R5653 VGND VGND.n2556 0.0229783
R5654 VGND.n2558 VGND 0.0229783
R5655 VGND VGND.n2563 0.0229783
R5656 VGND.n2565 VGND 0.0229783
R5657 VGND VGND.n2570 0.0229783
R5658 VGND.n2572 VGND 0.0229783
R5659 VGND VGND.n2577 0.0229783
R5660 VGND.n2579 VGND 0.0229783
R5661 VGND VGND.n2584 0.0229783
R5662 VGND VGND.n2586 0.0229783
R5663 VGND VGND.n2588 0.0229783
R5664 VGND VGND.n2590 0.0229783
R5665 VGND.n2599 VGND 0.0229783
R5666 VGND.n2598 VGND 0.0229783
R5667 VGND.n659 VGND 0.0229783
R5668 VGND.n658 VGND 0.0229783
R5669 VGND VGND.n657 0.0229783
R5670 VGND.n656 VGND 0.0229783
R5671 VGND.n655 VGND 0.0229783
R5672 VGND.n654 VGND 0.0229783
R5673 VGND.n652 VGND 0.0229783
R5674 VGND VGND.n651 0.0229783
R5675 VGND.n650 VGND 0.0229783
R5676 VGND.n2275 VGND.n2073 0.0221569
R5677 VGND.n2526 VGND.n2525 0.0215388
R5678 VGND.n1703 VGND.n1542 0.017549
R5679 VGND.n2380 VGND.n738 0.0142311
R5680 VGND.n2380 VGND.n2379 0.0142311
R5681 VGND.n2765 VGND.n2764 0.0129412
R5682 VGND.n2765 VGND.n10 0.0120196
R5683 VGND.n1917 VGND.n1156 0.00816304
R5684 VGND.n1700 VGND.n1542 0.00741176
R5685 VGND.n2071 VGND.n840 0.00305435
R5686 VGND.n1438 VGND.n1437 0.00280392
R5687 VGND.n1914 VGND.n1913 0.00280392
R5688 VGND.n2279 VGND.n2073 0.00280392
R5689 VGND.n2767 VGND.n2766 0.000653482
R5690 VGND.n1916 VGND.n1915 0.000531323
R5691 VGND.n2072 VGND.n9 0.000531323
R5692 VGND.n2766 VGND.n9 0.000531323
R5693 VGND.n2072 VGND.n839 0.000525058
R5694 VGND.n1915 VGND.n839 0.000506265
R5695 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t8 568.956
R5696 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t9 568.956
R5697 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n3 292.5
R5698 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n9 292.5
R5699 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n12 197.272
R5700 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n2 112.829
R5701 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n6 112.829
R5702 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n4 111.059
R5703 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t1 63.8431
R5704 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t2 63.8431
R5705 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t3 63.8431
R5706 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t0 63.8431
R5707 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n7 59.1064
R5708 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n5 53.4593
R5709 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n8 51.9534
R5710 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n1 44.4312
R5711 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t6 38.8894
R5712 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t7 38.8894
R5713 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t5 38.8894
R5714 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.t4 38.8894
R5715 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 20.3299
R5716 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 20.3299
R5717 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n11 20.3299
R5718 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 20.3299
R5719 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n10 20.3299
R5720 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 17.6946
R5721 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 17.6946
R5722 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 12.325
R5723 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 12.323
R5724 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 10.3476
R5725 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n0 8.26099
R5726 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.168144
R5727 VPWR.n1174 VPWR.n1068 3277.03
R5728 VPWR.n1174 VPWR.n1173 2602.71
R5729 VPWR VPWR.n1172 667.92
R5730 VPWR.n1512 VPWR.t127 574.351
R5731 VPWR.n1511 VPWR.t205 574.351
R5732 VPWR.n1117 VPWR.t168 574.351
R5733 VPWR.n1017 VPWR.t199 572.875
R5734 VPWR.n2072 VPWR.t29 568.956
R5735 VPWR.n2137 VPWR.t195 568.956
R5736 VPWR.n2082 VPWR.t59 568.956
R5737 VPWR.n2203 VPWR.t105 568.956
R5738 VPWR.n2148 VPWR.t74 568.956
R5739 VPWR.n2269 VPWR.t152 568.956
R5740 VPWR.n2214 VPWR.t144 568.956
R5741 VPWR.n1435 VPWR.t133 568.956
R5742 VPWR.n1314 VPWR.t82 568.956
R5743 VPWR.n1277 VPWR.t67 568.956
R5744 VPWR.n1248 VPWR.t124 568.956
R5745 VPWR.n1724 VPWR.t97 568.956
R5746 VPWR.n1612 VPWR.t185 568.956
R5747 VPWR.n1528 VPWR.t78 568.956
R5748 VPWR.n1523 VPWR.t208 568.956
R5749 VPWR.n1524 VPWR.t160 568.956
R5750 VPWR.n1525 VPWR.t109 568.956
R5751 VPWR.n1526 VPWR.t63 568.956
R5752 VPWR.n1527 VPWR.t51 568.956
R5753 VPWR.n1586 VPWR.t156 568.956
R5754 VPWR.n1581 VPWR.t40 568.956
R5755 VPWR.n1582 VPWR.t116 568.956
R5756 VPWR.n1583 VPWR.t174 568.956
R5757 VPWR.n1584 VPWR.t89 568.956
R5758 VPWR.n1585 VPWR.t148 568.956
R5759 VPWR.n952 VPWR.t202 568.956
R5760 VPWR.n931 VPWR.t33 568.956
R5761 VPWR.n780 VPWR.t189 568.956
R5762 VPWR.n954 VPWR.t93 568.956
R5763 VPWR.n1900 VPWR.t130 568.956
R5764 VPWR.n1779 VPWR.t113 568.956
R5765 VPWR.n1742 VPWR.t70 568.956
R5766 VPWR.n327 VPWR.t171 568.956
R5767 VPWR.n1940 VPWR.t85 568.956
R5768 VPWR.n622 VPWR.t101 568.956
R5769 VPWR.n601 VPWR.t182 568.956
R5770 VPWR.n450 VPWR.t192 568.956
R5771 VPWR.n624 VPWR.t48 568.956
R5772 VPWR.n1103 VPWR.t136 568.956
R5773 VPWR.n1166 VPWR.t140 568.956
R5774 VPWR.n1130 VPWR.t120 568.956
R5775 VPWR.n1007 VPWR.t44 568.956
R5776 VPWR.n1028 VPWR.t36 568.956
R5777 VPWR.n1064 VPWR.t178 568.956
R5778 VPWR.n2335 VPWR.t164 568.956
R5779 VPWR.n2280 VPWR.t55 568.956
R5780 VPWR.n1172 VPWR.n1068 425.372
R5781 VPWR.n1980 VPWR.t290 361.738
R5782 VPWR.n1981 VPWR.t332 361.738
R5783 VPWR.n1983 VPWR.t230 361.738
R5784 VPWR.n1985 VPWR.t14 361.738
R5785 VPWR.n1987 VPWR.t595 361.738
R5786 VPWR.n1989 VPWR.t311 361.738
R5787 VPWR.n1991 VPWR.t16 361.738
R5788 VPWR.n1996 VPWR.t227 361.738
R5789 VPWR.n1998 VPWR.t20 361.738
R5790 VPWR.n156 VPWR.t279 361.738
R5791 VPWR.n157 VPWR.t340 361.738
R5792 VPWR.n159 VPWR.t260 361.738
R5793 VPWR.n161 VPWR.t265 361.738
R5794 VPWR.n163 VPWR.t259 361.738
R5795 VPWR.n165 VPWR.t513 361.738
R5796 VPWR.n167 VPWR.t435 361.738
R5797 VPWR.n169 VPWR.t502 361.738
R5798 VPWR.n116 VPWR.t283 361.738
R5799 VPWR.n117 VPWR.t438 361.738
R5800 VPWR.n119 VPWR.t238 361.738
R5801 VPWR.n121 VPWR.t243 361.738
R5802 VPWR.n123 VPWR.t237 361.738
R5803 VPWR.n125 VPWR.t579 361.738
R5804 VPWR.n127 VPWR.t457 361.738
R5805 VPWR.n129 VPWR.t503 361.738
R5806 VPWR.n76 VPWR.t271 361.738
R5807 VPWR.n77 VPWR.t356 361.738
R5808 VPWR.n79 VPWR.t239 361.738
R5809 VPWR.n81 VPWR.t256 361.738
R5810 VPWR.n83 VPWR.t240 361.738
R5811 VPWR.n85 VPWR.t548 361.738
R5812 VPWR.n87 VPWR.t466 361.738
R5813 VPWR.n89 VPWR.t498 361.738
R5814 VPWR.n1212 VPWR.t333 361.738
R5815 VPWR.n1214 VPWR.t212 361.738
R5816 VPWR.n1216 VPWR.t8 361.738
R5817 VPWR.n1218 VPWR.t7 361.738
R5818 VPWR.n1220 VPWR.t268 361.738
R5819 VPWR.n1222 VPWR.t269 361.738
R5820 VPWR.n1224 VPWR.t232 361.738
R5821 VPWR.n1229 VPWR.t526 361.738
R5822 VPWR.n1231 VPWR.t524 361.738
R5823 VPWR.n1233 VPWR.t231 361.738
R5824 VPWR.n1235 VPWR.t325 361.738
R5825 VPWR.n1237 VPWR.t522 361.738
R5826 VPWR.n1513 VPWR.t3 361.738
R5827 VPWR.n1515 VPWR.t597 361.738
R5828 VPWR.n1517 VPWR.t5 361.738
R5829 VPWR.n1519 VPWR.t281 361.738
R5830 VPWR.n1521 VPWR.t373 361.738
R5831 VPWR.n1545 VPWR.t442 361.738
R5832 VPWR.n1556 VPWR.t446 361.738
R5833 VPWR.n1561 VPWR.t444 361.738
R5834 VPWR.n1563 VPWR.t387 361.738
R5835 VPWR.n1568 VPWR.t391 361.738
R5836 VPWR.n1570 VPWR.t383 361.738
R5837 VPWR.n745 VPWR.t216 361.738
R5838 VPWR.n747 VPWR.t303 361.738
R5839 VPWR.n749 VPWR.t270 361.738
R5840 VPWR.n751 VPWR.t274 361.738
R5841 VPWR.n753 VPWR.t326 361.738
R5842 VPWR.n755 VPWR.t327 361.738
R5843 VPWR.n757 VPWR.t249 361.738
R5844 VPWR.n762 VPWR.t533 361.738
R5845 VPWR.n764 VPWR.t534 361.738
R5846 VPWR.n766 VPWR.t248 361.738
R5847 VPWR.n768 VPWR.t261 361.738
R5848 VPWR.n770 VPWR.t527 361.738
R5849 VPWR.n291 VPWR.t317 361.738
R5850 VPWR.n293 VPWR.t250 361.738
R5851 VPWR.n295 VPWR.t225 361.738
R5852 VPWR.n297 VPWR.t224 361.738
R5853 VPWR.n299 VPWR.t306 361.738
R5854 VPWR.n301 VPWR.t307 361.738
R5855 VPWR.n303 VPWR.t304 361.738
R5856 VPWR.n308 VPWR.t519 361.738
R5857 VPWR.n310 VPWR.t530 361.738
R5858 VPWR.n312 VPWR.t305 361.738
R5859 VPWR.n314 VPWR.t28 361.738
R5860 VPWR.n316 VPWR.t538 361.738
R5861 VPWR.n415 VPWR.t315 361.738
R5862 VPWR.n417 VPWR.t314 361.738
R5863 VPWR.n419 VPWR.t12 361.738
R5864 VPWR.n421 VPWR.t293 361.738
R5865 VPWR.n423 VPWR.t11 361.738
R5866 VPWR.n425 VPWR.t10 361.738
R5867 VPWR.n427 VPWR.t244 361.738
R5868 VPWR.n432 VPWR.t529 361.738
R5869 VPWR.n434 VPWR.t520 361.738
R5870 VPWR.n436 VPWR.t245 361.738
R5871 VPWR.n438 VPWR.t273 361.738
R5872 VPWR.n440 VPWR.t541 361.738
R5873 VPWR.n1109 VPWR.t247 361.738
R5874 VPWR.n1115 VPWR.t302 361.738
R5875 VPWR.n1116 VPWR.t324 361.738
R5876 VPWR.n1120 VPWR.t428 361.738
R5877 VPWR.n29 VPWR.t251 361.738
R5878 VPWR.n30 VPWR.t367 361.738
R5879 VPWR.n32 VPWR.t286 361.738
R5880 VPWR.n34 VPWR.t337 361.738
R5881 VPWR.n36 VPWR.t287 361.738
R5882 VPWR.n38 VPWR.t575 361.738
R5883 VPWR.n40 VPWR.t453 361.738
R5884 VPWR.n42 VPWR.t499 361.738
R5885 VPWR.n370 VPWR.t459 361.738
R5886 VPWR.n369 VPWR.t461 361.738
R5887 VPWR.n375 VPWR.t464 361.738
R5888 VPWR.n374 VPWR.t465 361.738
R5889 VPWR.n380 VPWR.t433 361.738
R5890 VPWR.n379 VPWR.t434 361.738
R5891 VPWR.n385 VPWR.t401 361.738
R5892 VPWR.n384 VPWR.t399 361.738
R5893 VPWR.n4 VPWR.t586 361.738
R5894 VPWR.n3 VPWR.t588 361.738
R5895 VPWR.n9 VPWR.t543 361.738
R5896 VPWR.n8 VPWR.t544 361.738
R5897 VPWR.n14 VPWR.t577 361.738
R5898 VPWR.n13 VPWR.t578 361.738
R5899 VPWR.n19 VPWR.t481 361.738
R5900 VPWR.n18 VPWR.t482 361.738
R5901 VPWR.n700 VPWR.t601 361.738
R5902 VPWR.n699 VPWR.t599 361.738
R5903 VPWR.n705 VPWR.t581 361.738
R5904 VPWR.n704 VPWR.t582 361.738
R5905 VPWR.n710 VPWR.t406 361.738
R5906 VPWR.n709 VPWR.t403 361.738
R5907 VPWR.n715 VPWR.t377 361.738
R5908 VPWR.n714 VPWR.t375 361.738
R5909 VPWR.n231 VPWR.t470 361.738
R5910 VPWR.n230 VPWR.t468 361.738
R5911 VPWR.n236 VPWR.t412 361.738
R5912 VPWR.n235 VPWR.t409 361.738
R5913 VPWR.n241 VPWR.t492 361.738
R5914 VPWR.n240 VPWR.t489 361.738
R5915 VPWR.n246 VPWR.t222 361.738
R5916 VPWR.n245 VPWR.t220 361.738
R5917 VPWR.n1251 VPWR.t22 360.264
R5918 VPWR.n1250 VPWR.t23 360.264
R5919 VPWR.n1256 VPWR.t487 360.264
R5920 VPWR.n1255 VPWR.t486 360.264
R5921 VPWR.n1261 VPWR.t566 360.264
R5922 VPWR.n1260 VPWR.t568 360.264
R5923 VPWR.n1266 VPWR.t590 360.264
R5924 VPWR.n1265 VPWR.t589 360.264
R5925 VPWR.n657 VPWR.t361 360.264
R5926 VPWR.n656 VPWR.t346 360.264
R5927 VPWR.n662 VPWR.t349 360.264
R5928 VPWR.n661 VPWR.t348 360.264
R5929 VPWR.n667 VPWR.t507 360.264
R5930 VPWR.n666 VPWR.t508 360.264
R5931 VPWR.n672 VPWR.t510 360.264
R5932 VPWR.n671 VPWR.t425 360.264
R5933 VPWR.n199 VPWR.t456 360.264
R5934 VPWR.n198 VPWR.t478 360.264
R5935 VPWR.n204 VPWR.t357 360.264
R5936 VPWR.n203 VPWR.t359 360.264
R5937 VPWR.n209 VPWR.t517 360.264
R5938 VPWR.n208 VPWR.t518 360.264
R5939 VPWR.n214 VPWR.t495 360.264
R5940 VPWR.n213 VPWR.t493 360.264
R5941 VPWR.n346 VPWR.t422 360.264
R5942 VPWR.n345 VPWR.t423 360.264
R5943 VPWR.n351 VPWR.t416 360.264
R5944 VPWR.n350 VPWR.t415 360.264
R5945 VPWR.n356 VPWR.t571 360.264
R5946 VPWR.n355 VPWR.t572 360.264
R5947 VPWR.n361 VPWR.t396 360.264
R5948 VPWR.n360 VPWR.t397 360.264
R5949 VPWR.n2080 VPWR.t62 360.264
R5950 VPWR.n177 VPWR.t217 360.264
R5951 VPWR.n178 VPWR.t419 360.264
R5952 VPWR.n180 VPWR.t275 360.264
R5953 VPWR.n182 VPWR.t272 360.264
R5954 VPWR.n184 VPWR.t276 360.264
R5955 VPWR.n186 VPWR.t352 360.264
R5956 VPWR.n188 VPWR.t355 360.264
R5957 VPWR.n190 VPWR.t477 360.264
R5958 VPWR.n192 VPWR.t61 360.264
R5959 VPWR.n2146 VPWR.t77 360.264
R5960 VPWR.n137 VPWR.t291 360.264
R5961 VPWR.n138 VPWR.t338 360.264
R5962 VPWR.n140 VPWR.t215 360.264
R5963 VPWR.n142 VPWR.t213 360.264
R5964 VPWR.n144 VPWR.t214 360.264
R5965 VPWR.n146 VPWR.t223 360.264
R5966 VPWR.n148 VPWR.t354 360.264
R5967 VPWR.n150 VPWR.t476 360.264
R5968 VPWR.n152 VPWR.t76 360.264
R5969 VPWR.n2212 VPWR.t147 360.264
R5970 VPWR.n97 VPWR.t295 360.264
R5971 VPWR.n98 VPWR.t339 360.264
R5972 VPWR.n100 VPWR.t253 360.264
R5973 VPWR.n102 VPWR.t262 360.264
R5974 VPWR.n104 VPWR.t252 360.264
R5975 VPWR.n106 VPWR.t549 360.264
R5976 VPWR.n108 VPWR.t424 360.264
R5977 VPWR.n110 VPWR.t504 360.264
R5978 VPWR.n112 VPWR.t146 360.264
R5979 VPWR.n1312 VPWR.t84 360.264
R5980 VPWR.n1280 VPWR.t69 360.264
R5981 VPWR.n1278 VPWR.t68 360.264
R5982 VPWR.n1282 VPWR.t264 360.264
R5983 VPWR.n1284 VPWR.t263 360.264
R5984 VPWR.n1286 VPWR.t321 360.264
R5985 VPWR.n1288 VPWR.t300 360.264
R5986 VPWR.n1290 VPWR.t319 360.264
R5987 VPWR.n1292 VPWR.t320 360.264
R5988 VPWR.n1294 VPWR.t392 360.264
R5989 VPWR.n1299 VPWR.t537 360.264
R5990 VPWR.n1301 VPWR.t531 360.264
R5991 VPWR.n1303 VPWR.t393 360.264
R5992 VPWR.n1305 VPWR.t233 360.264
R5993 VPWR.n1307 VPWR.t542 360.264
R5994 VPWR.n1309 VPWR.t83 360.264
R5995 VPWR.n949 VPWR.t204 360.264
R5996 VPWR.n741 VPWR.t35 360.264
R5997 VPWR.n950 VPWR.t203 360.264
R5998 VPWR.n726 VPWR.t266 360.264
R5999 VPWR.n727 VPWR.t328 360.264
R6000 VPWR.n728 VPWR.t322 360.264
R6001 VPWR.n729 VPWR.t267 360.264
R6002 VPWR.n730 VPWR.t277 360.264
R6003 VPWR.n731 VPWR.t278 360.264
R6004 VPWR.n732 VPWR.t408 360.264
R6005 VPWR.n735 VPWR.t539 360.264
R6006 VPWR.n736 VPWR.t528 360.264
R6007 VPWR.n737 VPWR.t407 360.264
R6008 VPWR.n738 VPWR.t312 360.264
R6009 VPWR.n739 VPWR.t521 360.264
R6010 VPWR.n933 VPWR.t34 360.264
R6011 VPWR.n1777 VPWR.t115 360.264
R6012 VPWR.n1745 VPWR.t73 360.264
R6013 VPWR.n1743 VPWR.t72 360.264
R6014 VPWR.n1747 VPWR.t284 360.264
R6015 VPWR.n1749 VPWR.t294 360.264
R6016 VPWR.n1751 VPWR.t292 360.264
R6017 VPWR.n1753 VPWR.t285 360.264
R6018 VPWR.n1755 VPWR.t299 360.264
R6019 VPWR.n1757 VPWR.t298 360.264
R6020 VPWR.n1759 VPWR.t342 360.264
R6021 VPWR.n1764 VPWR.t540 360.264
R6022 VPWR.n1766 VPWR.t523 360.264
R6023 VPWR.n1768 VPWR.t341 360.264
R6024 VPWR.n1770 VPWR.t288 360.264
R6025 VPWR.n1772 VPWR.t532 360.264
R6026 VPWR.n1774 VPWR.t114 360.264
R6027 VPWR.n619 VPWR.t104 360.264
R6028 VPWR.n411 VPWR.t184 360.264
R6029 VPWR.n620 VPWR.t103 360.264
R6030 VPWR.n396 VPWR.t313 360.264
R6031 VPWR.n397 VPWR.t318 360.264
R6032 VPWR.n398 VPWR.t334 360.264
R6033 VPWR.n399 VPWR.t316 360.264
R6034 VPWR.n400 VPWR.t258 360.264
R6035 VPWR.n401 VPWR.t257 360.264
R6036 VPWR.n402 VPWR.t437 360.264
R6037 VPWR.n405 VPWR.t535 360.264
R6038 VPWR.n406 VPWR.t536 360.264
R6039 VPWR.n407 VPWR.t436 360.264
R6040 VPWR.n408 VPWR.t308 360.264
R6041 VPWR.n409 VPWR.t525 360.264
R6042 VPWR.n603 VPWR.t183 360.264
R6043 VPWR.n1009 VPWR.t47 360.264
R6044 VPWR.n1026 VPWR.t39 360.264
R6045 VPWR.n1066 VPWR.t181 360.264
R6046 VPWR.n998 VPWR.t46 360.264
R6047 VPWR.n1011 VPWR.t336 360.264
R6048 VPWR.n1015 VPWR.t242 360.264
R6049 VPWR.n1016 VPWR.t255 360.264
R6050 VPWR.n1020 VPWR.t430 360.264
R6051 VPWR.n1013 VPWR.t38 360.264
R6052 VPWR.n984 VPWR.t180 360.264
R6053 VPWR.n2278 VPWR.t58 360.264
R6054 VPWR.n50 VPWR.t309 360.264
R6055 VPWR.n51 VPWR.t343 360.264
R6056 VPWR.n53 VPWR.t297 360.264
R6057 VPWR.n55 VPWR.t282 360.264
R6058 VPWR.n57 VPWR.t296 360.264
R6059 VPWR.n59 VPWR.t414 360.264
R6060 VPWR.n61 VPWR.t379 360.264
R6061 VPWR.n63 VPWR.t505 360.264
R6062 VPWR.n65 VPWR.t57 360.264
R6063 VPWR.n2074 VPWR.t32 356.344
R6064 VPWR.n2002 VPWR.t31 356.344
R6065 VPWR.n2139 VPWR.t198 356.344
R6066 VPWR.n173 VPWR.t197 356.344
R6067 VPWR.n2205 VPWR.t108 356.344
R6068 VPWR.n133 VPWR.t107 356.344
R6069 VPWR.n2271 VPWR.t155 356.344
R6070 VPWR.n93 VPWR.t154 356.344
R6071 VPWR.n1436 VPWR.t135 356.344
R6072 VPWR.n1441 VPWR.t134 356.344
R6073 VPWR.n1211 VPWR.t126 356.344
R6074 VPWR.n1239 VPWR.t125 356.344
R6075 VPWR.n1725 VPWR.t100 356.344
R6076 VPWR.n1730 VPWR.t99 356.344
R6077 VPWR.n1510 VPWR.t188 356.344
R6078 VPWR.n1603 VPWR.t187 356.344
R6079 VPWR.n1530 VPWR.t80 356.344
R6080 VPWR.n1588 VPWR.t158 356.344
R6081 VPWR.n743 VPWR.t191 356.344
R6082 VPWR.n955 VPWR.t96 356.344
R6083 VPWR.n960 VPWR.t95 356.344
R6084 VPWR.n772 VPWR.t190 356.344
R6085 VPWR.n1901 VPWR.t132 356.344
R6086 VPWR.n1906 VPWR.t131 356.344
R6087 VPWR.n290 VPWR.t173 356.344
R6088 VPWR.n318 VPWR.t172 356.344
R6089 VPWR.n1943 VPWR.t88 356.344
R6090 VPWR.n1916 VPWR.t87 356.344
R6091 VPWR.n1948 VPWR.t330 356.344
R6092 VPWR.n1953 VPWR.t235 356.344
R6093 VPWR.n1958 VPWR.t501 356.344
R6094 VPWR.n413 VPWR.t194 356.344
R6095 VPWR.n625 VPWR.t50 356.344
R6096 VPWR.n630 VPWR.t49 356.344
R6097 VPWR.n442 VPWR.t193 356.344
R6098 VPWR.n1105 VPWR.t139 356.344
R6099 VPWR.n1093 VPWR.t138 356.344
R6100 VPWR.n1168 VPWR.t143 356.344
R6101 VPWR.n1071 VPWR.t142 356.344
R6102 VPWR.n1089 VPWR.t123 356.344
R6103 VPWR.n1111 VPWR.t122 356.344
R6104 VPWR.n2337 VPWR.t167 356.344
R6105 VPWR.n46 VPWR.t166 356.344
R6106 VPWR.n1994 VPWR.n1993 297.897
R6107 VPWR.n1227 VPWR.n1226 297.897
R6108 VPWR.n1548 VPWR.n1547 297.897
R6109 VPWR.n1551 VPWR.n1550 297.897
R6110 VPWR.n1554 VPWR.n1553 297.897
R6111 VPWR.n1559 VPWR.n1558 297.897
R6112 VPWR.n1566 VPWR.n1565 297.897
R6113 VPWR.n1573 VPWR.n1572 297.897
R6114 VPWR.n1576 VPWR.n1575 297.897
R6115 VPWR.n1579 VPWR.n1578 297.897
R6116 VPWR.n760 VPWR.n759 297.897
R6117 VPWR.n306 VPWR.n305 297.897
R6118 VPWR.n430 VPWR.n429 297.897
R6119 VPWR.n1119 VPWR.n1118 297.897
R6120 VPWR.n372 VPWR.n371 297.896
R6121 VPWR.n377 VPWR.n376 297.896
R6122 VPWR.n382 VPWR.n381 297.896
R6123 VPWR.n387 VPWR.n386 297.896
R6124 VPWR.n6 VPWR.n5 297.896
R6125 VPWR.n11 VPWR.n10 297.896
R6126 VPWR.n16 VPWR.n15 297.896
R6127 VPWR.n21 VPWR.n20 297.896
R6128 VPWR.n702 VPWR.n701 297.896
R6129 VPWR.n707 VPWR.n706 297.896
R6130 VPWR.n712 VPWR.n711 297.896
R6131 VPWR.n717 VPWR.n716 297.896
R6132 VPWR.n233 VPWR.n232 297.896
R6133 VPWR.n238 VPWR.n237 297.896
R6134 VPWR.n243 VPWR.n242 297.896
R6135 VPWR.n248 VPWR.n247 297.896
R6136 VPWR.n1253 VPWR.n1252 296.421
R6137 VPWR.n1258 VPWR.n1257 296.421
R6138 VPWR.n1263 VPWR.n1262 296.421
R6139 VPWR.n1268 VPWR.n1267 296.421
R6140 VPWR.n659 VPWR.n658 296.421
R6141 VPWR.n664 VPWR.n663 296.421
R6142 VPWR.n669 VPWR.n668 296.421
R6143 VPWR.n674 VPWR.n673 296.421
R6144 VPWR.n201 VPWR.n200 296.421
R6145 VPWR.n206 VPWR.n205 296.421
R6146 VPWR.n211 VPWR.n210 296.421
R6147 VPWR.n216 VPWR.n215 296.421
R6148 VPWR.n348 VPWR.n347 296.421
R6149 VPWR.n353 VPWR.n352 296.421
R6150 VPWR.n358 VPWR.n357 296.421
R6151 VPWR.n363 VPWR.n362 296.421
R6152 VPWR.n1297 VPWR.n1296 296.421
R6153 VPWR.n734 VPWR.n733 296.421
R6154 VPWR.n1762 VPWR.n1761 296.421
R6155 VPWR.n404 VPWR.n403 296.421
R6156 VPWR.n1019 VPWR.n1018 296.421
R6157 VPWR.n1532 VPWR.n1531 292.5
R6158 VPWR.n1534 VPWR.n1533 292.5
R6159 VPWR.n1536 VPWR.n1535 292.5
R6160 VPWR.n1538 VPWR.n1537 292.5
R6161 VPWR.n1540 VPWR.n1539 292.5
R6162 VPWR.n1542 VPWR.n1541 292.5
R6163 VPWR.n1590 VPWR.n1589 292.5
R6164 VPWR.n1592 VPWR.n1591 292.5
R6165 VPWR.n1594 VPWR.n1593 292.5
R6166 VPWR.n1596 VPWR.n1595 292.5
R6167 VPWR.n1598 VPWR.n1597 292.5
R6168 VPWR.n1600 VPWR.n1599 292.5
R6169 VPWR.t289 VPWR.n2021 243.056
R6170 VPWR.n2070 VPWR.t30 243.056
R6171 VPWR.t98 VPWR.n1454 243.056
R6172 VPWR.t186 VPWR.n1614 243.056
R6173 VPWR.t86 VPWR.n1919 243.056
R6174 VPWR.t500 VPWR.n1926 243.056
R6175 VPWR.t137 VPWR.n1095 243.056
R6176 VPWR.n1164 VPWR.t141 243.056
R6177 VPWR.t45 VPWR.n999 243.056
R6178 VPWR.n1062 VPWR.t179 243.056
R6179 VPWR.n2078 VPWR 228.48
R6180 VPWR.n1429 VPWR 226.279
R6181 VPWR VPWR.n929 226.279
R6182 VPWR.n1894 VPWR 226.279
R6183 VPWR VPWR.n599 226.279
R6184 VPWR.n2144 VPWR.n2143 225.024
R6185 VPWR.n2210 VPWR.n2209 225.024
R6186 VPWR.n2276 VPWR.n2275 225.024
R6187 VPWR.n2134 VPWR.t60 198.453
R6188 VPWR.n2134 VPWR.t196 198.453
R6189 VPWR.n2200 VPWR.t75 198.453
R6190 VPWR.n2200 VPWR.t106 198.453
R6191 VPWR.n2266 VPWR.t145 198.453
R6192 VPWR.n2266 VPWR.t153 198.453
R6193 VPWR.n2332 VPWR.t56 198.453
R6194 VPWR.n2332 VPWR.t165 198.453
R6195 VPWR.n2021 VPWR 192.822
R6196 VPWR.n2133 VPWR 192.822
R6197 VPWR.n2199 VPWR 192.822
R6198 VPWR.n2265 VPWR 192.822
R6199 VPWR.n2331 VPWR 192.822
R6200 VPWR.n1434 VPWR.n1178 190.215
R6201 VPWR.n1723 VPWR.n1454 190.215
R6202 VPWR.n953 VPWR.n725 190.215
R6203 VPWR.n1899 VPWR.n257 190.215
R6204 VPWR.n1939 VPWR.n1919 190.215
R6205 VPWR.n623 VPWR.n395 190.215
R6206 VPWR.n1102 VPWR.n1095 190.215
R6207 VPWR.n1006 VPWR.n999 190.215
R6208 VPWR VPWR.n2070 187.607
R6209 VPWR VPWR.n2135 187.607
R6210 VPWR VPWR.n2201 187.607
R6211 VPWR VPWR.n2267 187.607
R6212 VPWR.n1614 VPWR 187.607
R6213 VPWR.n1926 VPWR 187.607
R6214 VPWR VPWR.n1164 187.607
R6215 VPWR VPWR.n1062 187.607
R6216 VPWR VPWR.n2333 187.607
R6217 VPWR.n2020 VPWR.n2019 185
R6218 VPWR.n2022 VPWR.n2020 185
R6219 VPWR.n2025 VPWR.n2024 185
R6220 VPWR.n2024 VPWR.n2023 185
R6221 VPWR.n2026 VPWR.n2018 185
R6222 VPWR.n2018 VPWR.n2017 185
R6223 VPWR.n2029 VPWR.n2028 185
R6224 VPWR.n2030 VPWR.n2029 185
R6225 VPWR.n2027 VPWR.n2016 185
R6226 VPWR.n2031 VPWR.n2016 185
R6227 VPWR.n2035 VPWR.n2034 185
R6228 VPWR.n2034 VPWR.n2033 185
R6229 VPWR.n2036 VPWR.n2015 185
R6230 VPWR.n2032 VPWR.n2015 185
R6231 VPWR.n2039 VPWR.n2038 185
R6232 VPWR.n2040 VPWR.n2039 185
R6233 VPWR.n2037 VPWR.n2014 185
R6234 VPWR.n2041 VPWR.n2014 185
R6235 VPWR.n2045 VPWR.n2044 185
R6236 VPWR.n2044 VPWR.n2043 185
R6237 VPWR.n2046 VPWR.n2013 185
R6238 VPWR.n2042 VPWR.n2013 185
R6239 VPWR.n2048 VPWR.n2047 185
R6240 VPWR.n2049 VPWR.n2048 185
R6241 VPWR.n2012 VPWR.n2011 185
R6242 VPWR.n2050 VPWR.n2012 185
R6243 VPWR.n2054 VPWR.n2053 185
R6244 VPWR.n2053 VPWR.n2052 185
R6245 VPWR.n2055 VPWR.n2010 185
R6246 VPWR.n2051 VPWR.n2010 185
R6247 VPWR.n2058 VPWR.n2057 185
R6248 VPWR.n2059 VPWR.n2058 185
R6249 VPWR.n2056 VPWR.n2009 185
R6250 VPWR.n2060 VPWR.n2009 185
R6251 VPWR.n2064 VPWR.n2063 185
R6252 VPWR.n2063 VPWR.n2062 185
R6253 VPWR.n2065 VPWR.n2008 185
R6254 VPWR.n2061 VPWR.n2008 185
R6255 VPWR.n2067 VPWR.n2066 185
R6256 VPWR.n2068 VPWR.n2067 185
R6257 VPWR.n2007 VPWR.n2006 185
R6258 VPWR.n2069 VPWR.n2007 185
R6259 VPWR.n2134 VPWR.n2133 185
R6260 VPWR.n2132 VPWR.n2095 185
R6261 VPWR.n2131 VPWR.n2130 185
R6262 VPWR.n2129 VPWR.n2128 185
R6263 VPWR.n2127 VPWR.n2126 185
R6264 VPWR.n2125 VPWR.n2124 185
R6265 VPWR.n2123 VPWR.n2122 185
R6266 VPWR.n2121 VPWR.n2120 185
R6267 VPWR.n2119 VPWR.n2118 185
R6268 VPWR.n2117 VPWR.n2116 185
R6269 VPWR.n2115 VPWR.n2114 185
R6270 VPWR.n2113 VPWR.n2112 185
R6271 VPWR.n2111 VPWR.n2110 185
R6272 VPWR.n2109 VPWR.n2108 185
R6273 VPWR.n2107 VPWR.n2106 185
R6274 VPWR.n2105 VPWR.n2104 185
R6275 VPWR.n2103 VPWR.n2102 185
R6276 VPWR.n2101 VPWR.n2100 185
R6277 VPWR.n2099 VPWR.n2098 185
R6278 VPWR.n2097 VPWR.n2096 185
R6279 VPWR.n2084 VPWR.n2083 185
R6280 VPWR.n2135 VPWR.n2134 185
R6281 VPWR.n2200 VPWR.n2199 185
R6282 VPWR.n2198 VPWR.n2161 185
R6283 VPWR.n2197 VPWR.n2196 185
R6284 VPWR.n2195 VPWR.n2194 185
R6285 VPWR.n2193 VPWR.n2192 185
R6286 VPWR.n2191 VPWR.n2190 185
R6287 VPWR.n2189 VPWR.n2188 185
R6288 VPWR.n2187 VPWR.n2186 185
R6289 VPWR.n2185 VPWR.n2184 185
R6290 VPWR.n2183 VPWR.n2182 185
R6291 VPWR.n2181 VPWR.n2180 185
R6292 VPWR.n2179 VPWR.n2178 185
R6293 VPWR.n2177 VPWR.n2176 185
R6294 VPWR.n2175 VPWR.n2174 185
R6295 VPWR.n2173 VPWR.n2172 185
R6296 VPWR.n2171 VPWR.n2170 185
R6297 VPWR.n2169 VPWR.n2168 185
R6298 VPWR.n2167 VPWR.n2166 185
R6299 VPWR.n2165 VPWR.n2164 185
R6300 VPWR.n2163 VPWR.n2162 185
R6301 VPWR.n2150 VPWR.n2149 185
R6302 VPWR.n2201 VPWR.n2200 185
R6303 VPWR.n2266 VPWR.n2265 185
R6304 VPWR.n2264 VPWR.n2227 185
R6305 VPWR.n2263 VPWR.n2262 185
R6306 VPWR.n2261 VPWR.n2260 185
R6307 VPWR.n2259 VPWR.n2258 185
R6308 VPWR.n2257 VPWR.n2256 185
R6309 VPWR.n2255 VPWR.n2254 185
R6310 VPWR.n2253 VPWR.n2252 185
R6311 VPWR.n2251 VPWR.n2250 185
R6312 VPWR.n2249 VPWR.n2248 185
R6313 VPWR.n2247 VPWR.n2246 185
R6314 VPWR.n2245 VPWR.n2244 185
R6315 VPWR.n2243 VPWR.n2242 185
R6316 VPWR.n2241 VPWR.n2240 185
R6317 VPWR.n2239 VPWR.n2238 185
R6318 VPWR.n2237 VPWR.n2236 185
R6319 VPWR.n2235 VPWR.n2234 185
R6320 VPWR.n2233 VPWR.n2232 185
R6321 VPWR.n2231 VPWR.n2230 185
R6322 VPWR.n2229 VPWR.n2228 185
R6323 VPWR.n2216 VPWR.n2215 185
R6324 VPWR.n2267 VPWR.n2266 185
R6325 VPWR.n1430 VPWR.n1178 185
R6326 VPWR.n1433 VPWR.n1432 185
R6327 VPWR.n1180 VPWR.n1179 185
R6328 VPWR.n1316 VPWR.n1315 185
R6329 VPWR.n1318 VPWR.n1317 185
R6330 VPWR.n1320 VPWR.n1319 185
R6331 VPWR.n1322 VPWR.n1321 185
R6332 VPWR.n1324 VPWR.n1323 185
R6333 VPWR.n1326 VPWR.n1325 185
R6334 VPWR.n1328 VPWR.n1327 185
R6335 VPWR.n1330 VPWR.n1329 185
R6336 VPWR.n1332 VPWR.n1331 185
R6337 VPWR.n1334 VPWR.n1333 185
R6338 VPWR.n1336 VPWR.n1335 185
R6339 VPWR.n1338 VPWR.n1337 185
R6340 VPWR.n1340 VPWR.n1339 185
R6341 VPWR.n1342 VPWR.n1341 185
R6342 VPWR.n1344 VPWR.n1343 185
R6343 VPWR.n1346 VPWR.n1345 185
R6344 VPWR.n1348 VPWR.n1347 185
R6345 VPWR.n1350 VPWR.n1349 185
R6346 VPWR.n1352 VPWR.n1351 185
R6347 VPWR.n1354 VPWR.n1353 185
R6348 VPWR.n1356 VPWR.n1355 185
R6349 VPWR.n1358 VPWR.n1357 185
R6350 VPWR.n1360 VPWR.n1359 185
R6351 VPWR.n1362 VPWR.n1361 185
R6352 VPWR.n1364 VPWR.n1363 185
R6353 VPWR.n1366 VPWR.n1365 185
R6354 VPWR.n1368 VPWR.n1367 185
R6355 VPWR.n1370 VPWR.n1369 185
R6356 VPWR.n1372 VPWR.n1371 185
R6357 VPWR.n1374 VPWR.n1373 185
R6358 VPWR.n1376 VPWR.n1375 185
R6359 VPWR.n1378 VPWR.n1377 185
R6360 VPWR.n1380 VPWR.n1379 185
R6361 VPWR.n1382 VPWR.n1381 185
R6362 VPWR.n1384 VPWR.n1383 185
R6363 VPWR.n1386 VPWR.n1385 185
R6364 VPWR.n1388 VPWR.n1387 185
R6365 VPWR.n1390 VPWR.n1389 185
R6366 VPWR.n1392 VPWR.n1391 185
R6367 VPWR.n1394 VPWR.n1393 185
R6368 VPWR.n1396 VPWR.n1395 185
R6369 VPWR.n1398 VPWR.n1397 185
R6370 VPWR.n1400 VPWR.n1399 185
R6371 VPWR.n1402 VPWR.n1401 185
R6372 VPWR.n1404 VPWR.n1403 185
R6373 VPWR.n1406 VPWR.n1405 185
R6374 VPWR.n1408 VPWR.n1407 185
R6375 VPWR.n1410 VPWR.n1409 185
R6376 VPWR.n1412 VPWR.n1411 185
R6377 VPWR.n1414 VPWR.n1413 185
R6378 VPWR.n1416 VPWR.n1415 185
R6379 VPWR.n1418 VPWR.n1417 185
R6380 VPWR.n1420 VPWR.n1419 185
R6381 VPWR.n1422 VPWR.n1421 185
R6382 VPWR.n1424 VPWR.n1423 185
R6383 VPWR.n1426 VPWR.n1425 185
R6384 VPWR.n1427 VPWR.n1209 185
R6385 VPWR.n1722 VPWR.n1721 185
R6386 VPWR.n1721 VPWR.n1720 185
R6387 VPWR.n1456 VPWR.n1455 185
R6388 VPWR.n1719 VPWR.n1456 185
R6389 VPWR.n1717 VPWR.n1716 185
R6390 VPWR.n1718 VPWR.n1717 185
R6391 VPWR.n1715 VPWR.n1458 185
R6392 VPWR.n1458 VPWR.n1457 185
R6393 VPWR.n1714 VPWR.n1713 185
R6394 VPWR.n1713 VPWR.n1712 185
R6395 VPWR.n1461 VPWR.n1459 185
R6396 VPWR.n1711 VPWR.n1459 185
R6397 VPWR.n1709 VPWR.n1708 185
R6398 VPWR.n1710 VPWR.n1709 185
R6399 VPWR.n1707 VPWR.n1460 185
R6400 VPWR.n1464 VPWR.n1460 185
R6401 VPWR.n1706 VPWR.n1705 185
R6402 VPWR.n1705 VPWR.n1704 185
R6403 VPWR.n1463 VPWR.n1462 185
R6404 VPWR.n1703 VPWR.n1463 185
R6405 VPWR.n1701 VPWR.n1700 185
R6406 VPWR.n1702 VPWR.n1701 185
R6407 VPWR.n1699 VPWR.n1466 185
R6408 VPWR.n1466 VPWR.n1465 185
R6409 VPWR.n1698 VPWR.n1697 185
R6410 VPWR.n1697 VPWR.n1696 185
R6411 VPWR.n1469 VPWR.n1467 185
R6412 VPWR.n1695 VPWR.n1467 185
R6413 VPWR.n1693 VPWR.n1692 185
R6414 VPWR.n1694 VPWR.n1693 185
R6415 VPWR.n1691 VPWR.n1468 185
R6416 VPWR.n1471 VPWR.n1468 185
R6417 VPWR.n1690 VPWR.n1689 185
R6418 VPWR.n1689 VPWR.n1688 185
R6419 VPWR.n1474 VPWR.n1470 185
R6420 VPWR.n1687 VPWR.n1470 185
R6421 VPWR.n1685 VPWR.n1684 185
R6422 VPWR.n1686 VPWR.n1685 185
R6423 VPWR.n1683 VPWR.n1473 185
R6424 VPWR.n1473 VPWR.n1472 185
R6425 VPWR.n1682 VPWR.n1681 185
R6426 VPWR.n1681 VPWR.n1680 185
R6427 VPWR.n1477 VPWR.n1475 185
R6428 VPWR.n1679 VPWR.n1475 185
R6429 VPWR.n1677 VPWR.n1676 185
R6430 VPWR.n1678 VPWR.n1677 185
R6431 VPWR.n1675 VPWR.n1476 185
R6432 VPWR.n1479 VPWR.n1476 185
R6433 VPWR.n1674 VPWR.n1673 185
R6434 VPWR.n1673 VPWR.n1672 185
R6435 VPWR.n1482 VPWR.n1478 185
R6436 VPWR.n1671 VPWR.n1478 185
R6437 VPWR.n1669 VPWR.n1668 185
R6438 VPWR.n1670 VPWR.n1669 185
R6439 VPWR.n1667 VPWR.n1481 185
R6440 VPWR.n1481 VPWR.n1480 185
R6441 VPWR.n1666 VPWR.n1665 185
R6442 VPWR.n1665 VPWR.n1664 185
R6443 VPWR.n1485 VPWR.n1483 185
R6444 VPWR.n1663 VPWR.n1483 185
R6445 VPWR.n1661 VPWR.n1660 185
R6446 VPWR.n1662 VPWR.n1661 185
R6447 VPWR.n1659 VPWR.n1484 185
R6448 VPWR.n1487 VPWR.n1484 185
R6449 VPWR.n1658 VPWR.n1657 185
R6450 VPWR.n1657 VPWR.n1656 185
R6451 VPWR.n1489 VPWR.n1486 185
R6452 VPWR.n1655 VPWR.n1486 185
R6453 VPWR.n1653 VPWR.n1652 185
R6454 VPWR.n1654 VPWR.n1653 185
R6455 VPWR.n1651 VPWR.n1488 185
R6456 VPWR.n1492 VPWR.n1488 185
R6457 VPWR.n1650 VPWR.n1649 185
R6458 VPWR.n1649 VPWR.n1648 185
R6459 VPWR.n1491 VPWR.n1490 185
R6460 VPWR.n1647 VPWR.n1491 185
R6461 VPWR.n1645 VPWR.n1644 185
R6462 VPWR.n1646 VPWR.n1645 185
R6463 VPWR.n1643 VPWR.n1493 185
R6464 VPWR.n1495 VPWR.n1493 185
R6465 VPWR.n1642 VPWR.n1641 185
R6466 VPWR.n1641 VPWR.n1640 185
R6467 VPWR.n1497 VPWR.n1494 185
R6468 VPWR.n1639 VPWR.n1494 185
R6469 VPWR.n1637 VPWR.n1636 185
R6470 VPWR.n1638 VPWR.n1637 185
R6471 VPWR.n1635 VPWR.n1496 185
R6472 VPWR.n1500 VPWR.n1496 185
R6473 VPWR.n1634 VPWR.n1633 185
R6474 VPWR.n1633 VPWR.n1632 185
R6475 VPWR.n1499 VPWR.n1498 185
R6476 VPWR.n1631 VPWR.n1499 185
R6477 VPWR.n1629 VPWR.n1628 185
R6478 VPWR.n1630 VPWR.n1629 185
R6479 VPWR.n1627 VPWR.n1501 185
R6480 VPWR.n1503 VPWR.n1501 185
R6481 VPWR.n1626 VPWR.n1625 185
R6482 VPWR.n1625 VPWR.n1624 185
R6483 VPWR.n1505 VPWR.n1502 185
R6484 VPWR.n1623 VPWR.n1502 185
R6485 VPWR.n1621 VPWR.n1620 185
R6486 VPWR.n1622 VPWR.n1621 185
R6487 VPWR.n1619 VPWR.n1504 185
R6488 VPWR.n1508 VPWR.n1504 185
R6489 VPWR.n1618 VPWR.n1617 185
R6490 VPWR.n1617 VPWR.n1616 185
R6491 VPWR.n1507 VPWR.n1506 185
R6492 VPWR.n1615 VPWR.n1507 185
R6493 VPWR.n928 VPWR.n725 185
R6494 VPWR.n813 VPWR.n812 185
R6495 VPWR.n815 VPWR.n814 185
R6496 VPWR.n817 VPWR.n816 185
R6497 VPWR.n819 VPWR.n818 185
R6498 VPWR.n821 VPWR.n820 185
R6499 VPWR.n823 VPWR.n822 185
R6500 VPWR.n825 VPWR.n824 185
R6501 VPWR.n827 VPWR.n826 185
R6502 VPWR.n829 VPWR.n828 185
R6503 VPWR.n831 VPWR.n830 185
R6504 VPWR.n833 VPWR.n832 185
R6505 VPWR.n835 VPWR.n834 185
R6506 VPWR.n837 VPWR.n836 185
R6507 VPWR.n839 VPWR.n838 185
R6508 VPWR.n841 VPWR.n840 185
R6509 VPWR.n843 VPWR.n842 185
R6510 VPWR.n845 VPWR.n844 185
R6511 VPWR.n847 VPWR.n846 185
R6512 VPWR.n849 VPWR.n848 185
R6513 VPWR.n851 VPWR.n850 185
R6514 VPWR.n853 VPWR.n852 185
R6515 VPWR.n855 VPWR.n854 185
R6516 VPWR.n857 VPWR.n856 185
R6517 VPWR.n859 VPWR.n858 185
R6518 VPWR.n861 VPWR.n860 185
R6519 VPWR.n863 VPWR.n862 185
R6520 VPWR.n865 VPWR.n864 185
R6521 VPWR.n867 VPWR.n866 185
R6522 VPWR.n869 VPWR.n868 185
R6523 VPWR.n871 VPWR.n870 185
R6524 VPWR.n873 VPWR.n872 185
R6525 VPWR.n875 VPWR.n874 185
R6526 VPWR.n877 VPWR.n876 185
R6527 VPWR.n879 VPWR.n878 185
R6528 VPWR.n881 VPWR.n880 185
R6529 VPWR.n883 VPWR.n882 185
R6530 VPWR.n885 VPWR.n884 185
R6531 VPWR.n887 VPWR.n886 185
R6532 VPWR.n889 VPWR.n888 185
R6533 VPWR.n891 VPWR.n890 185
R6534 VPWR.n893 VPWR.n892 185
R6535 VPWR.n895 VPWR.n894 185
R6536 VPWR.n897 VPWR.n896 185
R6537 VPWR.n899 VPWR.n898 185
R6538 VPWR.n901 VPWR.n900 185
R6539 VPWR.n903 VPWR.n902 185
R6540 VPWR.n905 VPWR.n904 185
R6541 VPWR.n907 VPWR.n906 185
R6542 VPWR.n909 VPWR.n908 185
R6543 VPWR.n911 VPWR.n910 185
R6544 VPWR.n913 VPWR.n912 185
R6545 VPWR.n915 VPWR.n914 185
R6546 VPWR.n917 VPWR.n916 185
R6547 VPWR.n919 VPWR.n918 185
R6548 VPWR.n921 VPWR.n920 185
R6549 VPWR.n923 VPWR.n922 185
R6550 VPWR.n924 VPWR.n811 185
R6551 VPWR.n926 VPWR.n925 185
R6552 VPWR.n782 VPWR.n781 185
R6553 VPWR.n1895 VPWR.n257 185
R6554 VPWR.n1898 VPWR.n1897 185
R6555 VPWR.n259 VPWR.n258 185
R6556 VPWR.n1781 VPWR.n1780 185
R6557 VPWR.n1783 VPWR.n1782 185
R6558 VPWR.n1785 VPWR.n1784 185
R6559 VPWR.n1787 VPWR.n1786 185
R6560 VPWR.n1789 VPWR.n1788 185
R6561 VPWR.n1791 VPWR.n1790 185
R6562 VPWR.n1793 VPWR.n1792 185
R6563 VPWR.n1795 VPWR.n1794 185
R6564 VPWR.n1797 VPWR.n1796 185
R6565 VPWR.n1799 VPWR.n1798 185
R6566 VPWR.n1801 VPWR.n1800 185
R6567 VPWR.n1803 VPWR.n1802 185
R6568 VPWR.n1805 VPWR.n1804 185
R6569 VPWR.n1807 VPWR.n1806 185
R6570 VPWR.n1809 VPWR.n1808 185
R6571 VPWR.n1811 VPWR.n1810 185
R6572 VPWR.n1813 VPWR.n1812 185
R6573 VPWR.n1815 VPWR.n1814 185
R6574 VPWR.n1817 VPWR.n1816 185
R6575 VPWR.n1819 VPWR.n1818 185
R6576 VPWR.n1821 VPWR.n1820 185
R6577 VPWR.n1823 VPWR.n1822 185
R6578 VPWR.n1825 VPWR.n1824 185
R6579 VPWR.n1827 VPWR.n1826 185
R6580 VPWR.n1829 VPWR.n1828 185
R6581 VPWR.n1831 VPWR.n1830 185
R6582 VPWR.n1833 VPWR.n1832 185
R6583 VPWR.n1835 VPWR.n1834 185
R6584 VPWR.n1837 VPWR.n1836 185
R6585 VPWR.n1839 VPWR.n1838 185
R6586 VPWR.n1841 VPWR.n1840 185
R6587 VPWR.n1843 VPWR.n1842 185
R6588 VPWR.n1845 VPWR.n1844 185
R6589 VPWR.n1847 VPWR.n1846 185
R6590 VPWR.n1849 VPWR.n1848 185
R6591 VPWR.n1851 VPWR.n1850 185
R6592 VPWR.n1853 VPWR.n1852 185
R6593 VPWR.n1855 VPWR.n1854 185
R6594 VPWR.n1857 VPWR.n1856 185
R6595 VPWR.n1859 VPWR.n1858 185
R6596 VPWR.n1861 VPWR.n1860 185
R6597 VPWR.n1863 VPWR.n1862 185
R6598 VPWR.n1865 VPWR.n1864 185
R6599 VPWR.n1867 VPWR.n1866 185
R6600 VPWR.n1869 VPWR.n1868 185
R6601 VPWR.n1871 VPWR.n1870 185
R6602 VPWR.n1873 VPWR.n1872 185
R6603 VPWR.n1875 VPWR.n1874 185
R6604 VPWR.n1877 VPWR.n1876 185
R6605 VPWR.n1879 VPWR.n1878 185
R6606 VPWR.n1881 VPWR.n1880 185
R6607 VPWR.n1883 VPWR.n1882 185
R6608 VPWR.n1885 VPWR.n1884 185
R6609 VPWR.n1887 VPWR.n1886 185
R6610 VPWR.n1889 VPWR.n1888 185
R6611 VPWR.n1891 VPWR.n1890 185
R6612 VPWR.n1892 VPWR.n288 185
R6613 VPWR.n1938 VPWR.n1937 185
R6614 VPWR.n1937 VPWR.n1936 185
R6615 VPWR.n1921 VPWR.n1920 185
R6616 VPWR.n1935 VPWR.n1921 185
R6617 VPWR.n1933 VPWR.n1932 185
R6618 VPWR.n1934 VPWR.n1933 185
R6619 VPWR.n1931 VPWR.n1923 185
R6620 VPWR.n1923 VPWR.n1922 185
R6621 VPWR.n1930 VPWR.n1929 185
R6622 VPWR.n1929 VPWR.n1928 185
R6623 VPWR.n1925 VPWR.n1924 185
R6624 VPWR.n1927 VPWR.n1925 185
R6625 VPWR.n598 VPWR.n395 185
R6626 VPWR.n483 VPWR.n482 185
R6627 VPWR.n485 VPWR.n484 185
R6628 VPWR.n487 VPWR.n486 185
R6629 VPWR.n489 VPWR.n488 185
R6630 VPWR.n491 VPWR.n490 185
R6631 VPWR.n493 VPWR.n492 185
R6632 VPWR.n495 VPWR.n494 185
R6633 VPWR.n497 VPWR.n496 185
R6634 VPWR.n499 VPWR.n498 185
R6635 VPWR.n501 VPWR.n500 185
R6636 VPWR.n503 VPWR.n502 185
R6637 VPWR.n505 VPWR.n504 185
R6638 VPWR.n507 VPWR.n506 185
R6639 VPWR.n509 VPWR.n508 185
R6640 VPWR.n511 VPWR.n510 185
R6641 VPWR.n513 VPWR.n512 185
R6642 VPWR.n515 VPWR.n514 185
R6643 VPWR.n517 VPWR.n516 185
R6644 VPWR.n519 VPWR.n518 185
R6645 VPWR.n521 VPWR.n520 185
R6646 VPWR.n523 VPWR.n522 185
R6647 VPWR.n525 VPWR.n524 185
R6648 VPWR.n527 VPWR.n526 185
R6649 VPWR.n529 VPWR.n528 185
R6650 VPWR.n531 VPWR.n530 185
R6651 VPWR.n533 VPWR.n532 185
R6652 VPWR.n535 VPWR.n534 185
R6653 VPWR.n537 VPWR.n536 185
R6654 VPWR.n539 VPWR.n538 185
R6655 VPWR.n541 VPWR.n540 185
R6656 VPWR.n543 VPWR.n542 185
R6657 VPWR.n545 VPWR.n544 185
R6658 VPWR.n547 VPWR.n546 185
R6659 VPWR.n549 VPWR.n548 185
R6660 VPWR.n551 VPWR.n550 185
R6661 VPWR.n553 VPWR.n552 185
R6662 VPWR.n555 VPWR.n554 185
R6663 VPWR.n557 VPWR.n556 185
R6664 VPWR.n559 VPWR.n558 185
R6665 VPWR.n561 VPWR.n560 185
R6666 VPWR.n563 VPWR.n562 185
R6667 VPWR.n565 VPWR.n564 185
R6668 VPWR.n567 VPWR.n566 185
R6669 VPWR.n569 VPWR.n568 185
R6670 VPWR.n571 VPWR.n570 185
R6671 VPWR.n573 VPWR.n572 185
R6672 VPWR.n575 VPWR.n574 185
R6673 VPWR.n577 VPWR.n576 185
R6674 VPWR.n579 VPWR.n578 185
R6675 VPWR.n581 VPWR.n580 185
R6676 VPWR.n583 VPWR.n582 185
R6677 VPWR.n585 VPWR.n584 185
R6678 VPWR.n587 VPWR.n586 185
R6679 VPWR.n589 VPWR.n588 185
R6680 VPWR.n591 VPWR.n590 185
R6681 VPWR.n593 VPWR.n592 185
R6682 VPWR.n594 VPWR.n481 185
R6683 VPWR.n596 VPWR.n595 185
R6684 VPWR.n452 VPWR.n451 185
R6685 VPWR.n1101 VPWR.n1100 185
R6686 VPWR.n1100 VPWR.n1099 185
R6687 VPWR.n1097 VPWR.n1096 185
R6688 VPWR.n1098 VPWR.n1097 185
R6689 VPWR.n1087 VPWR.n1086 185
R6690 VPWR.n1086 VPWR.n1085 185
R6691 VPWR.n1133 VPWR.n1132 185
R6692 VPWR.n1134 VPWR.n1133 185
R6693 VPWR.n1084 VPWR.n1083 185
R6694 VPWR.n1135 VPWR.n1084 185
R6695 VPWR.n1138 VPWR.n1137 185
R6696 VPWR.n1137 VPWR.n1136 185
R6697 VPWR.n1139 VPWR.n1082 185
R6698 VPWR.n1082 VPWR.n1081 185
R6699 VPWR.n1142 VPWR.n1141 185
R6700 VPWR.n1143 VPWR.n1142 185
R6701 VPWR.n1140 VPWR.n1080 185
R6702 VPWR.n1144 VPWR.n1080 185
R6703 VPWR.n1148 VPWR.n1147 185
R6704 VPWR.n1147 VPWR.n1146 185
R6705 VPWR.n1149 VPWR.n1079 185
R6706 VPWR.n1145 VPWR.n1079 185
R6707 VPWR.n1152 VPWR.n1151 185
R6708 VPWR.n1153 VPWR.n1152 185
R6709 VPWR.n1150 VPWR.n1078 185
R6710 VPWR.n1154 VPWR.n1078 185
R6711 VPWR.n1158 VPWR.n1157 185
R6712 VPWR.n1157 VPWR.n1156 185
R6713 VPWR.n1159 VPWR.n1077 185
R6714 VPWR.n1155 VPWR.n1077 185
R6715 VPWR.n1161 VPWR.n1160 185
R6716 VPWR.n1162 VPWR.n1161 185
R6717 VPWR.n1076 VPWR.n1075 185
R6718 VPWR.n1163 VPWR.n1076 185
R6719 VPWR.n1005 VPWR.n1004 185
R6720 VPWR.n1004 VPWR.n1003 185
R6721 VPWR.n1001 VPWR.n1000 185
R6722 VPWR.n1002 VPWR.n1001 185
R6723 VPWR.n997 VPWR.n996 185
R6724 VPWR.n996 VPWR.n995 185
R6725 VPWR.n1031 VPWR.n1030 185
R6726 VPWR.n1032 VPWR.n1031 185
R6727 VPWR.n994 VPWR.n993 185
R6728 VPWR.n1033 VPWR.n994 185
R6729 VPWR.n1036 VPWR.n1035 185
R6730 VPWR.n1035 VPWR.n1034 185
R6731 VPWR.n1037 VPWR.n992 185
R6732 VPWR.n992 VPWR.n991 185
R6733 VPWR.n1040 VPWR.n1039 185
R6734 VPWR.n1041 VPWR.n1040 185
R6735 VPWR.n1038 VPWR.n990 185
R6736 VPWR.n1042 VPWR.n990 185
R6737 VPWR.n1046 VPWR.n1045 185
R6738 VPWR.n1045 VPWR.n1044 185
R6739 VPWR.n1047 VPWR.n989 185
R6740 VPWR.n1043 VPWR.n989 185
R6741 VPWR.n1050 VPWR.n1049 185
R6742 VPWR.n1051 VPWR.n1050 185
R6743 VPWR.n1048 VPWR.n988 185
R6744 VPWR.n1052 VPWR.n988 185
R6745 VPWR.n1056 VPWR.n1055 185
R6746 VPWR.n1055 VPWR.n1054 185
R6747 VPWR.n1057 VPWR.n987 185
R6748 VPWR.n1053 VPWR.n987 185
R6749 VPWR.n1059 VPWR.n1058 185
R6750 VPWR.n1060 VPWR.n1059 185
R6751 VPWR.n986 VPWR.n985 185
R6752 VPWR.n1061 VPWR.n986 185
R6753 VPWR.n2332 VPWR.n2331 185
R6754 VPWR.n2330 VPWR.n2293 185
R6755 VPWR.n2329 VPWR.n2328 185
R6756 VPWR.n2327 VPWR.n2326 185
R6757 VPWR.n2325 VPWR.n2324 185
R6758 VPWR.n2323 VPWR.n2322 185
R6759 VPWR.n2321 VPWR.n2320 185
R6760 VPWR.n2319 VPWR.n2318 185
R6761 VPWR.n2317 VPWR.n2316 185
R6762 VPWR.n2315 VPWR.n2314 185
R6763 VPWR.n2313 VPWR.n2312 185
R6764 VPWR.n2311 VPWR.n2310 185
R6765 VPWR.n2309 VPWR.n2308 185
R6766 VPWR.n2307 VPWR.n2306 185
R6767 VPWR.n2305 VPWR.n2304 185
R6768 VPWR.n2303 VPWR.n2302 185
R6769 VPWR.n2301 VPWR.n2300 185
R6770 VPWR.n2299 VPWR.n2298 185
R6771 VPWR.n2297 VPWR.n2296 185
R6772 VPWR.n2295 VPWR.n2294 185
R6773 VPWR.n2282 VPWR.n2281 185
R6774 VPWR.n2333 VPWR.n2332 185
R6775 VPWR.n1529 VPWR.t565 131.389
R6776 VPWR.n1587 VPWR.t554 131.389
R6777 VPWR VPWR.n1529 128.754
R6778 VPWR VPWR.n1587 128.754
R6779 VPWR.n2023 VPWR.n2022 116.112
R6780 VPWR.n2030 VPWR.n2017 116.112
R6781 VPWR.n2033 VPWR.n2032 116.112
R6782 VPWR.n2041 VPWR.n2040 116.112
R6783 VPWR.n2043 VPWR.n2042 116.112
R6784 VPWR.n2052 VPWR.n2050 116.112
R6785 VPWR.n2060 VPWR.n2059 116.112
R6786 VPWR.n2062 VPWR.n2061 116.112
R6787 VPWR.n2069 VPWR.n2068 116.112
R6788 VPWR.n1720 VPWR.n1719 116.112
R6789 VPWR.n1718 VPWR.n1457 116.112
R6790 VPWR.n1711 VPWR.n1710 116.112
R6791 VPWR.n1704 VPWR.n1703 116.112
R6792 VPWR.n1702 VPWR.n1465 116.112
R6793 VPWR.n1686 VPWR.n1472 116.112
R6794 VPWR.n1670 VPWR.n1480 116.112
R6795 VPWR.n1656 VPWR.n1487 116.112
R6796 VPWR.n1648 VPWR.n1647 116.112
R6797 VPWR.n1632 VPWR.n1631 116.112
R6798 VPWR.n1616 VPWR.n1615 116.112
R6799 VPWR.n1936 VPWR.n1935 116.112
R6800 VPWR.n1934 VPWR.n1922 116.112
R6801 VPWR.n1928 VPWR.n1927 116.112
R6802 VPWR.n1099 VPWR.n1098 116.112
R6803 VPWR.n1134 VPWR.n1085 116.112
R6804 VPWR.n1136 VPWR.n1135 116.112
R6805 VPWR.n1143 VPWR.n1081 116.112
R6806 VPWR.n1146 VPWR.n1145 116.112
R6807 VPWR.n1156 VPWR.n1155 116.112
R6808 VPWR.n1163 VPWR.n1162 116.112
R6809 VPWR.n1003 VPWR.n1002 116.112
R6810 VPWR.n1032 VPWR.n995 116.112
R6811 VPWR.n1034 VPWR.n1033 116.112
R6812 VPWR.n1041 VPWR.n991 116.112
R6813 VPWR.n1044 VPWR.n1043 116.112
R6814 VPWR.n1054 VPWR.n1053 116.112
R6815 VPWR.n1061 VPWR.n1060 116.112
R6816 VPWR.n2341 VPWR 112.511
R6817 VPWR.n2021 VPWR.n2020 97.7783
R6818 VPWR.n2024 VPWR.n2020 97.7783
R6819 VPWR.n2024 VPWR.n2018 97.7783
R6820 VPWR.n2029 VPWR.n2018 97.7783
R6821 VPWR.n2029 VPWR.n2016 97.7783
R6822 VPWR.n2034 VPWR.n2016 97.7783
R6823 VPWR.n2034 VPWR.n2015 97.7783
R6824 VPWR.n2039 VPWR.n2015 97.7783
R6825 VPWR.n2039 VPWR.n2014 97.7783
R6826 VPWR.n2044 VPWR.n2014 97.7783
R6827 VPWR.n2044 VPWR.n2013 97.7783
R6828 VPWR.n2048 VPWR.n2013 97.7783
R6829 VPWR.n2048 VPWR.n2012 97.7783
R6830 VPWR.n2053 VPWR.n2012 97.7783
R6831 VPWR.n2053 VPWR.n2010 97.7783
R6832 VPWR.n2058 VPWR.n2010 97.7783
R6833 VPWR.n2058 VPWR.n2009 97.7783
R6834 VPWR.n2063 VPWR.n2009 97.7783
R6835 VPWR.n2063 VPWR.n2008 97.7783
R6836 VPWR.n2067 VPWR.n2008 97.7783
R6837 VPWR.n2067 VPWR.n2007 97.7783
R6838 VPWR.n2070 VPWR.n2007 97.7783
R6839 VPWR.n2133 VPWR.n2095 97.7783
R6840 VPWR.n2130 VPWR.n2129 97.7783
R6841 VPWR.n2126 VPWR.n2125 97.7783
R6842 VPWR.n2122 VPWR.n2121 97.7783
R6843 VPWR.n2118 VPWR.n2117 97.7783
R6844 VPWR.n2114 VPWR.n2113 97.7783
R6845 VPWR.n2110 VPWR.n2109 97.7783
R6846 VPWR.n2106 VPWR.n2105 97.7783
R6847 VPWR.n2102 VPWR.n2101 97.7783
R6848 VPWR.n2098 VPWR.n2097 97.7783
R6849 VPWR.n2135 VPWR.n2084 97.7783
R6850 VPWR.n2199 VPWR.n2161 97.7783
R6851 VPWR.n2196 VPWR.n2195 97.7783
R6852 VPWR.n2192 VPWR.n2191 97.7783
R6853 VPWR.n2188 VPWR.n2187 97.7783
R6854 VPWR.n2184 VPWR.n2183 97.7783
R6855 VPWR.n2180 VPWR.n2179 97.7783
R6856 VPWR.n2176 VPWR.n2175 97.7783
R6857 VPWR.n2172 VPWR.n2171 97.7783
R6858 VPWR.n2168 VPWR.n2167 97.7783
R6859 VPWR.n2164 VPWR.n2163 97.7783
R6860 VPWR.n2201 VPWR.n2150 97.7783
R6861 VPWR.n2265 VPWR.n2227 97.7783
R6862 VPWR.n2262 VPWR.n2261 97.7783
R6863 VPWR.n2258 VPWR.n2257 97.7783
R6864 VPWR.n2254 VPWR.n2253 97.7783
R6865 VPWR.n2250 VPWR.n2249 97.7783
R6866 VPWR.n2246 VPWR.n2245 97.7783
R6867 VPWR.n2242 VPWR.n2241 97.7783
R6868 VPWR.n2238 VPWR.n2237 97.7783
R6869 VPWR.n2234 VPWR.n2233 97.7783
R6870 VPWR.n2230 VPWR.n2229 97.7783
R6871 VPWR.n2267 VPWR.n2216 97.7783
R6872 VPWR.n1432 VPWR.n1178 97.7783
R6873 VPWR.n1315 VPWR.n1180 97.7783
R6874 VPWR.n1319 VPWR.n1318 97.7783
R6875 VPWR.n1323 VPWR.n1322 97.7783
R6876 VPWR.n1327 VPWR.n1326 97.7783
R6877 VPWR.n1331 VPWR.n1330 97.7783
R6878 VPWR.n1335 VPWR.n1334 97.7783
R6879 VPWR.n1339 VPWR.n1338 97.7783
R6880 VPWR.n1343 VPWR.n1342 97.7783
R6881 VPWR.n1347 VPWR.n1346 97.7783
R6882 VPWR.n1351 VPWR.n1350 97.7783
R6883 VPWR.n1355 VPWR.n1354 97.7783
R6884 VPWR.n1359 VPWR.n1358 97.7783
R6885 VPWR.n1363 VPWR.n1362 97.7783
R6886 VPWR.n1367 VPWR.n1366 97.7783
R6887 VPWR.n1371 VPWR.n1370 97.7783
R6888 VPWR.n1375 VPWR.n1374 97.7783
R6889 VPWR.n1379 VPWR.n1378 97.7783
R6890 VPWR.n1383 VPWR.n1382 97.7783
R6891 VPWR.n1387 VPWR.n1386 97.7783
R6892 VPWR.n1391 VPWR.n1390 97.7783
R6893 VPWR.n1395 VPWR.n1394 97.7783
R6894 VPWR.n1399 VPWR.n1398 97.7783
R6895 VPWR.n1403 VPWR.n1402 97.7783
R6896 VPWR.n1407 VPWR.n1406 97.7783
R6897 VPWR.n1411 VPWR.n1410 97.7783
R6898 VPWR.n1415 VPWR.n1414 97.7783
R6899 VPWR.n1419 VPWR.n1418 97.7783
R6900 VPWR.n1423 VPWR.n1422 97.7783
R6901 VPWR.n1425 VPWR.n1209 97.7783
R6902 VPWR.n1721 VPWR.n1454 97.7783
R6903 VPWR.n1721 VPWR.n1456 97.7783
R6904 VPWR.n1717 VPWR.n1456 97.7783
R6905 VPWR.n1717 VPWR.n1458 97.7783
R6906 VPWR.n1713 VPWR.n1458 97.7783
R6907 VPWR.n1713 VPWR.n1459 97.7783
R6908 VPWR.n1709 VPWR.n1459 97.7783
R6909 VPWR.n1709 VPWR.n1460 97.7783
R6910 VPWR.n1705 VPWR.n1460 97.7783
R6911 VPWR.n1705 VPWR.n1463 97.7783
R6912 VPWR.n1701 VPWR.n1463 97.7783
R6913 VPWR.n1701 VPWR.n1466 97.7783
R6914 VPWR.n1697 VPWR.n1466 97.7783
R6915 VPWR.n1697 VPWR.n1467 97.7783
R6916 VPWR.n1693 VPWR.n1467 97.7783
R6917 VPWR.n1693 VPWR.n1468 97.7783
R6918 VPWR.n1689 VPWR.n1468 97.7783
R6919 VPWR.n1689 VPWR.n1470 97.7783
R6920 VPWR.n1685 VPWR.n1470 97.7783
R6921 VPWR.n1685 VPWR.n1473 97.7783
R6922 VPWR.n1681 VPWR.n1473 97.7783
R6923 VPWR.n1681 VPWR.n1475 97.7783
R6924 VPWR.n1677 VPWR.n1475 97.7783
R6925 VPWR.n1677 VPWR.n1476 97.7783
R6926 VPWR.n1673 VPWR.n1476 97.7783
R6927 VPWR.n1673 VPWR.n1478 97.7783
R6928 VPWR.n1669 VPWR.n1478 97.7783
R6929 VPWR.n1669 VPWR.n1481 97.7783
R6930 VPWR.n1665 VPWR.n1481 97.7783
R6931 VPWR.n1665 VPWR.n1483 97.7783
R6932 VPWR.n1661 VPWR.n1483 97.7783
R6933 VPWR.n1661 VPWR.n1484 97.7783
R6934 VPWR.n1657 VPWR.n1484 97.7783
R6935 VPWR.n1657 VPWR.n1486 97.7783
R6936 VPWR.n1653 VPWR.n1486 97.7783
R6937 VPWR.n1653 VPWR.n1488 97.7783
R6938 VPWR.n1649 VPWR.n1488 97.7783
R6939 VPWR.n1649 VPWR.n1491 97.7783
R6940 VPWR.n1645 VPWR.n1491 97.7783
R6941 VPWR.n1645 VPWR.n1493 97.7783
R6942 VPWR.n1641 VPWR.n1493 97.7783
R6943 VPWR.n1641 VPWR.n1494 97.7783
R6944 VPWR.n1637 VPWR.n1494 97.7783
R6945 VPWR.n1637 VPWR.n1496 97.7783
R6946 VPWR.n1633 VPWR.n1496 97.7783
R6947 VPWR.n1633 VPWR.n1499 97.7783
R6948 VPWR.n1629 VPWR.n1499 97.7783
R6949 VPWR.n1629 VPWR.n1501 97.7783
R6950 VPWR.n1625 VPWR.n1501 97.7783
R6951 VPWR.n1625 VPWR.n1502 97.7783
R6952 VPWR.n1621 VPWR.n1502 97.7783
R6953 VPWR.n1621 VPWR.n1504 97.7783
R6954 VPWR.n1617 VPWR.n1504 97.7783
R6955 VPWR.n1617 VPWR.n1507 97.7783
R6956 VPWR.n1614 VPWR.n1507 97.7783
R6957 VPWR.n812 VPWR.n725 97.7783
R6958 VPWR.n816 VPWR.n815 97.7783
R6959 VPWR.n820 VPWR.n819 97.7783
R6960 VPWR.n824 VPWR.n823 97.7783
R6961 VPWR.n828 VPWR.n827 97.7783
R6962 VPWR.n832 VPWR.n831 97.7783
R6963 VPWR.n836 VPWR.n835 97.7783
R6964 VPWR.n840 VPWR.n839 97.7783
R6965 VPWR.n844 VPWR.n843 97.7783
R6966 VPWR.n848 VPWR.n847 97.7783
R6967 VPWR.n852 VPWR.n851 97.7783
R6968 VPWR.n856 VPWR.n855 97.7783
R6969 VPWR.n860 VPWR.n859 97.7783
R6970 VPWR.n864 VPWR.n863 97.7783
R6971 VPWR.n868 VPWR.n867 97.7783
R6972 VPWR.n872 VPWR.n871 97.7783
R6973 VPWR.n876 VPWR.n875 97.7783
R6974 VPWR.n880 VPWR.n879 97.7783
R6975 VPWR.n884 VPWR.n883 97.7783
R6976 VPWR.n888 VPWR.n887 97.7783
R6977 VPWR.n892 VPWR.n891 97.7783
R6978 VPWR.n896 VPWR.n895 97.7783
R6979 VPWR.n900 VPWR.n899 97.7783
R6980 VPWR.n904 VPWR.n903 97.7783
R6981 VPWR.n908 VPWR.n907 97.7783
R6982 VPWR.n912 VPWR.n911 97.7783
R6983 VPWR.n916 VPWR.n915 97.7783
R6984 VPWR.n920 VPWR.n919 97.7783
R6985 VPWR.n922 VPWR.n811 97.7783
R6986 VPWR.n926 VPWR.n782 97.7783
R6987 VPWR.n1897 VPWR.n257 97.7783
R6988 VPWR.n1780 VPWR.n259 97.7783
R6989 VPWR.n1784 VPWR.n1783 97.7783
R6990 VPWR.n1788 VPWR.n1787 97.7783
R6991 VPWR.n1792 VPWR.n1791 97.7783
R6992 VPWR.n1796 VPWR.n1795 97.7783
R6993 VPWR.n1800 VPWR.n1799 97.7783
R6994 VPWR.n1804 VPWR.n1803 97.7783
R6995 VPWR.n1808 VPWR.n1807 97.7783
R6996 VPWR.n1812 VPWR.n1811 97.7783
R6997 VPWR.n1816 VPWR.n1815 97.7783
R6998 VPWR.n1820 VPWR.n1819 97.7783
R6999 VPWR.n1824 VPWR.n1823 97.7783
R7000 VPWR.n1828 VPWR.n1827 97.7783
R7001 VPWR.n1832 VPWR.n1831 97.7783
R7002 VPWR.n1836 VPWR.n1835 97.7783
R7003 VPWR.n1840 VPWR.n1839 97.7783
R7004 VPWR.n1844 VPWR.n1843 97.7783
R7005 VPWR.n1848 VPWR.n1847 97.7783
R7006 VPWR.n1852 VPWR.n1851 97.7783
R7007 VPWR.n1856 VPWR.n1855 97.7783
R7008 VPWR.n1860 VPWR.n1859 97.7783
R7009 VPWR.n1864 VPWR.n1863 97.7783
R7010 VPWR.n1868 VPWR.n1867 97.7783
R7011 VPWR.n1872 VPWR.n1871 97.7783
R7012 VPWR.n1876 VPWR.n1875 97.7783
R7013 VPWR.n1880 VPWR.n1879 97.7783
R7014 VPWR.n1884 VPWR.n1883 97.7783
R7015 VPWR.n1888 VPWR.n1887 97.7783
R7016 VPWR.n1890 VPWR.n288 97.7783
R7017 VPWR.n1937 VPWR.n1919 97.7783
R7018 VPWR.n1937 VPWR.n1921 97.7783
R7019 VPWR.n1933 VPWR.n1921 97.7783
R7020 VPWR.n1933 VPWR.n1923 97.7783
R7021 VPWR.n1929 VPWR.n1923 97.7783
R7022 VPWR.n1929 VPWR.n1925 97.7783
R7023 VPWR.n1926 VPWR.n1925 97.7783
R7024 VPWR.n482 VPWR.n395 97.7783
R7025 VPWR.n486 VPWR.n485 97.7783
R7026 VPWR.n490 VPWR.n489 97.7783
R7027 VPWR.n494 VPWR.n493 97.7783
R7028 VPWR.n498 VPWR.n497 97.7783
R7029 VPWR.n502 VPWR.n501 97.7783
R7030 VPWR.n506 VPWR.n505 97.7783
R7031 VPWR.n510 VPWR.n509 97.7783
R7032 VPWR.n514 VPWR.n513 97.7783
R7033 VPWR.n518 VPWR.n517 97.7783
R7034 VPWR.n522 VPWR.n521 97.7783
R7035 VPWR.n526 VPWR.n525 97.7783
R7036 VPWR.n530 VPWR.n529 97.7783
R7037 VPWR.n534 VPWR.n533 97.7783
R7038 VPWR.n538 VPWR.n537 97.7783
R7039 VPWR.n542 VPWR.n541 97.7783
R7040 VPWR.n546 VPWR.n545 97.7783
R7041 VPWR.n550 VPWR.n549 97.7783
R7042 VPWR.n554 VPWR.n553 97.7783
R7043 VPWR.n558 VPWR.n557 97.7783
R7044 VPWR.n562 VPWR.n561 97.7783
R7045 VPWR.n566 VPWR.n565 97.7783
R7046 VPWR.n570 VPWR.n569 97.7783
R7047 VPWR.n574 VPWR.n573 97.7783
R7048 VPWR.n578 VPWR.n577 97.7783
R7049 VPWR.n582 VPWR.n581 97.7783
R7050 VPWR.n586 VPWR.n585 97.7783
R7051 VPWR.n590 VPWR.n589 97.7783
R7052 VPWR.n592 VPWR.n481 97.7783
R7053 VPWR.n596 VPWR.n452 97.7783
R7054 VPWR.n1100 VPWR.n1095 97.7783
R7055 VPWR.n1100 VPWR.n1097 97.7783
R7056 VPWR.n1097 VPWR.n1086 97.7783
R7057 VPWR.n1133 VPWR.n1086 97.7783
R7058 VPWR.n1133 VPWR.n1084 97.7783
R7059 VPWR.n1137 VPWR.n1084 97.7783
R7060 VPWR.n1137 VPWR.n1082 97.7783
R7061 VPWR.n1142 VPWR.n1082 97.7783
R7062 VPWR.n1142 VPWR.n1080 97.7783
R7063 VPWR.n1147 VPWR.n1080 97.7783
R7064 VPWR.n1147 VPWR.n1079 97.7783
R7065 VPWR.n1152 VPWR.n1079 97.7783
R7066 VPWR.n1152 VPWR.n1078 97.7783
R7067 VPWR.n1157 VPWR.n1078 97.7783
R7068 VPWR.n1157 VPWR.n1077 97.7783
R7069 VPWR.n1161 VPWR.n1077 97.7783
R7070 VPWR.n1161 VPWR.n1076 97.7783
R7071 VPWR.n1164 VPWR.n1076 97.7783
R7072 VPWR.n1004 VPWR.n999 97.7783
R7073 VPWR.n1004 VPWR.n1001 97.7783
R7074 VPWR.n1001 VPWR.n996 97.7783
R7075 VPWR.n1031 VPWR.n996 97.7783
R7076 VPWR.n1031 VPWR.n994 97.7783
R7077 VPWR.n1035 VPWR.n994 97.7783
R7078 VPWR.n1035 VPWR.n992 97.7783
R7079 VPWR.n1040 VPWR.n992 97.7783
R7080 VPWR.n1040 VPWR.n990 97.7783
R7081 VPWR.n1045 VPWR.n990 97.7783
R7082 VPWR.n1045 VPWR.n989 97.7783
R7083 VPWR.n1050 VPWR.n989 97.7783
R7084 VPWR.n1050 VPWR.n988 97.7783
R7085 VPWR.n1055 VPWR.n988 97.7783
R7086 VPWR.n1055 VPWR.n987 97.7783
R7087 VPWR.n1059 VPWR.n987 97.7783
R7088 VPWR.n1059 VPWR.n986 97.7783
R7089 VPWR.n1062 VPWR.n986 97.7783
R7090 VPWR.n2331 VPWR.n2293 97.7783
R7091 VPWR.n2328 VPWR.n2327 97.7783
R7092 VPWR.n2324 VPWR.n2323 97.7783
R7093 VPWR.n2320 VPWR.n2319 97.7783
R7094 VPWR.n2316 VPWR.n2315 97.7783
R7095 VPWR.n2312 VPWR.n2311 97.7783
R7096 VPWR.n2308 VPWR.n2307 97.7783
R7097 VPWR.n2304 VPWR.n2303 97.7783
R7098 VPWR.n2300 VPWR.n2299 97.7783
R7099 VPWR.n2296 VPWR.n2295 97.7783
R7100 VPWR.n2333 VPWR.n2282 97.7783
R7101 VPWR.n1430 VPWR.t21 74.6187
R7102 VPWR.n1430 VPWR.t6 74.6187
R7103 VPWR.n928 VPWR.t17 74.6187
R7104 VPWR.n928 VPWR.t94 74.6187
R7105 VPWR.n1895 VPWR.t71 74.6187
R7106 VPWR.n1895 VPWR.t27 74.6187
R7107 VPWR.n598 VPWR.t102 74.6187
R7108 VPWR.n598 VPWR.t9 74.6187
R7109 VPWR.n2134 VPWR.n2085 73.1661
R7110 VPWR.n2134 VPWR.n2086 73.1661
R7111 VPWR.n2134 VPWR.n2087 73.1661
R7112 VPWR.n2134 VPWR.n2088 73.1661
R7113 VPWR.n2134 VPWR.n2089 73.1661
R7114 VPWR.n2134 VPWR.n2090 73.1661
R7115 VPWR.n2134 VPWR.n2091 73.1661
R7116 VPWR.n2134 VPWR.n2092 73.1661
R7117 VPWR.n2134 VPWR.n2093 73.1661
R7118 VPWR.n2134 VPWR.n2094 73.1661
R7119 VPWR.n2200 VPWR.n2151 73.1661
R7120 VPWR.n2200 VPWR.n2152 73.1661
R7121 VPWR.n2200 VPWR.n2153 73.1661
R7122 VPWR.n2200 VPWR.n2154 73.1661
R7123 VPWR.n2200 VPWR.n2155 73.1661
R7124 VPWR.n2200 VPWR.n2156 73.1661
R7125 VPWR.n2200 VPWR.n2157 73.1661
R7126 VPWR.n2200 VPWR.n2158 73.1661
R7127 VPWR.n2200 VPWR.n2159 73.1661
R7128 VPWR.n2200 VPWR.n2160 73.1661
R7129 VPWR.n2266 VPWR.n2217 73.1661
R7130 VPWR.n2266 VPWR.n2218 73.1661
R7131 VPWR.n2266 VPWR.n2219 73.1661
R7132 VPWR.n2266 VPWR.n2220 73.1661
R7133 VPWR.n2266 VPWR.n2221 73.1661
R7134 VPWR.n2266 VPWR.n2222 73.1661
R7135 VPWR.n2266 VPWR.n2223 73.1661
R7136 VPWR.n2266 VPWR.n2224 73.1661
R7137 VPWR.n2266 VPWR.n2225 73.1661
R7138 VPWR.n2266 VPWR.n2226 73.1661
R7139 VPWR.n1431 VPWR.n1430 73.1661
R7140 VPWR.n1430 VPWR.n1181 73.1661
R7141 VPWR.n1430 VPWR.n1182 73.1661
R7142 VPWR.n1430 VPWR.n1183 73.1661
R7143 VPWR.n1430 VPWR.n1184 73.1661
R7144 VPWR.n1430 VPWR.n1185 73.1661
R7145 VPWR.n1430 VPWR.n1186 73.1661
R7146 VPWR.n1430 VPWR.n1187 73.1661
R7147 VPWR.n1430 VPWR.n1188 73.1661
R7148 VPWR.n1430 VPWR.n1189 73.1661
R7149 VPWR.n1430 VPWR.n1190 73.1661
R7150 VPWR.n1430 VPWR.n1191 73.1661
R7151 VPWR.n1430 VPWR.n1192 73.1661
R7152 VPWR.n1430 VPWR.n1193 73.1661
R7153 VPWR.n1430 VPWR.n1194 73.1661
R7154 VPWR.n1430 VPWR.n1195 73.1661
R7155 VPWR.n1430 VPWR.n1196 73.1661
R7156 VPWR.n1430 VPWR.n1197 73.1661
R7157 VPWR.n1430 VPWR.n1198 73.1661
R7158 VPWR.n1430 VPWR.n1199 73.1661
R7159 VPWR.n1430 VPWR.n1200 73.1661
R7160 VPWR.n1430 VPWR.n1201 73.1661
R7161 VPWR.n1430 VPWR.n1202 73.1661
R7162 VPWR.n1430 VPWR.n1203 73.1661
R7163 VPWR.n1430 VPWR.n1204 73.1661
R7164 VPWR.n1430 VPWR.n1205 73.1661
R7165 VPWR.n1430 VPWR.n1206 73.1661
R7166 VPWR.n1430 VPWR.n1207 73.1661
R7167 VPWR.n1430 VPWR.n1208 73.1661
R7168 VPWR.n1430 VPWR.n1429 73.1661
R7169 VPWR.n928 VPWR.n783 73.1661
R7170 VPWR.n928 VPWR.n784 73.1661
R7171 VPWR.n928 VPWR.n785 73.1661
R7172 VPWR.n928 VPWR.n786 73.1661
R7173 VPWR.n928 VPWR.n787 73.1661
R7174 VPWR.n928 VPWR.n788 73.1661
R7175 VPWR.n928 VPWR.n789 73.1661
R7176 VPWR.n928 VPWR.n790 73.1661
R7177 VPWR.n928 VPWR.n791 73.1661
R7178 VPWR.n928 VPWR.n792 73.1661
R7179 VPWR.n928 VPWR.n793 73.1661
R7180 VPWR.n928 VPWR.n794 73.1661
R7181 VPWR.n928 VPWR.n795 73.1661
R7182 VPWR.n928 VPWR.n796 73.1661
R7183 VPWR.n928 VPWR.n797 73.1661
R7184 VPWR.n928 VPWR.n798 73.1661
R7185 VPWR.n928 VPWR.n799 73.1661
R7186 VPWR.n928 VPWR.n800 73.1661
R7187 VPWR.n928 VPWR.n801 73.1661
R7188 VPWR.n928 VPWR.n802 73.1661
R7189 VPWR.n928 VPWR.n803 73.1661
R7190 VPWR.n928 VPWR.n804 73.1661
R7191 VPWR.n928 VPWR.n805 73.1661
R7192 VPWR.n928 VPWR.n806 73.1661
R7193 VPWR.n928 VPWR.n807 73.1661
R7194 VPWR.n928 VPWR.n808 73.1661
R7195 VPWR.n928 VPWR.n809 73.1661
R7196 VPWR.n928 VPWR.n810 73.1661
R7197 VPWR.n928 VPWR.n927 73.1661
R7198 VPWR.n929 VPWR.n928 73.1661
R7199 VPWR.n1896 VPWR.n1895 73.1661
R7200 VPWR.n1895 VPWR.n260 73.1661
R7201 VPWR.n1895 VPWR.n261 73.1661
R7202 VPWR.n1895 VPWR.n262 73.1661
R7203 VPWR.n1895 VPWR.n263 73.1661
R7204 VPWR.n1895 VPWR.n264 73.1661
R7205 VPWR.n1895 VPWR.n265 73.1661
R7206 VPWR.n1895 VPWR.n266 73.1661
R7207 VPWR.n1895 VPWR.n267 73.1661
R7208 VPWR.n1895 VPWR.n268 73.1661
R7209 VPWR.n1895 VPWR.n269 73.1661
R7210 VPWR.n1895 VPWR.n270 73.1661
R7211 VPWR.n1895 VPWR.n271 73.1661
R7212 VPWR.n1895 VPWR.n272 73.1661
R7213 VPWR.n1895 VPWR.n273 73.1661
R7214 VPWR.n1895 VPWR.n274 73.1661
R7215 VPWR.n1895 VPWR.n275 73.1661
R7216 VPWR.n1895 VPWR.n276 73.1661
R7217 VPWR.n1895 VPWR.n277 73.1661
R7218 VPWR.n1895 VPWR.n278 73.1661
R7219 VPWR.n1895 VPWR.n279 73.1661
R7220 VPWR.n1895 VPWR.n280 73.1661
R7221 VPWR.n1895 VPWR.n281 73.1661
R7222 VPWR.n1895 VPWR.n282 73.1661
R7223 VPWR.n1895 VPWR.n283 73.1661
R7224 VPWR.n1895 VPWR.n284 73.1661
R7225 VPWR.n1895 VPWR.n285 73.1661
R7226 VPWR.n1895 VPWR.n286 73.1661
R7227 VPWR.n1895 VPWR.n287 73.1661
R7228 VPWR.n1895 VPWR.n1894 73.1661
R7229 VPWR.n598 VPWR.n453 73.1661
R7230 VPWR.n598 VPWR.n454 73.1661
R7231 VPWR.n598 VPWR.n455 73.1661
R7232 VPWR.n598 VPWR.n456 73.1661
R7233 VPWR.n598 VPWR.n457 73.1661
R7234 VPWR.n598 VPWR.n458 73.1661
R7235 VPWR.n598 VPWR.n459 73.1661
R7236 VPWR.n598 VPWR.n460 73.1661
R7237 VPWR.n598 VPWR.n461 73.1661
R7238 VPWR.n598 VPWR.n462 73.1661
R7239 VPWR.n598 VPWR.n463 73.1661
R7240 VPWR.n598 VPWR.n464 73.1661
R7241 VPWR.n598 VPWR.n465 73.1661
R7242 VPWR.n598 VPWR.n466 73.1661
R7243 VPWR.n598 VPWR.n467 73.1661
R7244 VPWR.n598 VPWR.n468 73.1661
R7245 VPWR.n598 VPWR.n469 73.1661
R7246 VPWR.n598 VPWR.n470 73.1661
R7247 VPWR.n598 VPWR.n471 73.1661
R7248 VPWR.n598 VPWR.n472 73.1661
R7249 VPWR.n598 VPWR.n473 73.1661
R7250 VPWR.n598 VPWR.n474 73.1661
R7251 VPWR.n598 VPWR.n475 73.1661
R7252 VPWR.n598 VPWR.n476 73.1661
R7253 VPWR.n598 VPWR.n477 73.1661
R7254 VPWR.n598 VPWR.n478 73.1661
R7255 VPWR.n598 VPWR.n479 73.1661
R7256 VPWR.n598 VPWR.n480 73.1661
R7257 VPWR.n598 VPWR.n597 73.1661
R7258 VPWR.n599 VPWR.n598 73.1661
R7259 VPWR.n2332 VPWR.n2283 73.1661
R7260 VPWR.n2332 VPWR.n2284 73.1661
R7261 VPWR.n2332 VPWR.n2285 73.1661
R7262 VPWR.n2332 VPWR.n2286 73.1661
R7263 VPWR.n2332 VPWR.n2287 73.1661
R7264 VPWR.n2332 VPWR.n2288 73.1661
R7265 VPWR.n2332 VPWR.n2289 73.1661
R7266 VPWR.n2332 VPWR.n2290 73.1661
R7267 VPWR.n2332 VPWR.n2291 73.1661
R7268 VPWR.n2332 VPWR.n2292 73.1661
R7269 VPWR.n1940 VPWR.n1939 69.1205
R7270 VPWR.n1530 VPWR 64.7534
R7271 VPWR.n1588 VPWR 64.7534
R7272 VPWR.n371 VPWR.t458 63.8431
R7273 VPWR.n371 VPWR.t460 63.8431
R7274 VPWR.n376 VPWR.t463 63.8431
R7275 VPWR.n376 VPWR.t462 63.8431
R7276 VPWR.n381 VPWR.t432 63.8431
R7277 VPWR.n381 VPWR.t431 63.8431
R7278 VPWR.n386 VPWR.t400 63.8431
R7279 VPWR.n386 VPWR.t402 63.8431
R7280 VPWR.n1993 VPWR.t1 63.8431
R7281 VPWR.n1993 VPWR.t551 63.8431
R7282 VPWR.n1252 VPWR.t24 63.8431
R7283 VPWR.n1252 VPWR.t25 63.8431
R7284 VPWR.n1257 VPWR.t485 63.8431
R7285 VPWR.n1257 VPWR.t488 63.8431
R7286 VPWR.n1262 VPWR.t569 63.8431
R7287 VPWR.n1262 VPWR.t567 63.8431
R7288 VPWR.n1267 VPWR.t592 63.8431
R7289 VPWR.n1267 VPWR.t591 63.8431
R7290 VPWR.n5 VPWR.t587 63.8431
R7291 VPWR.n5 VPWR.t585 63.8431
R7292 VPWR.n10 VPWR.t545 63.8431
R7293 VPWR.n10 VPWR.t546 63.8431
R7294 VPWR.n15 VPWR.t576 63.8431
R7295 VPWR.n15 VPWR.t574 63.8431
R7296 VPWR.n20 VPWR.t479 63.8431
R7297 VPWR.n20 VPWR.t480 63.8431
R7298 VPWR.n1296 VPWR.t413 63.8431
R7299 VPWR.n1296 VPWR.t26 63.8431
R7300 VPWR.n1226 VPWR.t593 63.8431
R7301 VPWR.n1226 VPWR.t514 63.8431
R7302 VPWR.n1541 VPWR.t211 63.8431
R7303 VPWR.n1541 VPWR.t369 63.8431
R7304 VPWR.n1531 VPWR.t81 63.8431
R7305 VPWR.n1531 VPWR.t53 63.8431
R7306 VPWR.n1533 VPWR.t54 63.8431
R7307 VPWR.n1533 VPWR.t65 63.8431
R7308 VPWR.n1535 VPWR.t66 63.8431
R7309 VPWR.n1535 VPWR.t111 63.8431
R7310 VPWR.n1537 VPWR.t112 63.8431
R7311 VPWR.n1537 VPWR.t162 63.8431
R7312 VPWR.n1539 VPWR.t163 63.8431
R7313 VPWR.n1539 VPWR.t210 63.8431
R7314 VPWR.n1547 VPWR.t440 63.8431
R7315 VPWR.n1547 VPWR.t452 63.8431
R7316 VPWR.n1550 VPWR.t562 63.8431
R7317 VPWR.n1550 VPWR.t129 63.8431
R7318 VPWR.n1553 VPWR.t558 63.8431
R7319 VPWR.n1553 VPWR.t553 63.8431
R7320 VPWR.n1558 VPWR.t450 63.8431
R7321 VPWR.n1558 VPWR.t448 63.8431
R7322 VPWR.n1565 VPWR.t381 63.8431
R7323 VPWR.n1565 VPWR.t345 63.8431
R7324 VPWR.n1572 VPWR.t385 63.8431
R7325 VPWR.n1572 VPWR.t389 63.8431
R7326 VPWR.n1575 VPWR.t560 63.8431
R7327 VPWR.n1575 VPWR.t207 63.8431
R7328 VPWR.n1578 VPWR.t564 63.8431
R7329 VPWR.n1578 VPWR.t556 63.8431
R7330 VPWR.n1599 VPWR.t43 63.8431
R7331 VPWR.n1599 VPWR.t371 63.8431
R7332 VPWR.n1589 VPWR.t159 63.8431
R7333 VPWR.n1589 VPWR.t150 63.8431
R7334 VPWR.n1591 VPWR.t151 63.8431
R7335 VPWR.n1591 VPWR.t91 63.8431
R7336 VPWR.n1593 VPWR.t92 63.8431
R7337 VPWR.n1593 VPWR.t176 63.8431
R7338 VPWR.n1595 VPWR.t177 63.8431
R7339 VPWR.n1595 VPWR.t118 63.8431
R7340 VPWR.n1597 VPWR.t119 63.8431
R7341 VPWR.n1597 VPWR.t42 63.8431
R7342 VPWR.n759 VPWR.t580 63.8431
R7343 VPWR.n759 VPWR.t394 63.8431
R7344 VPWR.n733 VPWR.t218 63.8431
R7345 VPWR.n733 VPWR.t18 63.8431
R7346 VPWR.n658 VPWR.t362 63.8431
R7347 VPWR.n658 VPWR.t347 63.8431
R7348 VPWR.n663 VPWR.t351 63.8431
R7349 VPWR.n663 VPWR.t350 63.8431
R7350 VPWR.n668 VPWR.t506 63.8431
R7351 VPWR.n668 VPWR.t509 63.8431
R7352 VPWR.n673 VPWR.t426 63.8431
R7353 VPWR.n673 VPWR.t511 63.8431
R7354 VPWR.n701 VPWR.t598 63.8431
R7355 VPWR.n701 VPWR.t600 63.8431
R7356 VPWR.n706 VPWR.t583 63.8431
R7357 VPWR.n706 VPWR.t584 63.8431
R7358 VPWR.n711 VPWR.t405 63.8431
R7359 VPWR.n711 VPWR.t404 63.8431
R7360 VPWR.n716 VPWR.t374 63.8431
R7361 VPWR.n716 VPWR.t376 63.8431
R7362 VPWR.n232 VPWR.t471 63.8431
R7363 VPWR.n232 VPWR.t469 63.8431
R7364 VPWR.n237 VPWR.t411 63.8431
R7365 VPWR.n237 VPWR.t410 63.8431
R7366 VPWR.n242 VPWR.t491 63.8431
R7367 VPWR.n242 VPWR.t490 63.8431
R7368 VPWR.n247 VPWR.t219 63.8431
R7369 VPWR.n247 VPWR.t221 63.8431
R7370 VPWR.n200 VPWR.t454 63.8431
R7371 VPWR.n200 VPWR.t455 63.8431
R7372 VPWR.n205 VPWR.t360 63.8431
R7373 VPWR.n205 VPWR.t358 63.8431
R7374 VPWR.n210 VPWR.t516 63.8431
R7375 VPWR.n210 VPWR.t515 63.8431
R7376 VPWR.n215 VPWR.t494 63.8431
R7377 VPWR.n215 VPWR.t496 63.8431
R7378 VPWR.n1761 VPWR.t353 63.8431
R7379 VPWR.n1761 VPWR.t236 63.8431
R7380 VPWR.n305 VPWR.t512 63.8431
R7381 VPWR.n305 VPWR.t467 63.8431
R7382 VPWR.n429 VPWR.t547 63.8431
R7383 VPWR.n429 VPWR.t483 63.8431
R7384 VPWR.n403 VPWR.t484 63.8431
R7385 VPWR.n403 VPWR.t378 63.8431
R7386 VPWR.n347 VPWR.t421 63.8431
R7387 VPWR.n347 VPWR.t420 63.8431
R7388 VPWR.n352 VPWR.t418 63.8431
R7389 VPWR.n352 VPWR.t417 63.8431
R7390 VPWR.n357 VPWR.t573 63.8431
R7391 VPWR.n357 VPWR.t570 63.8431
R7392 VPWR.n362 VPWR.t398 63.8431
R7393 VPWR.n362 VPWR.t395 63.8431
R7394 VPWR.n1118 VPWR.t170 63.8431
R7395 VPWR.n1118 VPWR.t364 63.8431
R7396 VPWR.n1018 VPWR.t201 63.8431
R7397 VPWR.n1018 VPWR.t475 63.8431
R7398 VPWR.n2072 VPWR.n2071 60.9887
R7399 VPWR.n2137 VPWR.n2136 60.9887
R7400 VPWR.n2203 VPWR.n2202 60.9887
R7401 VPWR.n2269 VPWR.n2268 60.9887
R7402 VPWR.n1428 VPWR.n1248 60.9887
R7403 VPWR.n1435 VPWR.n1434 60.9887
R7404 VPWR.n1613 VPWR.n1612 60.9887
R7405 VPWR.n1724 VPWR.n1723 60.9887
R7406 VPWR.n954 VPWR.n953 60.9887
R7407 VPWR.n930 VPWR.n780 60.9887
R7408 VPWR.n1893 VPWR.n327 60.9887
R7409 VPWR.n1900 VPWR.n1899 60.9887
R7410 VPWR.n624 VPWR.n623 60.9887
R7411 VPWR.n600 VPWR.n450 60.9887
R7412 VPWR.n1166 VPWR.n1165 60.9887
R7413 VPWR.n1131 VPWR.n1130 60.9887
R7414 VPWR.n1103 VPWR.n1102 60.9887
R7415 VPWR.n2335 VPWR.n2334 60.9887
R7416 VPWR.n2022 VPWR.t289 58.0561
R7417 VPWR.n2023 VPWR.t331 58.0561
R7418 VPWR.t331 VPWR.n2017 58.0561
R7419 VPWR.t229 VPWR.n2030 58.0561
R7420 VPWR.n2031 VPWR.t229 58.0561
R7421 VPWR.t13 VPWR.n2031 58.0561
R7422 VPWR.n2033 VPWR.t13 58.0561
R7423 VPWR.n2032 VPWR.t594 58.0561
R7424 VPWR.n2040 VPWR.t594 58.0561
R7425 VPWR.t310 VPWR.n2041 58.0561
R7426 VPWR.n2043 VPWR.t310 58.0561
R7427 VPWR.n2042 VPWR.t228 58.0561
R7428 VPWR.n2049 VPWR.t228 58.0561
R7429 VPWR.t15 VPWR.n2049 58.0561
R7430 VPWR.n2050 VPWR.t15 58.0561
R7431 VPWR.n2052 VPWR.t0 58.0561
R7432 VPWR.t0 VPWR.n2051 58.0561
R7433 VPWR.n2051 VPWR.t550 58.0561
R7434 VPWR.n2059 VPWR.t550 58.0561
R7435 VPWR.t226 VPWR.n2060 58.0561
R7436 VPWR.n2062 VPWR.t226 58.0561
R7437 VPWR.n2061 VPWR.t19 58.0561
R7438 VPWR.n2068 VPWR.t19 58.0561
R7439 VPWR.t30 VPWR.n2069 58.0561
R7440 VPWR.n1720 VPWR.t98 58.0561
R7441 VPWR.n1719 VPWR.t2 58.0561
R7442 VPWR.t2 VPWR.n1718 58.0561
R7443 VPWR.t497 VPWR.n1457 58.0561
R7444 VPWR.n1712 VPWR.t497 58.0561
R7445 VPWR.n1712 VPWR.t596 58.0561
R7446 VPWR.t596 VPWR.n1711 58.0561
R7447 VPWR.n1710 VPWR.t4 58.0561
R7448 VPWR.n1464 VPWR.t4 58.0561
R7449 VPWR.t280 VPWR.n1464 58.0561
R7450 VPWR.n1704 VPWR.t280 58.0561
R7451 VPWR.n1703 VPWR.t372 58.0561
R7452 VPWR.t372 VPWR.n1702 58.0561
R7453 VPWR.t79 VPWR.n1465 58.0561
R7454 VPWR.n1696 VPWR.t79 58.0561
R7455 VPWR.n1696 VPWR.t52 58.0561
R7456 VPWR.t52 VPWR.n1695 58.0561
R7457 VPWR.n1695 VPWR.t64 58.0561
R7458 VPWR.t64 VPWR.n1694 58.0561
R7459 VPWR.n1694 VPWR.t110 58.0561
R7460 VPWR.n1471 VPWR.t110 58.0561
R7461 VPWR.t161 VPWR.n1471 58.0561
R7462 VPWR.n1688 VPWR.t161 58.0561
R7463 VPWR.n1688 VPWR.t209 58.0561
R7464 VPWR.t209 VPWR.n1687 58.0561
R7465 VPWR.n1687 VPWR.t368 58.0561
R7466 VPWR.t368 VPWR.n1686 58.0561
R7467 VPWR.t441 VPWR.n1472 58.0561
R7468 VPWR.n1680 VPWR.t441 58.0561
R7469 VPWR.n1680 VPWR.t439 58.0561
R7470 VPWR.t439 VPWR.n1679 58.0561
R7471 VPWR.n1679 VPWR.t451 58.0561
R7472 VPWR.t451 VPWR.n1678 58.0561
R7473 VPWR.n1678 VPWR.t561 58.0561
R7474 VPWR.n1479 VPWR.t561 58.0561
R7475 VPWR.t128 VPWR.n1479 58.0561
R7476 VPWR.n1672 VPWR.t128 58.0561
R7477 VPWR.n1672 VPWR.t557 58.0561
R7478 VPWR.t557 VPWR.n1671 58.0561
R7479 VPWR.n1671 VPWR.t552 58.0561
R7480 VPWR.t552 VPWR.n1670 58.0561
R7481 VPWR.t445 VPWR.n1480 58.0561
R7482 VPWR.n1664 VPWR.t445 58.0561
R7483 VPWR.n1664 VPWR.t449 58.0561
R7484 VPWR.t449 VPWR.n1663 58.0561
R7485 VPWR.n1663 VPWR.t447 58.0561
R7486 VPWR.t447 VPWR.n1662 58.0561
R7487 VPWR.n1662 VPWR.t443 58.0561
R7488 VPWR.n1487 VPWR.t443 58.0561
R7489 VPWR.n1656 VPWR.t386 58.0561
R7490 VPWR.t386 VPWR.n1655 58.0561
R7491 VPWR.n1655 VPWR.t380 58.0561
R7492 VPWR.t380 VPWR.n1654 58.0561
R7493 VPWR.n1654 VPWR.t344 58.0561
R7494 VPWR.n1492 VPWR.t344 58.0561
R7495 VPWR.t390 VPWR.n1492 58.0561
R7496 VPWR.n1648 VPWR.t390 58.0561
R7497 VPWR.n1647 VPWR.t382 58.0561
R7498 VPWR.t382 VPWR.n1646 58.0561
R7499 VPWR.n1646 VPWR.t384 58.0561
R7500 VPWR.n1495 VPWR.t384 58.0561
R7501 VPWR.t388 VPWR.n1495 58.0561
R7502 VPWR.n1640 VPWR.t388 58.0561
R7503 VPWR.n1640 VPWR.t559 58.0561
R7504 VPWR.t559 VPWR.n1639 58.0561
R7505 VPWR.n1639 VPWR.t206 58.0561
R7506 VPWR.t206 VPWR.n1638 58.0561
R7507 VPWR.n1638 VPWR.t563 58.0561
R7508 VPWR.n1500 VPWR.t563 58.0561
R7509 VPWR.t555 VPWR.n1500 58.0561
R7510 VPWR.n1632 VPWR.t555 58.0561
R7511 VPWR.n1631 VPWR.t157 58.0561
R7512 VPWR.t157 VPWR.n1630 58.0561
R7513 VPWR.n1630 VPWR.t149 58.0561
R7514 VPWR.n1503 VPWR.t149 58.0561
R7515 VPWR.t90 VPWR.n1503 58.0561
R7516 VPWR.n1624 VPWR.t90 58.0561
R7517 VPWR.n1624 VPWR.t175 58.0561
R7518 VPWR.t175 VPWR.n1623 58.0561
R7519 VPWR.n1623 VPWR.t117 58.0561
R7520 VPWR.t117 VPWR.n1622 58.0561
R7521 VPWR.n1622 VPWR.t41 58.0561
R7522 VPWR.n1508 VPWR.t41 58.0561
R7523 VPWR.t370 VPWR.n1508 58.0561
R7524 VPWR.n1616 VPWR.t370 58.0561
R7525 VPWR.n1615 VPWR.t186 58.0561
R7526 VPWR.n1936 VPWR.t86 58.0561
R7527 VPWR.n1935 VPWR.t329 58.0561
R7528 VPWR.t329 VPWR.n1934 58.0561
R7529 VPWR.t234 VPWR.n1922 58.0561
R7530 VPWR.n1928 VPWR.t234 58.0561
R7531 VPWR.n1927 VPWR.t500 58.0561
R7532 VPWR.n1099 VPWR.t137 58.0561
R7533 VPWR.n1098 VPWR.t246 58.0561
R7534 VPWR.t246 VPWR.n1085 58.0561
R7535 VPWR.t121 VPWR.n1134 58.0561
R7536 VPWR.n1135 VPWR.t121 58.0561
R7537 VPWR.n1136 VPWR.t301 58.0561
R7538 VPWR.t301 VPWR.n1081 58.0561
R7539 VPWR.t323 VPWR.n1143 58.0561
R7540 VPWR.n1144 VPWR.t323 58.0561
R7541 VPWR.t365 VPWR.n1144 58.0561
R7542 VPWR.n1146 VPWR.t365 58.0561
R7543 VPWR.n1145 VPWR.t366 58.0561
R7544 VPWR.n1153 VPWR.t366 58.0561
R7545 VPWR.t169 VPWR.n1153 58.0561
R7546 VPWR.n1154 VPWR.t169 58.0561
R7547 VPWR.t363 VPWR.n1154 58.0561
R7548 VPWR.n1156 VPWR.t363 58.0561
R7549 VPWR.n1155 VPWR.t427 58.0561
R7550 VPWR.n1162 VPWR.t427 58.0561
R7551 VPWR.t141 VPWR.n1163 58.0561
R7552 VPWR.n1003 VPWR.t45 58.0561
R7553 VPWR.n1002 VPWR.t335 58.0561
R7554 VPWR.t335 VPWR.n995 58.0561
R7555 VPWR.t37 VPWR.n1032 58.0561
R7556 VPWR.n1033 VPWR.t37 58.0561
R7557 VPWR.n1034 VPWR.t241 58.0561
R7558 VPWR.t241 VPWR.n991 58.0561
R7559 VPWR.t254 VPWR.n1041 58.0561
R7560 VPWR.n1042 VPWR.t254 58.0561
R7561 VPWR.t473 VPWR.n1042 58.0561
R7562 VPWR.n1044 VPWR.t473 58.0561
R7563 VPWR.n1043 VPWR.t472 58.0561
R7564 VPWR.n1051 VPWR.t472 58.0561
R7565 VPWR.t200 VPWR.n1051 58.0561
R7566 VPWR.n1052 VPWR.t200 58.0561
R7567 VPWR.t474 VPWR.n1052 58.0561
R7568 VPWR.n1054 VPWR.t474 58.0561
R7569 VPWR.n1053 VPWR.t429 58.0561
R7570 VPWR.n1060 VPWR.t429 58.0561
R7571 VPWR.t179 VPWR.n1061 58.0561
R7572 VPWR.n1949 VPWR 46.7832
R7573 VPWR.n1954 VPWR 46.7832
R7574 VPWR.n1959 VPWR 46.7832
R7575 VPWR.n2082 VPWR.n2081 43.2946
R7576 VPWR.n2148 VPWR.n2147 43.2946
R7577 VPWR.n2214 VPWR.n2213 43.2946
R7578 VPWR.n1279 VPWR.n1277 43.2946
R7579 VPWR.n1314 VPWR.n1313 43.2946
R7580 VPWR.n932 VPWR.n931 43.2946
R7581 VPWR.n952 VPWR.n951 43.2946
R7582 VPWR.n1744 VPWR.n1742 43.2946
R7583 VPWR.n1779 VPWR.n1778 43.2946
R7584 VPWR.n602 VPWR.n601 43.2946
R7585 VPWR.n622 VPWR.n621 43.2946
R7586 VPWR.n1028 VPWR.n1027 43.2946
R7587 VPWR.n1065 VPWR.n1064 43.2946
R7588 VPWR.n1008 VPWR.n1007 43.2946
R7589 VPWR.n2280 VPWR.n2279 43.2946
R7590 VPWR.n2136 VPWR 40.6593
R7591 VPWR.n2202 VPWR 40.6593
R7592 VPWR.n2268 VPWR 40.6593
R7593 VPWR.n1434 VPWR 40.6593
R7594 VPWR.n1428 VPWR 40.6593
R7595 VPWR VPWR.n930 40.6593
R7596 VPWR.n953 VPWR 40.6593
R7597 VPWR.n1899 VPWR 40.6593
R7598 VPWR.n1893 VPWR 40.6593
R7599 VPWR VPWR.n600 40.6593
R7600 VPWR.n623 VPWR 40.6593
R7601 VPWR.n1029 VPWR 40.6593
R7602 VPWR VPWR.n1063 40.6593
R7603 VPWR VPWR.n1006 40.6593
R7604 VPWR.n2334 VPWR 40.6593
R7605 VPWR.n1918 VPWR 39.2538
R7606 VPWR.n1942 VPWR 39.2538
R7607 VPWR.n2095 VPWR.n2085 38.6708
R7608 VPWR.n2129 VPWR.n2086 38.6708
R7609 VPWR.n2125 VPWR.n2087 38.6708
R7610 VPWR.n2121 VPWR.n2088 38.6708
R7611 VPWR.n2117 VPWR.n2089 38.6708
R7612 VPWR.n2113 VPWR.n2090 38.6708
R7613 VPWR.n2109 VPWR.n2091 38.6708
R7614 VPWR.n2105 VPWR.n2092 38.6708
R7615 VPWR.n2101 VPWR.n2093 38.6708
R7616 VPWR.n2097 VPWR.n2094 38.6708
R7617 VPWR.n2130 VPWR.n2085 38.6708
R7618 VPWR.n2126 VPWR.n2086 38.6708
R7619 VPWR.n2122 VPWR.n2087 38.6708
R7620 VPWR.n2118 VPWR.n2088 38.6708
R7621 VPWR.n2114 VPWR.n2089 38.6708
R7622 VPWR.n2110 VPWR.n2090 38.6708
R7623 VPWR.n2106 VPWR.n2091 38.6708
R7624 VPWR.n2102 VPWR.n2092 38.6708
R7625 VPWR.n2098 VPWR.n2093 38.6708
R7626 VPWR.n2094 VPWR.n2084 38.6708
R7627 VPWR.n2161 VPWR.n2151 38.6708
R7628 VPWR.n2195 VPWR.n2152 38.6708
R7629 VPWR.n2191 VPWR.n2153 38.6708
R7630 VPWR.n2187 VPWR.n2154 38.6708
R7631 VPWR.n2183 VPWR.n2155 38.6708
R7632 VPWR.n2179 VPWR.n2156 38.6708
R7633 VPWR.n2175 VPWR.n2157 38.6708
R7634 VPWR.n2171 VPWR.n2158 38.6708
R7635 VPWR.n2167 VPWR.n2159 38.6708
R7636 VPWR.n2163 VPWR.n2160 38.6708
R7637 VPWR.n2196 VPWR.n2151 38.6708
R7638 VPWR.n2192 VPWR.n2152 38.6708
R7639 VPWR.n2188 VPWR.n2153 38.6708
R7640 VPWR.n2184 VPWR.n2154 38.6708
R7641 VPWR.n2180 VPWR.n2155 38.6708
R7642 VPWR.n2176 VPWR.n2156 38.6708
R7643 VPWR.n2172 VPWR.n2157 38.6708
R7644 VPWR.n2168 VPWR.n2158 38.6708
R7645 VPWR.n2164 VPWR.n2159 38.6708
R7646 VPWR.n2160 VPWR.n2150 38.6708
R7647 VPWR.n2227 VPWR.n2217 38.6708
R7648 VPWR.n2261 VPWR.n2218 38.6708
R7649 VPWR.n2257 VPWR.n2219 38.6708
R7650 VPWR.n2253 VPWR.n2220 38.6708
R7651 VPWR.n2249 VPWR.n2221 38.6708
R7652 VPWR.n2245 VPWR.n2222 38.6708
R7653 VPWR.n2241 VPWR.n2223 38.6708
R7654 VPWR.n2237 VPWR.n2224 38.6708
R7655 VPWR.n2233 VPWR.n2225 38.6708
R7656 VPWR.n2229 VPWR.n2226 38.6708
R7657 VPWR.n2262 VPWR.n2217 38.6708
R7658 VPWR.n2258 VPWR.n2218 38.6708
R7659 VPWR.n2254 VPWR.n2219 38.6708
R7660 VPWR.n2250 VPWR.n2220 38.6708
R7661 VPWR.n2246 VPWR.n2221 38.6708
R7662 VPWR.n2242 VPWR.n2222 38.6708
R7663 VPWR.n2238 VPWR.n2223 38.6708
R7664 VPWR.n2234 VPWR.n2224 38.6708
R7665 VPWR.n2230 VPWR.n2225 38.6708
R7666 VPWR.n2226 VPWR.n2216 38.6708
R7667 VPWR.n1432 VPWR.n1431 38.6708
R7668 VPWR.n1315 VPWR.n1181 38.6708
R7669 VPWR.n1319 VPWR.n1182 38.6708
R7670 VPWR.n1323 VPWR.n1183 38.6708
R7671 VPWR.n1327 VPWR.n1184 38.6708
R7672 VPWR.n1331 VPWR.n1185 38.6708
R7673 VPWR.n1335 VPWR.n1186 38.6708
R7674 VPWR.n1339 VPWR.n1187 38.6708
R7675 VPWR.n1343 VPWR.n1188 38.6708
R7676 VPWR.n1347 VPWR.n1189 38.6708
R7677 VPWR.n1351 VPWR.n1190 38.6708
R7678 VPWR.n1355 VPWR.n1191 38.6708
R7679 VPWR.n1359 VPWR.n1192 38.6708
R7680 VPWR.n1363 VPWR.n1193 38.6708
R7681 VPWR.n1367 VPWR.n1194 38.6708
R7682 VPWR.n1371 VPWR.n1195 38.6708
R7683 VPWR.n1375 VPWR.n1196 38.6708
R7684 VPWR.n1379 VPWR.n1197 38.6708
R7685 VPWR.n1383 VPWR.n1198 38.6708
R7686 VPWR.n1387 VPWR.n1199 38.6708
R7687 VPWR.n1391 VPWR.n1200 38.6708
R7688 VPWR.n1395 VPWR.n1201 38.6708
R7689 VPWR.n1399 VPWR.n1202 38.6708
R7690 VPWR.n1403 VPWR.n1203 38.6708
R7691 VPWR.n1407 VPWR.n1204 38.6708
R7692 VPWR.n1411 VPWR.n1205 38.6708
R7693 VPWR.n1415 VPWR.n1206 38.6708
R7694 VPWR.n1419 VPWR.n1207 38.6708
R7695 VPWR.n1423 VPWR.n1208 38.6708
R7696 VPWR.n1429 VPWR.n1209 38.6708
R7697 VPWR.n1431 VPWR.n1180 38.6708
R7698 VPWR.n1318 VPWR.n1181 38.6708
R7699 VPWR.n1322 VPWR.n1182 38.6708
R7700 VPWR.n1326 VPWR.n1183 38.6708
R7701 VPWR.n1330 VPWR.n1184 38.6708
R7702 VPWR.n1334 VPWR.n1185 38.6708
R7703 VPWR.n1338 VPWR.n1186 38.6708
R7704 VPWR.n1342 VPWR.n1187 38.6708
R7705 VPWR.n1346 VPWR.n1188 38.6708
R7706 VPWR.n1350 VPWR.n1189 38.6708
R7707 VPWR.n1354 VPWR.n1190 38.6708
R7708 VPWR.n1358 VPWR.n1191 38.6708
R7709 VPWR.n1362 VPWR.n1192 38.6708
R7710 VPWR.n1366 VPWR.n1193 38.6708
R7711 VPWR.n1370 VPWR.n1194 38.6708
R7712 VPWR.n1374 VPWR.n1195 38.6708
R7713 VPWR.n1378 VPWR.n1196 38.6708
R7714 VPWR.n1382 VPWR.n1197 38.6708
R7715 VPWR.n1386 VPWR.n1198 38.6708
R7716 VPWR.n1390 VPWR.n1199 38.6708
R7717 VPWR.n1394 VPWR.n1200 38.6708
R7718 VPWR.n1398 VPWR.n1201 38.6708
R7719 VPWR.n1402 VPWR.n1202 38.6708
R7720 VPWR.n1406 VPWR.n1203 38.6708
R7721 VPWR.n1410 VPWR.n1204 38.6708
R7722 VPWR.n1414 VPWR.n1205 38.6708
R7723 VPWR.n1418 VPWR.n1206 38.6708
R7724 VPWR.n1422 VPWR.n1207 38.6708
R7725 VPWR.n1425 VPWR.n1208 38.6708
R7726 VPWR.n812 VPWR.n783 38.6708
R7727 VPWR.n816 VPWR.n784 38.6708
R7728 VPWR.n820 VPWR.n785 38.6708
R7729 VPWR.n824 VPWR.n786 38.6708
R7730 VPWR.n828 VPWR.n787 38.6708
R7731 VPWR.n832 VPWR.n788 38.6708
R7732 VPWR.n836 VPWR.n789 38.6708
R7733 VPWR.n840 VPWR.n790 38.6708
R7734 VPWR.n844 VPWR.n791 38.6708
R7735 VPWR.n848 VPWR.n792 38.6708
R7736 VPWR.n852 VPWR.n793 38.6708
R7737 VPWR.n856 VPWR.n794 38.6708
R7738 VPWR.n860 VPWR.n795 38.6708
R7739 VPWR.n864 VPWR.n796 38.6708
R7740 VPWR.n868 VPWR.n797 38.6708
R7741 VPWR.n872 VPWR.n798 38.6708
R7742 VPWR.n876 VPWR.n799 38.6708
R7743 VPWR.n880 VPWR.n800 38.6708
R7744 VPWR.n884 VPWR.n801 38.6708
R7745 VPWR.n888 VPWR.n802 38.6708
R7746 VPWR.n892 VPWR.n803 38.6708
R7747 VPWR.n896 VPWR.n804 38.6708
R7748 VPWR.n900 VPWR.n805 38.6708
R7749 VPWR.n904 VPWR.n806 38.6708
R7750 VPWR.n908 VPWR.n807 38.6708
R7751 VPWR.n912 VPWR.n808 38.6708
R7752 VPWR.n916 VPWR.n809 38.6708
R7753 VPWR.n920 VPWR.n810 38.6708
R7754 VPWR.n927 VPWR.n811 38.6708
R7755 VPWR.n929 VPWR.n782 38.6708
R7756 VPWR.n815 VPWR.n783 38.6708
R7757 VPWR.n819 VPWR.n784 38.6708
R7758 VPWR.n823 VPWR.n785 38.6708
R7759 VPWR.n827 VPWR.n786 38.6708
R7760 VPWR.n831 VPWR.n787 38.6708
R7761 VPWR.n835 VPWR.n788 38.6708
R7762 VPWR.n839 VPWR.n789 38.6708
R7763 VPWR.n843 VPWR.n790 38.6708
R7764 VPWR.n847 VPWR.n791 38.6708
R7765 VPWR.n851 VPWR.n792 38.6708
R7766 VPWR.n855 VPWR.n793 38.6708
R7767 VPWR.n859 VPWR.n794 38.6708
R7768 VPWR.n863 VPWR.n795 38.6708
R7769 VPWR.n867 VPWR.n796 38.6708
R7770 VPWR.n871 VPWR.n797 38.6708
R7771 VPWR.n875 VPWR.n798 38.6708
R7772 VPWR.n879 VPWR.n799 38.6708
R7773 VPWR.n883 VPWR.n800 38.6708
R7774 VPWR.n887 VPWR.n801 38.6708
R7775 VPWR.n891 VPWR.n802 38.6708
R7776 VPWR.n895 VPWR.n803 38.6708
R7777 VPWR.n899 VPWR.n804 38.6708
R7778 VPWR.n903 VPWR.n805 38.6708
R7779 VPWR.n907 VPWR.n806 38.6708
R7780 VPWR.n911 VPWR.n807 38.6708
R7781 VPWR.n915 VPWR.n808 38.6708
R7782 VPWR.n919 VPWR.n809 38.6708
R7783 VPWR.n922 VPWR.n810 38.6708
R7784 VPWR.n927 VPWR.n926 38.6708
R7785 VPWR.n1897 VPWR.n1896 38.6708
R7786 VPWR.n1780 VPWR.n260 38.6708
R7787 VPWR.n1784 VPWR.n261 38.6708
R7788 VPWR.n1788 VPWR.n262 38.6708
R7789 VPWR.n1792 VPWR.n263 38.6708
R7790 VPWR.n1796 VPWR.n264 38.6708
R7791 VPWR.n1800 VPWR.n265 38.6708
R7792 VPWR.n1804 VPWR.n266 38.6708
R7793 VPWR.n1808 VPWR.n267 38.6708
R7794 VPWR.n1812 VPWR.n268 38.6708
R7795 VPWR.n1816 VPWR.n269 38.6708
R7796 VPWR.n1820 VPWR.n270 38.6708
R7797 VPWR.n1824 VPWR.n271 38.6708
R7798 VPWR.n1828 VPWR.n272 38.6708
R7799 VPWR.n1832 VPWR.n273 38.6708
R7800 VPWR.n1836 VPWR.n274 38.6708
R7801 VPWR.n1840 VPWR.n275 38.6708
R7802 VPWR.n1844 VPWR.n276 38.6708
R7803 VPWR.n1848 VPWR.n277 38.6708
R7804 VPWR.n1852 VPWR.n278 38.6708
R7805 VPWR.n1856 VPWR.n279 38.6708
R7806 VPWR.n1860 VPWR.n280 38.6708
R7807 VPWR.n1864 VPWR.n281 38.6708
R7808 VPWR.n1868 VPWR.n282 38.6708
R7809 VPWR.n1872 VPWR.n283 38.6708
R7810 VPWR.n1876 VPWR.n284 38.6708
R7811 VPWR.n1880 VPWR.n285 38.6708
R7812 VPWR.n1884 VPWR.n286 38.6708
R7813 VPWR.n1888 VPWR.n287 38.6708
R7814 VPWR.n1894 VPWR.n288 38.6708
R7815 VPWR.n1896 VPWR.n259 38.6708
R7816 VPWR.n1783 VPWR.n260 38.6708
R7817 VPWR.n1787 VPWR.n261 38.6708
R7818 VPWR.n1791 VPWR.n262 38.6708
R7819 VPWR.n1795 VPWR.n263 38.6708
R7820 VPWR.n1799 VPWR.n264 38.6708
R7821 VPWR.n1803 VPWR.n265 38.6708
R7822 VPWR.n1807 VPWR.n266 38.6708
R7823 VPWR.n1811 VPWR.n267 38.6708
R7824 VPWR.n1815 VPWR.n268 38.6708
R7825 VPWR.n1819 VPWR.n269 38.6708
R7826 VPWR.n1823 VPWR.n270 38.6708
R7827 VPWR.n1827 VPWR.n271 38.6708
R7828 VPWR.n1831 VPWR.n272 38.6708
R7829 VPWR.n1835 VPWR.n273 38.6708
R7830 VPWR.n1839 VPWR.n274 38.6708
R7831 VPWR.n1843 VPWR.n275 38.6708
R7832 VPWR.n1847 VPWR.n276 38.6708
R7833 VPWR.n1851 VPWR.n277 38.6708
R7834 VPWR.n1855 VPWR.n278 38.6708
R7835 VPWR.n1859 VPWR.n279 38.6708
R7836 VPWR.n1863 VPWR.n280 38.6708
R7837 VPWR.n1867 VPWR.n281 38.6708
R7838 VPWR.n1871 VPWR.n282 38.6708
R7839 VPWR.n1875 VPWR.n283 38.6708
R7840 VPWR.n1879 VPWR.n284 38.6708
R7841 VPWR.n1883 VPWR.n285 38.6708
R7842 VPWR.n1887 VPWR.n286 38.6708
R7843 VPWR.n1890 VPWR.n287 38.6708
R7844 VPWR.n482 VPWR.n453 38.6708
R7845 VPWR.n486 VPWR.n454 38.6708
R7846 VPWR.n490 VPWR.n455 38.6708
R7847 VPWR.n494 VPWR.n456 38.6708
R7848 VPWR.n498 VPWR.n457 38.6708
R7849 VPWR.n502 VPWR.n458 38.6708
R7850 VPWR.n506 VPWR.n459 38.6708
R7851 VPWR.n510 VPWR.n460 38.6708
R7852 VPWR.n514 VPWR.n461 38.6708
R7853 VPWR.n518 VPWR.n462 38.6708
R7854 VPWR.n522 VPWR.n463 38.6708
R7855 VPWR.n526 VPWR.n464 38.6708
R7856 VPWR.n530 VPWR.n465 38.6708
R7857 VPWR.n534 VPWR.n466 38.6708
R7858 VPWR.n538 VPWR.n467 38.6708
R7859 VPWR.n542 VPWR.n468 38.6708
R7860 VPWR.n546 VPWR.n469 38.6708
R7861 VPWR.n550 VPWR.n470 38.6708
R7862 VPWR.n554 VPWR.n471 38.6708
R7863 VPWR.n558 VPWR.n472 38.6708
R7864 VPWR.n562 VPWR.n473 38.6708
R7865 VPWR.n566 VPWR.n474 38.6708
R7866 VPWR.n570 VPWR.n475 38.6708
R7867 VPWR.n574 VPWR.n476 38.6708
R7868 VPWR.n578 VPWR.n477 38.6708
R7869 VPWR.n582 VPWR.n478 38.6708
R7870 VPWR.n586 VPWR.n479 38.6708
R7871 VPWR.n590 VPWR.n480 38.6708
R7872 VPWR.n597 VPWR.n481 38.6708
R7873 VPWR.n599 VPWR.n452 38.6708
R7874 VPWR.n485 VPWR.n453 38.6708
R7875 VPWR.n489 VPWR.n454 38.6708
R7876 VPWR.n493 VPWR.n455 38.6708
R7877 VPWR.n497 VPWR.n456 38.6708
R7878 VPWR.n501 VPWR.n457 38.6708
R7879 VPWR.n505 VPWR.n458 38.6708
R7880 VPWR.n509 VPWR.n459 38.6708
R7881 VPWR.n513 VPWR.n460 38.6708
R7882 VPWR.n517 VPWR.n461 38.6708
R7883 VPWR.n521 VPWR.n462 38.6708
R7884 VPWR.n525 VPWR.n463 38.6708
R7885 VPWR.n529 VPWR.n464 38.6708
R7886 VPWR.n533 VPWR.n465 38.6708
R7887 VPWR.n537 VPWR.n466 38.6708
R7888 VPWR.n541 VPWR.n467 38.6708
R7889 VPWR.n545 VPWR.n468 38.6708
R7890 VPWR.n549 VPWR.n469 38.6708
R7891 VPWR.n553 VPWR.n470 38.6708
R7892 VPWR.n557 VPWR.n471 38.6708
R7893 VPWR.n561 VPWR.n472 38.6708
R7894 VPWR.n565 VPWR.n473 38.6708
R7895 VPWR.n569 VPWR.n474 38.6708
R7896 VPWR.n573 VPWR.n475 38.6708
R7897 VPWR.n577 VPWR.n476 38.6708
R7898 VPWR.n581 VPWR.n477 38.6708
R7899 VPWR.n585 VPWR.n478 38.6708
R7900 VPWR.n589 VPWR.n479 38.6708
R7901 VPWR.n592 VPWR.n480 38.6708
R7902 VPWR.n597 VPWR.n596 38.6708
R7903 VPWR.n2293 VPWR.n2283 38.6708
R7904 VPWR.n2327 VPWR.n2284 38.6708
R7905 VPWR.n2323 VPWR.n2285 38.6708
R7906 VPWR.n2319 VPWR.n2286 38.6708
R7907 VPWR.n2315 VPWR.n2287 38.6708
R7908 VPWR.n2311 VPWR.n2288 38.6708
R7909 VPWR.n2307 VPWR.n2289 38.6708
R7910 VPWR.n2303 VPWR.n2290 38.6708
R7911 VPWR.n2299 VPWR.n2291 38.6708
R7912 VPWR.n2295 VPWR.n2292 38.6708
R7913 VPWR.n2328 VPWR.n2283 38.6708
R7914 VPWR.n2324 VPWR.n2284 38.6708
R7915 VPWR.n2320 VPWR.n2285 38.6708
R7916 VPWR.n2316 VPWR.n2286 38.6708
R7917 VPWR.n2312 VPWR.n2287 38.6708
R7918 VPWR.n2308 VPWR.n2288 38.6708
R7919 VPWR.n2304 VPWR.n2289 38.6708
R7920 VPWR.n2300 VPWR.n2290 38.6708
R7921 VPWR.n2296 VPWR.n2291 38.6708
R7922 VPWR.n2292 VPWR.n2282 38.6708
R7923 VPWR.n2210 VPWR.n114 38.3102
R7924 VPWR.n638 VPWR.n114 37.1032
R7925 VPWR.n2342 VPWR.n28 37.1032
R7926 VPWR.n2078 VPWR.n1979 36.2684
R7927 VPWR.n2144 VPWR.n154 36.2684
R7928 VPWR.n2276 VPWR.n74 36.2684
R7929 VPWR.n2342 VPWR.n2341 35.5276
R7930 VPWR.n1978 VPWR.n195 35.0614
R7931 VPWR.n691 VPWR.n690 35.0614
R7932 VPWR.n2073 VPWR.n2005 35.0123
R7933 VPWR.n2075 VPWR.n2073 35.0123
R7934 VPWR.n2138 VPWR.n176 35.0123
R7935 VPWR.n2140 VPWR.n2138 35.0123
R7936 VPWR.n2204 VPWR.n136 35.0123
R7937 VPWR.n2206 VPWR.n2204 35.0123
R7938 VPWR.n2270 VPWR.n96 35.0123
R7939 VPWR.n2272 VPWR.n2270 35.0123
R7940 VPWR.n1442 VPWR.n1440 35.0123
R7941 VPWR.n1247 VPWR.n1246 35.0123
R7942 VPWR.n1247 VPWR.n1210 35.0123
R7943 VPWR.n1440 VPWR.n1439 35.0123
R7944 VPWR.n1731 VPWR.n1729 35.0123
R7945 VPWR.n1611 VPWR.n1610 35.0123
R7946 VPWR.n1611 VPWR.n1509 35.0123
R7947 VPWR.n1729 VPWR.n1728 35.0123
R7948 VPWR.n779 VPWR.n778 35.0123
R7949 VPWR.n961 VPWR.n959 35.0123
R7950 VPWR.n959 VPWR.n958 35.0123
R7951 VPWR.n779 VPWR.n742 35.0123
R7952 VPWR.n1907 VPWR.n1905 35.0123
R7953 VPWR.n326 VPWR.n325 35.0123
R7954 VPWR.n326 VPWR.n289 35.0123
R7955 VPWR.n1905 VPWR.n1904 35.0123
R7956 VPWR.n449 VPWR.n448 35.0123
R7957 VPWR.n631 VPWR.n629 35.0123
R7958 VPWR.n629 VPWR.n628 35.0123
R7959 VPWR.n449 VPWR.n412 35.0123
R7960 VPWR.n1104 VPWR.n1094 35.0123
R7961 VPWR.n1169 VPWR.n1167 35.0123
R7962 VPWR.n1167 VPWR.n1074 35.0123
R7963 VPWR.n1129 VPWR.n1128 35.0123
R7964 VPWR.n1129 VPWR.n1088 35.0123
R7965 VPWR.n1106 VPWR.n1104 35.0123
R7966 VPWR.n2336 VPWR.n49 35.0123
R7967 VPWR.n2338 VPWR.n2336 35.0123
R7968 VPWR.n2143 VPWR.n155 33.4858
R7969 VPWR.n2209 VPWR.n115 33.4858
R7970 VPWR.n2275 VPWR.n75 33.4858
R7971 VPWR.n1941 VPWR.n1918 32.0005
R7972 VPWR.n1942 VPWR.n1941 32.0005
R7973 VPWR.n1941 VPWR 26.8805
R7974 VPWR VPWR.n1940 23.0405
R7975 VPWR.n2073 VPWR 22.9652
R7976 VPWR.n2138 VPWR 22.9652
R7977 VPWR.n2204 VPWR 22.9652
R7978 VPWR.n2270 VPWR 22.9652
R7979 VPWR VPWR.n1247 22.9652
R7980 VPWR.n1440 VPWR 22.9652
R7981 VPWR VPWR.n1611 22.9652
R7982 VPWR.n1729 VPWR 22.9652
R7983 VPWR.n959 VPWR 22.9652
R7984 VPWR VPWR.n779 22.9652
R7985 VPWR VPWR.n326 22.9652
R7986 VPWR.n1905 VPWR 22.9652
R7987 VPWR.n629 VPWR 22.9652
R7988 VPWR VPWR.n449 22.9652
R7989 VPWR.n1167 VPWR 22.9652
R7990 VPWR VPWR.n1129 22.9652
R7991 VPWR.n1104 VPWR 22.9652
R7992 VPWR.n2336 VPWR 22.9652
R7993 VPWR.n2081 VPWR 21.4593
R7994 VPWR.n2081 VPWR 21.4593
R7995 VPWR.n2147 VPWR 21.4593
R7996 VPWR.n2147 VPWR 21.4593
R7997 VPWR.n2213 VPWR 21.4593
R7998 VPWR.n2213 VPWR 21.4593
R7999 VPWR.n1313 VPWR 21.4593
R8000 VPWR VPWR.n1279 21.4593
R8001 VPWR.n1279 VPWR 21.4593
R8002 VPWR.n1313 VPWR 21.4593
R8003 VPWR.n951 VPWR 21.4593
R8004 VPWR.n932 VPWR 21.4593
R8005 VPWR VPWR.n932 21.4593
R8006 VPWR.n951 VPWR 21.4593
R8007 VPWR.n1778 VPWR 21.4593
R8008 VPWR VPWR.n1744 21.4593
R8009 VPWR.n1744 VPWR 21.4593
R8010 VPWR.n1778 VPWR 21.4593
R8011 VPWR.n621 VPWR 21.4593
R8012 VPWR.n602 VPWR 21.4593
R8013 VPWR VPWR.n602 21.4593
R8014 VPWR.n621 VPWR 21.4593
R8015 VPWR VPWR.n1008 21.4593
R8016 VPWR.n1027 VPWR 21.4593
R8017 VPWR.n1027 VPWR 21.4593
R8018 VPWR VPWR.n1065 21.4593
R8019 VPWR.n1065 VPWR 21.4593
R8020 VPWR.n1008 VPWR 21.4593
R8021 VPWR.n2279 VPWR 21.4593
R8022 VPWR.n2279 VPWR 21.4593
R8023 VPWR VPWR.n2072 20.3299
R8024 VPWR VPWR.n2082 20.3299
R8025 VPWR VPWR.n2137 20.3299
R8026 VPWR VPWR.n2148 20.3299
R8027 VPWR VPWR.n2203 20.3299
R8028 VPWR VPWR.n2214 20.3299
R8029 VPWR VPWR.n2269 20.3299
R8030 VPWR.n1277 VPWR 20.3299
R8031 VPWR.n1248 VPWR 20.3299
R8032 VPWR VPWR.n1314 20.3299
R8033 VPWR VPWR.n1435 20.3299
R8034 VPWR.n1612 VPWR 20.3299
R8035 VPWR VPWR.n1724 20.3299
R8036 VPWR.n1523 VPWR 20.3299
R8037 VPWR.n1524 VPWR.n1523 20.3299
R8038 VPWR.n1524 VPWR 20.3299
R8039 VPWR.n1525 VPWR.n1524 20.3299
R8040 VPWR.n1525 VPWR 20.3299
R8041 VPWR.n1526 VPWR.n1525 20.3299
R8042 VPWR.n1526 VPWR 20.3299
R8043 VPWR.n1527 VPWR.n1526 20.3299
R8044 VPWR.n1527 VPWR 20.3299
R8045 VPWR.n1528 VPWR.n1527 20.3299
R8046 VPWR VPWR.n1528 20.3299
R8047 VPWR.n1530 VPWR 20.3299
R8048 VPWR.n1529 VPWR 20.3299
R8049 VPWR.n1532 VPWR.n1530 20.3299
R8050 VPWR.n1532 VPWR 20.3299
R8051 VPWR.n1534 VPWR.n1532 20.3299
R8052 VPWR.n1534 VPWR 20.3299
R8053 VPWR.n1536 VPWR.n1534 20.3299
R8054 VPWR.n1536 VPWR 20.3299
R8055 VPWR.n1538 VPWR.n1536 20.3299
R8056 VPWR.n1538 VPWR 20.3299
R8057 VPWR.n1540 VPWR.n1538 20.3299
R8058 VPWR.n1540 VPWR 20.3299
R8059 VPWR.n1542 VPWR.n1540 20.3299
R8060 VPWR.n1581 VPWR 20.3299
R8061 VPWR.n1582 VPWR.n1581 20.3299
R8062 VPWR.n1582 VPWR 20.3299
R8063 VPWR.n1583 VPWR.n1582 20.3299
R8064 VPWR.n1583 VPWR 20.3299
R8065 VPWR.n1584 VPWR.n1583 20.3299
R8066 VPWR.n1584 VPWR 20.3299
R8067 VPWR.n1585 VPWR.n1584 20.3299
R8068 VPWR.n1585 VPWR 20.3299
R8069 VPWR.n1586 VPWR.n1585 20.3299
R8070 VPWR VPWR.n1586 20.3299
R8071 VPWR.n1588 VPWR 20.3299
R8072 VPWR.n1587 VPWR 20.3299
R8073 VPWR.n1590 VPWR.n1588 20.3299
R8074 VPWR.n1590 VPWR 20.3299
R8075 VPWR.n1592 VPWR.n1590 20.3299
R8076 VPWR.n1592 VPWR 20.3299
R8077 VPWR.n1594 VPWR.n1592 20.3299
R8078 VPWR.n1594 VPWR 20.3299
R8079 VPWR.n1596 VPWR.n1594 20.3299
R8080 VPWR.n1596 VPWR 20.3299
R8081 VPWR.n1598 VPWR.n1596 20.3299
R8082 VPWR.n1598 VPWR 20.3299
R8083 VPWR.n1600 VPWR.n1598 20.3299
R8084 VPWR VPWR.n954 20.3299
R8085 VPWR.n780 VPWR 20.3299
R8086 VPWR.n931 VPWR 20.3299
R8087 VPWR VPWR.n952 20.3299
R8088 VPWR.n1742 VPWR 20.3299
R8089 VPWR.n327 VPWR 20.3299
R8090 VPWR VPWR.n1779 20.3299
R8091 VPWR VPWR.n1900 20.3299
R8092 VPWR VPWR.n624 20.3299
R8093 VPWR.n450 VPWR 20.3299
R8094 VPWR.n601 VPWR 20.3299
R8095 VPWR VPWR.n622 20.3299
R8096 VPWR VPWR.n1166 20.3299
R8097 VPWR.n1130 VPWR 20.3299
R8098 VPWR VPWR.n1103 20.3299
R8099 VPWR VPWR.n1028 20.3299
R8100 VPWR.n1064 VPWR 20.3299
R8101 VPWR.n1007 VPWR 20.3299
R8102 VPWR VPWR.n2280 20.3299
R8103 VPWR VPWR.n2335 20.3299
R8104 VPWR.n1174 VPWR 18.6711
R8105 VPWR.n1017 VPWR 15.2133
R8106 VPWR VPWR.n2080 15.2133
R8107 VPWR.n177 VPWR 15.2133
R8108 VPWR.n178 VPWR 15.2133
R8109 VPWR.n180 VPWR 15.2133
R8110 VPWR.n182 VPWR 15.2133
R8111 VPWR.n184 VPWR 15.2133
R8112 VPWR.n186 VPWR 15.2133
R8113 VPWR.n188 VPWR 15.2133
R8114 VPWR.n190 VPWR 15.2133
R8115 VPWR.n192 VPWR 15.2133
R8116 VPWR VPWR.n2146 15.2133
R8117 VPWR.n137 VPWR 15.2133
R8118 VPWR.n138 VPWR 15.2133
R8119 VPWR.n140 VPWR 15.2133
R8120 VPWR.n142 VPWR 15.2133
R8121 VPWR.n144 VPWR 15.2133
R8122 VPWR.n146 VPWR 15.2133
R8123 VPWR.n148 VPWR 15.2133
R8124 VPWR.n150 VPWR 15.2133
R8125 VPWR.n152 VPWR 15.2133
R8126 VPWR VPWR.n2212 15.2133
R8127 VPWR.n97 VPWR 15.2133
R8128 VPWR.n98 VPWR 15.2133
R8129 VPWR.n100 VPWR 15.2133
R8130 VPWR.n102 VPWR 15.2133
R8131 VPWR.n104 VPWR 15.2133
R8132 VPWR.n106 VPWR 15.2133
R8133 VPWR.n108 VPWR 15.2133
R8134 VPWR.n110 VPWR 15.2133
R8135 VPWR.n112 VPWR 15.2133
R8136 VPWR VPWR.n1312 15.2133
R8137 VPWR.n1280 VPWR 15.2133
R8138 VPWR VPWR.n1278 15.2133
R8139 VPWR.n1282 VPWR 15.2133
R8140 VPWR.n1284 VPWR 15.2133
R8141 VPWR.n1286 VPWR 15.2133
R8142 VPWR.n1288 VPWR 15.2133
R8143 VPWR.n1290 VPWR 15.2133
R8144 VPWR.n1292 VPWR 15.2133
R8145 VPWR.n1294 VPWR 15.2133
R8146 VPWR.n1297 VPWR 15.2133
R8147 VPWR.n1299 VPWR 15.2133
R8148 VPWR.n1301 VPWR 15.2133
R8149 VPWR.n1303 VPWR 15.2133
R8150 VPWR.n1305 VPWR 15.2133
R8151 VPWR.n1307 VPWR 15.2133
R8152 VPWR.n1309 VPWR 15.2133
R8153 VPWR VPWR.n949 15.2133
R8154 VPWR VPWR.n741 15.2133
R8155 VPWR.n933 VPWR 15.2133
R8156 VPWR VPWR.n950 15.2133
R8157 VPWR.n726 VPWR 15.2133
R8158 VPWR.n727 VPWR 15.2133
R8159 VPWR.n728 VPWR 15.2133
R8160 VPWR.n729 VPWR 15.2133
R8161 VPWR.n730 VPWR 15.2133
R8162 VPWR.n731 VPWR 15.2133
R8163 VPWR.n732 VPWR 15.2133
R8164 VPWR.n734 VPWR 15.2133
R8165 VPWR.n735 VPWR 15.2133
R8166 VPWR.n736 VPWR 15.2133
R8167 VPWR.n737 VPWR 15.2133
R8168 VPWR.n738 VPWR 15.2133
R8169 VPWR.n739 VPWR 15.2133
R8170 VPWR VPWR.n1777 15.2133
R8171 VPWR.n1745 VPWR 15.2133
R8172 VPWR VPWR.n1743 15.2133
R8173 VPWR.n1747 VPWR 15.2133
R8174 VPWR.n1749 VPWR 15.2133
R8175 VPWR.n1751 VPWR 15.2133
R8176 VPWR.n1753 VPWR 15.2133
R8177 VPWR.n1755 VPWR 15.2133
R8178 VPWR.n1757 VPWR 15.2133
R8179 VPWR.n1759 VPWR 15.2133
R8180 VPWR.n1762 VPWR 15.2133
R8181 VPWR.n1764 VPWR 15.2133
R8182 VPWR.n1766 VPWR 15.2133
R8183 VPWR.n1768 VPWR 15.2133
R8184 VPWR.n1770 VPWR 15.2133
R8185 VPWR.n1772 VPWR 15.2133
R8186 VPWR.n1774 VPWR 15.2133
R8187 VPWR VPWR.n619 15.2133
R8188 VPWR VPWR.n411 15.2133
R8189 VPWR.n603 VPWR 15.2133
R8190 VPWR VPWR.n620 15.2133
R8191 VPWR.n396 VPWR 15.2133
R8192 VPWR.n397 VPWR 15.2133
R8193 VPWR.n398 VPWR 15.2133
R8194 VPWR.n399 VPWR 15.2133
R8195 VPWR.n400 VPWR 15.2133
R8196 VPWR.n401 VPWR 15.2133
R8197 VPWR.n402 VPWR 15.2133
R8198 VPWR.n404 VPWR 15.2133
R8199 VPWR.n405 VPWR 15.2133
R8200 VPWR.n406 VPWR 15.2133
R8201 VPWR.n407 VPWR 15.2133
R8202 VPWR.n408 VPWR 15.2133
R8203 VPWR.n409 VPWR 15.2133
R8204 VPWR.n1009 VPWR 15.2133
R8205 VPWR VPWR.n1026 15.2133
R8206 VPWR.n1013 VPWR 15.2133
R8207 VPWR.n1066 VPWR 15.2133
R8208 VPWR VPWR.n984 15.2133
R8209 VPWR VPWR.n998 15.2133
R8210 VPWR.n1011 VPWR 15.2133
R8211 VPWR.n1015 VPWR 15.2133
R8212 VPWR.n1016 VPWR 15.2133
R8213 VPWR.n1019 VPWR 15.2133
R8214 VPWR.n1020 VPWR 15.2133
R8215 VPWR VPWR.n2278 15.2133
R8216 VPWR.n50 VPWR 15.2133
R8217 VPWR.n51 VPWR 15.2133
R8218 VPWR.n53 VPWR 15.2133
R8219 VPWR.n55 VPWR 15.2133
R8220 VPWR.n57 VPWR 15.2133
R8221 VPWR.n59 VPWR 15.2133
R8222 VPWR.n61 VPWR 15.2133
R8223 VPWR.n63 VPWR 15.2133
R8224 VPWR.n65 VPWR 15.2133
R8225 VPWR.n1253 VPWR 15.2129
R8226 VPWR.n1251 VPWR 15.2129
R8227 VPWR.n1250 VPWR 15.2129
R8228 VPWR.n1258 VPWR 15.2129
R8229 VPWR.n1256 VPWR 15.2129
R8230 VPWR.n1255 VPWR 15.2129
R8231 VPWR.n1263 VPWR 15.2129
R8232 VPWR.n1261 VPWR 15.2129
R8233 VPWR.n1260 VPWR 15.2129
R8234 VPWR.n1268 VPWR 15.2129
R8235 VPWR.n1266 VPWR 15.2129
R8236 VPWR.n1265 VPWR 15.2129
R8237 VPWR.n659 VPWR 15.2129
R8238 VPWR.n657 VPWR 15.2129
R8239 VPWR.n656 VPWR 15.2129
R8240 VPWR.n664 VPWR 15.2129
R8241 VPWR.n662 VPWR 15.2129
R8242 VPWR.n661 VPWR 15.2129
R8243 VPWR.n669 VPWR 15.2129
R8244 VPWR.n667 VPWR 15.2129
R8245 VPWR.n666 VPWR 15.2129
R8246 VPWR.n674 VPWR 15.2129
R8247 VPWR.n672 VPWR 15.2129
R8248 VPWR.n671 VPWR 15.2129
R8249 VPWR.n201 VPWR 15.2129
R8250 VPWR.n199 VPWR 15.2129
R8251 VPWR.n198 VPWR 15.2129
R8252 VPWR.n206 VPWR 15.2129
R8253 VPWR.n204 VPWR 15.2129
R8254 VPWR.n203 VPWR 15.2129
R8255 VPWR.n211 VPWR 15.2129
R8256 VPWR.n209 VPWR 15.2129
R8257 VPWR.n208 VPWR 15.2129
R8258 VPWR.n216 VPWR 15.2129
R8259 VPWR.n214 VPWR 15.2129
R8260 VPWR.n213 VPWR 15.2129
R8261 VPWR.n348 VPWR 15.2129
R8262 VPWR.n346 VPWR 15.2129
R8263 VPWR.n345 VPWR 15.2129
R8264 VPWR.n353 VPWR 15.2129
R8265 VPWR.n351 VPWR 15.2129
R8266 VPWR.n350 VPWR 15.2129
R8267 VPWR.n358 VPWR 15.2129
R8268 VPWR.n356 VPWR 15.2129
R8269 VPWR.n355 VPWR 15.2129
R8270 VPWR.n363 VPWR 15.2129
R8271 VPWR.n361 VPWR 15.2129
R8272 VPWR.n360 VPWR 15.2129
R8273 VPWR.n2003 VPWR.n2002 12.8005
R8274 VPWR.n2074 VPWR.n2001 12.8005
R8275 VPWR.n174 VPWR.n173 12.8005
R8276 VPWR.n2139 VPWR.n172 12.8005
R8277 VPWR.n134 VPWR.n133 12.8005
R8278 VPWR.n2205 VPWR.n132 12.8005
R8279 VPWR.n94 VPWR.n93 12.8005
R8280 VPWR.n2271 VPWR.n92 12.8005
R8281 VPWR.n1441 VPWR.n1177 12.8005
R8282 VPWR.n1244 VPWR.n1211 12.8005
R8283 VPWR.n1240 VPWR.n1239 12.8005
R8284 VPWR.n1437 VPWR.n1436 12.8005
R8285 VPWR.n1730 VPWR.n1453 12.8005
R8286 VPWR.n1608 VPWR.n1510 12.8005
R8287 VPWR.n1604 VPWR.n1603 12.8005
R8288 VPWR.n1726 VPWR.n1725 12.8005
R8289 VPWR.n744 VPWR.n743 12.8005
R8290 VPWR.n960 VPWR.n724 12.8005
R8291 VPWR.n956 VPWR.n955 12.8005
R8292 VPWR.n773 VPWR.n772 12.8005
R8293 VPWR.n1906 VPWR.n256 12.8005
R8294 VPWR.n323 VPWR.n290 12.8005
R8295 VPWR.n319 VPWR.n318 12.8005
R8296 VPWR.n1902 VPWR.n1901 12.8005
R8297 VPWR.n1916 VPWR.n1915 12.8005
R8298 VPWR.n1943 VPWR.n1914 12.8005
R8299 VPWR.n1948 VPWR.n1947 12.8005
R8300 VPWR.n1953 VPWR.n1952 12.8005
R8301 VPWR.n1958 VPWR.n1957 12.8005
R8302 VPWR.n414 VPWR.n413 12.8005
R8303 VPWR.n630 VPWR.n394 12.8005
R8304 VPWR.n626 VPWR.n625 12.8005
R8305 VPWR.n443 VPWR.n442 12.8005
R8306 VPWR.n1093 VPWR.n1092 12.8005
R8307 VPWR.n1168 VPWR.n1070 12.8005
R8308 VPWR.n1072 VPWR.n1071 12.8005
R8309 VPWR.n1126 VPWR.n1089 12.8005
R8310 VPWR.n1112 VPWR.n1111 12.8005
R8311 VPWR.n1105 VPWR.n1091 12.8005
R8312 VPWR.n1173 VPWR 12.8005
R8313 VPWR.n47 VPWR.n46 12.8005
R8314 VPWR.n2337 VPWR.n45 12.8005
R8315 VPWR.n372 VPWR 10.6653
R8316 VPWR.n370 VPWR 10.6653
R8317 VPWR.n369 VPWR 10.6653
R8318 VPWR.n377 VPWR 10.6653
R8319 VPWR.n375 VPWR 10.6653
R8320 VPWR.n374 VPWR 10.6653
R8321 VPWR.n382 VPWR 10.6653
R8322 VPWR.n380 VPWR 10.6653
R8323 VPWR.n379 VPWR 10.6653
R8324 VPWR.n387 VPWR 10.6653
R8325 VPWR.n385 VPWR 10.6653
R8326 VPWR.n384 VPWR 10.6653
R8327 VPWR.n6 VPWR 10.6653
R8328 VPWR.n4 VPWR 10.6653
R8329 VPWR.n3 VPWR 10.6653
R8330 VPWR.n11 VPWR 10.6653
R8331 VPWR.n9 VPWR 10.6653
R8332 VPWR.n8 VPWR 10.6653
R8333 VPWR.n16 VPWR 10.6653
R8334 VPWR.n14 VPWR 10.6653
R8335 VPWR.n13 VPWR 10.6653
R8336 VPWR.n21 VPWR 10.6653
R8337 VPWR.n19 VPWR 10.6653
R8338 VPWR.n18 VPWR 10.6653
R8339 VPWR.n702 VPWR 10.6653
R8340 VPWR.n700 VPWR 10.6653
R8341 VPWR.n699 VPWR 10.6653
R8342 VPWR.n707 VPWR 10.6653
R8343 VPWR.n705 VPWR 10.6653
R8344 VPWR.n704 VPWR 10.6653
R8345 VPWR.n712 VPWR 10.6653
R8346 VPWR.n710 VPWR 10.6653
R8347 VPWR.n709 VPWR 10.6653
R8348 VPWR.n717 VPWR 10.6653
R8349 VPWR.n715 VPWR 10.6653
R8350 VPWR.n714 VPWR 10.6653
R8351 VPWR.n233 VPWR 10.6653
R8352 VPWR.n231 VPWR 10.6653
R8353 VPWR.n230 VPWR 10.6653
R8354 VPWR.n238 VPWR 10.6653
R8355 VPWR.n236 VPWR 10.6653
R8356 VPWR.n235 VPWR 10.6653
R8357 VPWR.n243 VPWR 10.6653
R8358 VPWR.n241 VPWR 10.6653
R8359 VPWR.n240 VPWR 10.6653
R8360 VPWR.n248 VPWR 10.6653
R8361 VPWR.n246 VPWR 10.6653
R8362 VPWR.n245 VPWR 10.6653
R8363 VPWR.n1980 VPWR 10.6647
R8364 VPWR.n1981 VPWR 10.6647
R8365 VPWR.n1983 VPWR 10.6647
R8366 VPWR.n1985 VPWR 10.6647
R8367 VPWR.n1987 VPWR 10.6647
R8368 VPWR.n1989 VPWR 10.6647
R8369 VPWR.n1991 VPWR 10.6647
R8370 VPWR.n1994 VPWR 10.6647
R8371 VPWR.n1996 VPWR 10.6647
R8372 VPWR.n1998 VPWR 10.6647
R8373 VPWR.n156 VPWR 10.6647
R8374 VPWR.n157 VPWR 10.6647
R8375 VPWR.n159 VPWR 10.6647
R8376 VPWR.n161 VPWR 10.6647
R8377 VPWR.n163 VPWR 10.6647
R8378 VPWR.n165 VPWR 10.6647
R8379 VPWR.n167 VPWR 10.6647
R8380 VPWR.n169 VPWR 10.6647
R8381 VPWR.n116 VPWR 10.6647
R8382 VPWR.n117 VPWR 10.6647
R8383 VPWR.n119 VPWR 10.6647
R8384 VPWR.n121 VPWR 10.6647
R8385 VPWR.n123 VPWR 10.6647
R8386 VPWR.n125 VPWR 10.6647
R8387 VPWR.n127 VPWR 10.6647
R8388 VPWR.n129 VPWR 10.6647
R8389 VPWR.n76 VPWR 10.6647
R8390 VPWR.n77 VPWR 10.6647
R8391 VPWR.n79 VPWR 10.6647
R8392 VPWR.n81 VPWR 10.6647
R8393 VPWR.n83 VPWR 10.6647
R8394 VPWR.n85 VPWR 10.6647
R8395 VPWR.n87 VPWR 10.6647
R8396 VPWR.n89 VPWR 10.6647
R8397 VPWR.n1212 VPWR 10.6647
R8398 VPWR.n1214 VPWR 10.6647
R8399 VPWR.n1216 VPWR 10.6647
R8400 VPWR.n1218 VPWR 10.6647
R8401 VPWR.n1220 VPWR 10.6647
R8402 VPWR.n1222 VPWR 10.6647
R8403 VPWR.n1224 VPWR 10.6647
R8404 VPWR.n1227 VPWR 10.6647
R8405 VPWR.n1229 VPWR 10.6647
R8406 VPWR.n1231 VPWR 10.6647
R8407 VPWR.n1233 VPWR 10.6647
R8408 VPWR.n1235 VPWR 10.6647
R8409 VPWR.n1237 VPWR 10.6647
R8410 VPWR.n1513 VPWR 10.6647
R8411 VPWR.n1515 VPWR 10.6647
R8412 VPWR.n1517 VPWR 10.6647
R8413 VPWR.n1519 VPWR 10.6647
R8414 VPWR.n1521 VPWR 10.6647
R8415 VPWR.n1543 VPWR 10.6647
R8416 VPWR.n1545 VPWR 10.6647
R8417 VPWR.n1548 VPWR 10.6647
R8418 VPWR.n1551 VPWR 10.6647
R8419 VPWR.n1554 VPWR 10.6647
R8420 VPWR.n1556 VPWR 10.6647
R8421 VPWR.n1559 VPWR 10.6647
R8422 VPWR.n1561 VPWR 10.6647
R8423 VPWR.n1563 VPWR 10.6647
R8424 VPWR.n1566 VPWR 10.6647
R8425 VPWR.n1568 VPWR 10.6647
R8426 VPWR.n1570 VPWR 10.6647
R8427 VPWR.n1573 VPWR 10.6647
R8428 VPWR.n1576 VPWR 10.6647
R8429 VPWR.n1579 VPWR 10.6647
R8430 VPWR.n1601 VPWR 10.6647
R8431 VPWR.n745 VPWR 10.6647
R8432 VPWR.n747 VPWR 10.6647
R8433 VPWR.n749 VPWR 10.6647
R8434 VPWR.n751 VPWR 10.6647
R8435 VPWR.n753 VPWR 10.6647
R8436 VPWR.n755 VPWR 10.6647
R8437 VPWR.n757 VPWR 10.6647
R8438 VPWR.n760 VPWR 10.6647
R8439 VPWR.n762 VPWR 10.6647
R8440 VPWR.n764 VPWR 10.6647
R8441 VPWR.n766 VPWR 10.6647
R8442 VPWR.n768 VPWR 10.6647
R8443 VPWR.n770 VPWR 10.6647
R8444 VPWR.n291 VPWR 10.6647
R8445 VPWR.n293 VPWR 10.6647
R8446 VPWR.n295 VPWR 10.6647
R8447 VPWR.n297 VPWR 10.6647
R8448 VPWR.n299 VPWR 10.6647
R8449 VPWR.n301 VPWR 10.6647
R8450 VPWR.n303 VPWR 10.6647
R8451 VPWR.n306 VPWR 10.6647
R8452 VPWR.n308 VPWR 10.6647
R8453 VPWR.n310 VPWR 10.6647
R8454 VPWR.n312 VPWR 10.6647
R8455 VPWR.n314 VPWR 10.6647
R8456 VPWR.n316 VPWR 10.6647
R8457 VPWR.n415 VPWR 10.6647
R8458 VPWR.n417 VPWR 10.6647
R8459 VPWR.n419 VPWR 10.6647
R8460 VPWR.n421 VPWR 10.6647
R8461 VPWR.n423 VPWR 10.6647
R8462 VPWR.n425 VPWR 10.6647
R8463 VPWR.n427 VPWR 10.6647
R8464 VPWR.n430 VPWR 10.6647
R8465 VPWR.n432 VPWR 10.6647
R8466 VPWR.n434 VPWR 10.6647
R8467 VPWR.n436 VPWR 10.6647
R8468 VPWR.n438 VPWR 10.6647
R8469 VPWR.n440 VPWR 10.6647
R8470 VPWR.n1109 VPWR 10.6647
R8471 VPWR.n1115 VPWR 10.6647
R8472 VPWR.n1116 VPWR 10.6647
R8473 VPWR.n1119 VPWR 10.6647
R8474 VPWR.n1120 VPWR 10.6647
R8475 VPWR.n29 VPWR 10.6647
R8476 VPWR.n30 VPWR 10.6647
R8477 VPWR.n32 VPWR 10.6647
R8478 VPWR.n34 VPWR 10.6647
R8479 VPWR.n36 VPWR 10.6647
R8480 VPWR.n38 VPWR 10.6647
R8481 VPWR.n40 VPWR 10.6647
R8482 VPWR.n42 VPWR 10.6647
R8483 VPWR.n1512 VPWR 10.6647
R8484 VPWR.n1511 VPWR 10.6647
R8485 VPWR.n1117 VPWR 10.6647
R8486 VPWR.n2025 VPWR.n2019 10.4301
R8487 VPWR.n2028 VPWR.n2026 10.4301
R8488 VPWR.n2036 VPWR.n2035 10.4301
R8489 VPWR.n2038 VPWR.n2037 10.4301
R8490 VPWR.n2046 VPWR.n2045 10.4301
R8491 VPWR.n2054 VPWR.n2011 10.4301
R8492 VPWR.n2057 VPWR.n2056 10.4301
R8493 VPWR.n2065 VPWR.n2064 10.4301
R8494 VPWR.n2066 VPWR.n2006 10.4301
R8495 VPWR.n2132 VPWR.n2131 10.4301
R8496 VPWR.n2127 VPWR.n2124 10.4301
R8497 VPWR.n2120 VPWR.n2119 10.4301
R8498 VPWR.n2116 VPWR.n2115 10.4301
R8499 VPWR.n2111 VPWR.n2108 10.4301
R8500 VPWR.n2104 VPWR.n2103 10.4301
R8501 VPWR.n2100 VPWR.n2099 10.4301
R8502 VPWR.n2096 VPWR.n2083 10.4301
R8503 VPWR.n2198 VPWR.n2197 10.4301
R8504 VPWR.n2193 VPWR.n2190 10.4301
R8505 VPWR.n2186 VPWR.n2185 10.4301
R8506 VPWR.n2182 VPWR.n2181 10.4301
R8507 VPWR.n2177 VPWR.n2174 10.4301
R8508 VPWR.n2170 VPWR.n2169 10.4301
R8509 VPWR.n2166 VPWR.n2165 10.4301
R8510 VPWR.n2162 VPWR.n2149 10.4301
R8511 VPWR.n2264 VPWR.n2263 10.4301
R8512 VPWR.n2259 VPWR.n2256 10.4301
R8513 VPWR.n2252 VPWR.n2251 10.4301
R8514 VPWR.n2248 VPWR.n2247 10.4301
R8515 VPWR.n2243 VPWR.n2240 10.4301
R8516 VPWR.n2236 VPWR.n2235 10.4301
R8517 VPWR.n2232 VPWR.n2231 10.4301
R8518 VPWR.n2228 VPWR.n2215 10.4301
R8519 VPWR.n1433 VPWR.n1179 10.4301
R8520 VPWR.n1317 VPWR.n1316 10.4301
R8521 VPWR.n1324 VPWR.n1321 10.4301
R8522 VPWR.n1328 VPWR.n1325 10.4301
R8523 VPWR.n1333 VPWR.n1332 10.4301
R8524 VPWR.n1337 VPWR.n1336 10.4301
R8525 VPWR.n1341 VPWR.n1340 10.4301
R8526 VPWR.n1352 VPWR.n1349 10.4301
R8527 VPWR.n1361 VPWR.n1360 10.4301
R8528 VPWR.n1372 VPWR.n1369 10.4301
R8529 VPWR.n1381 VPWR.n1380 10.4301
R8530 VPWR.n1392 VPWR.n1389 10.4301
R8531 VPWR.n1400 VPWR.n1397 10.4301
R8532 VPWR.n1408 VPWR.n1405 10.4301
R8533 VPWR.n1412 VPWR.n1409 10.4301
R8534 VPWR.n1416 VPWR.n1413 10.4301
R8535 VPWR.n1420 VPWR.n1417 10.4301
R8536 VPWR.n1424 VPWR.n1421 10.4301
R8537 VPWR.n1427 VPWR.n1426 10.4301
R8538 VPWR.n1722 VPWR.n1455 10.4301
R8539 VPWR.n1716 VPWR.n1715 10.4301
R8540 VPWR.n1708 VPWR.n1461 10.4301
R8541 VPWR.n1706 VPWR.n1462 10.4301
R8542 VPWR.n1700 VPWR.n1699 10.4301
R8543 VPWR.n1684 VPWR.n1683 10.4301
R8544 VPWR.n1668 VPWR.n1667 10.4301
R8545 VPWR.n1659 VPWR.n1658 10.4301
R8546 VPWR.n1650 VPWR.n1490 10.4301
R8547 VPWR.n1634 VPWR.n1498 10.4301
R8548 VPWR.n1618 VPWR.n1506 10.4301
R8549 VPWR.n814 VPWR.n813 10.4301
R8550 VPWR.n818 VPWR.n817 10.4301
R8551 VPWR.n825 VPWR.n822 10.4301
R8552 VPWR.n829 VPWR.n826 10.4301
R8553 VPWR.n834 VPWR.n833 10.4301
R8554 VPWR.n838 VPWR.n837 10.4301
R8555 VPWR.n842 VPWR.n841 10.4301
R8556 VPWR.n853 VPWR.n850 10.4301
R8557 VPWR.n862 VPWR.n861 10.4301
R8558 VPWR.n873 VPWR.n870 10.4301
R8559 VPWR.n882 VPWR.n881 10.4301
R8560 VPWR.n893 VPWR.n890 10.4301
R8561 VPWR.n901 VPWR.n898 10.4301
R8562 VPWR.n909 VPWR.n906 10.4301
R8563 VPWR.n913 VPWR.n910 10.4301
R8564 VPWR.n917 VPWR.n914 10.4301
R8565 VPWR.n921 VPWR.n918 10.4301
R8566 VPWR.n924 VPWR.n923 10.4301
R8567 VPWR.n925 VPWR.n781 10.4301
R8568 VPWR.n1898 VPWR.n258 10.4301
R8569 VPWR.n1782 VPWR.n1781 10.4301
R8570 VPWR.n1789 VPWR.n1786 10.4301
R8571 VPWR.n1793 VPWR.n1790 10.4301
R8572 VPWR.n1798 VPWR.n1797 10.4301
R8573 VPWR.n1802 VPWR.n1801 10.4301
R8574 VPWR.n1806 VPWR.n1805 10.4301
R8575 VPWR.n1817 VPWR.n1814 10.4301
R8576 VPWR.n1826 VPWR.n1825 10.4301
R8577 VPWR.n1837 VPWR.n1834 10.4301
R8578 VPWR.n1846 VPWR.n1845 10.4301
R8579 VPWR.n1857 VPWR.n1854 10.4301
R8580 VPWR.n1865 VPWR.n1862 10.4301
R8581 VPWR.n1873 VPWR.n1870 10.4301
R8582 VPWR.n1877 VPWR.n1874 10.4301
R8583 VPWR.n1881 VPWR.n1878 10.4301
R8584 VPWR.n1885 VPWR.n1882 10.4301
R8585 VPWR.n1889 VPWR.n1886 10.4301
R8586 VPWR.n1892 VPWR.n1891 10.4301
R8587 VPWR.n1938 VPWR.n1920 10.4301
R8588 VPWR.n1932 VPWR.n1931 10.4301
R8589 VPWR.n1930 VPWR.n1924 10.4301
R8590 VPWR.n484 VPWR.n483 10.4301
R8591 VPWR.n488 VPWR.n487 10.4301
R8592 VPWR.n495 VPWR.n492 10.4301
R8593 VPWR.n499 VPWR.n496 10.4301
R8594 VPWR.n504 VPWR.n503 10.4301
R8595 VPWR.n508 VPWR.n507 10.4301
R8596 VPWR.n512 VPWR.n511 10.4301
R8597 VPWR.n523 VPWR.n520 10.4301
R8598 VPWR.n532 VPWR.n531 10.4301
R8599 VPWR.n543 VPWR.n540 10.4301
R8600 VPWR.n552 VPWR.n551 10.4301
R8601 VPWR.n563 VPWR.n560 10.4301
R8602 VPWR.n571 VPWR.n568 10.4301
R8603 VPWR.n579 VPWR.n576 10.4301
R8604 VPWR.n583 VPWR.n580 10.4301
R8605 VPWR.n587 VPWR.n584 10.4301
R8606 VPWR.n591 VPWR.n588 10.4301
R8607 VPWR.n594 VPWR.n593 10.4301
R8608 VPWR.n595 VPWR.n451 10.4301
R8609 VPWR.n1101 VPWR.n1096 10.4301
R8610 VPWR.n1132 VPWR.n1087 10.4301
R8611 VPWR.n1138 VPWR.n1083 10.4301
R8612 VPWR.n1141 VPWR.n1139 10.4301
R8613 VPWR.n1149 VPWR.n1148 10.4301
R8614 VPWR.n1159 VPWR.n1158 10.4301
R8615 VPWR.n1160 VPWR.n1075 10.4301
R8616 VPWR.n1005 VPWR.n1000 10.4301
R8617 VPWR.n1030 VPWR.n997 10.4301
R8618 VPWR.n1036 VPWR.n993 10.4301
R8619 VPWR.n1039 VPWR.n1037 10.4301
R8620 VPWR.n1047 VPWR.n1046 10.4301
R8621 VPWR.n1057 VPWR.n1056 10.4301
R8622 VPWR.n1058 VPWR.n985 10.4301
R8623 VPWR.n2330 VPWR.n2329 10.4301
R8624 VPWR.n2325 VPWR.n2322 10.4301
R8625 VPWR.n2318 VPWR.n2317 10.4301
R8626 VPWR.n2314 VPWR.n2313 10.4301
R8627 VPWR.n2309 VPWR.n2306 10.4301
R8628 VPWR.n2302 VPWR.n2301 10.4301
R8629 VPWR.n2298 VPWR.n2297 10.4301
R8630 VPWR.n2294 VPWR.n2281 10.4301
R8631 VPWR.n1022 VPWR.n1017 9.57565
R8632 VPWR.n1915 VPWR.n1913 9.3947
R8633 VPWR.n1945 VPWR.n1914 9.3947
R8634 VPWR.n1950 VPWR.n1947 9.3947
R8635 VPWR.n1955 VPWR.n1952 9.3947
R8636 VPWR.n1960 VPWR.n1957 9.3947
R8637 VPWR.n2004 VPWR.n2003 9.39464
R8638 VPWR.n2076 VPWR.n2001 9.39464
R8639 VPWR.n2076 VPWR.n2075 9.39464
R8640 VPWR.n2005 VPWR.n2004 9.39464
R8641 VPWR.n175 VPWR.n174 9.39464
R8642 VPWR.n2141 VPWR.n172 9.39464
R8643 VPWR.n2141 VPWR.n2140 9.39464
R8644 VPWR.n176 VPWR.n175 9.39464
R8645 VPWR.n135 VPWR.n134 9.39464
R8646 VPWR.n2207 VPWR.n132 9.39464
R8647 VPWR.n2207 VPWR.n2206 9.39464
R8648 VPWR.n136 VPWR.n135 9.39464
R8649 VPWR.n95 VPWR.n94 9.39464
R8650 VPWR.n2273 VPWR.n92 9.39464
R8651 VPWR.n2273 VPWR.n2272 9.39464
R8652 VPWR.n96 VPWR.n95 9.39464
R8653 VPWR.n1443 VPWR.n1177 9.39464
R8654 VPWR.n1245 VPWR.n1244 9.39464
R8655 VPWR.n1246 VPWR.n1245 9.39464
R8656 VPWR.n1241 VPWR.n1240 9.39464
R8657 VPWR.n1438 VPWR.n1437 9.39464
R8658 VPWR.n1439 VPWR.n1438 9.39464
R8659 VPWR.n1732 VPWR.n1453 9.39464
R8660 VPWR.n1609 VPWR.n1608 9.39464
R8661 VPWR.n1610 VPWR.n1609 9.39464
R8662 VPWR.n1605 VPWR.n1604 9.39464
R8663 VPWR.n1727 VPWR.n1726 9.39464
R8664 VPWR.n1728 VPWR.n1727 9.39464
R8665 VPWR.n1605 VPWR.n1509 9.39464
R8666 VPWR.n1732 VPWR.n1731 9.39464
R8667 VPWR.n777 VPWR.n744 9.39464
R8668 VPWR.n778 VPWR.n777 9.39464
R8669 VPWR.n962 VPWR.n724 9.39464
R8670 VPWR.n957 VPWR.n956 9.39464
R8671 VPWR.n958 VPWR.n957 9.39464
R8672 VPWR.n962 VPWR.n961 9.39464
R8673 VPWR.n774 VPWR.n742 9.39464
R8674 VPWR.n774 VPWR.n773 9.39464
R8675 VPWR.n1908 VPWR.n256 9.39464
R8676 VPWR.n324 VPWR.n323 9.39464
R8677 VPWR.n325 VPWR.n324 9.39464
R8678 VPWR.n320 VPWR.n319 9.39464
R8679 VPWR.n1903 VPWR.n1902 9.39464
R8680 VPWR.n1904 VPWR.n1903 9.39464
R8681 VPWR.n320 VPWR.n289 9.39464
R8682 VPWR.n1908 VPWR.n1907 9.39464
R8683 VPWR.n447 VPWR.n414 9.39464
R8684 VPWR.n448 VPWR.n447 9.39464
R8685 VPWR.n632 VPWR.n394 9.39464
R8686 VPWR.n627 VPWR.n626 9.39464
R8687 VPWR.n628 VPWR.n627 9.39464
R8688 VPWR.n632 VPWR.n631 9.39464
R8689 VPWR.n444 VPWR.n412 9.39464
R8690 VPWR.n444 VPWR.n443 9.39464
R8691 VPWR.n1092 VPWR.n1090 9.39464
R8692 VPWR.n1170 VPWR.n1070 9.39464
R8693 VPWR.n1170 VPWR.n1169 9.39464
R8694 VPWR.n1073 VPWR.n1072 9.39464
R8695 VPWR.n1127 VPWR.n1126 9.39464
R8696 VPWR.n1128 VPWR.n1127 9.39464
R8697 VPWR.n1113 VPWR.n1112 9.39464
R8698 VPWR.n1107 VPWR.n1091 9.39464
R8699 VPWR.n1107 VPWR.n1106 9.39464
R8700 VPWR.n1113 VPWR.n1088 9.39464
R8701 VPWR.n1074 VPWR.n1073 9.39464
R8702 VPWR.n1094 VPWR.n1090 9.39464
R8703 VPWR.n1241 VPWR.n1210 9.39464
R8704 VPWR.n1443 VPWR.n1442 9.39464
R8705 VPWR.n48 VPWR.n47 9.39464
R8706 VPWR.n2339 VPWR.n45 9.39464
R8707 VPWR.n2339 VPWR.n2338 9.39464
R8708 VPWR.n49 VPWR.n48 9.39464
R8709 VPWR.n1917 VPWR.n1913 9.39457
R8710 VPWR.n1945 VPWR.n1944 9.39457
R8711 VPWR.n1950 VPWR.n1949 9.39457
R8712 VPWR.n1955 VPWR.n1954 9.39457
R8713 VPWR.n1960 VPWR.n1959 9.39457
R8714 VPWR.n1010 VPWR.n998 9.38993
R8715 VPWR VPWR.n177 9.36745
R8716 VPWR VPWR.n137 9.36745
R8717 VPWR VPWR.n97 9.36745
R8718 VPWR VPWR.n50 9.36745
R8719 VPWR.n193 VPWR.n192 9.34497
R8720 VPWR.n153 VPWR.n152 9.34497
R8721 VPWR.n113 VPWR.n112 9.34497
R8722 VPWR.n1310 VPWR.n1309 9.34497
R8723 VPWR.n1775 VPWR.n1774 9.34497
R8724 VPWR.n66 VPWR.n65 9.34497
R8725 VPWR.n2080 VPWR.n2079 9.34497
R8726 VPWR.n179 VPWR.n178 9.34497
R8727 VPWR.n181 VPWR.n180 9.34497
R8728 VPWR.n183 VPWR.n182 9.34497
R8729 VPWR.n185 VPWR.n184 9.34497
R8730 VPWR.n187 VPWR.n186 9.34497
R8731 VPWR.n189 VPWR.n188 9.34497
R8732 VPWR.n191 VPWR.n190 9.34497
R8733 VPWR.n2146 VPWR.n2145 9.34497
R8734 VPWR.n139 VPWR.n138 9.34497
R8735 VPWR.n141 VPWR.n140 9.34497
R8736 VPWR.n143 VPWR.n142 9.34497
R8737 VPWR.n145 VPWR.n144 9.34497
R8738 VPWR.n147 VPWR.n146 9.34497
R8739 VPWR.n149 VPWR.n148 9.34497
R8740 VPWR.n151 VPWR.n150 9.34497
R8741 VPWR.n2212 VPWR.n2211 9.34497
R8742 VPWR.n99 VPWR.n98 9.34497
R8743 VPWR.n101 VPWR.n100 9.34497
R8744 VPWR.n103 VPWR.n102 9.34497
R8745 VPWR.n105 VPWR.n104 9.34497
R8746 VPWR.n107 VPWR.n106 9.34497
R8747 VPWR.n109 VPWR.n108 9.34497
R8748 VPWR.n111 VPWR.n110 9.34497
R8749 VPWR.n1312 VPWR.n1311 9.34497
R8750 VPWR.n1278 VPWR.n1276 9.34497
R8751 VPWR.n1283 VPWR.n1282 9.34497
R8752 VPWR.n1285 VPWR.n1284 9.34497
R8753 VPWR.n1287 VPWR.n1286 9.34497
R8754 VPWR.n1289 VPWR.n1288 9.34497
R8755 VPWR.n1291 VPWR.n1290 9.34497
R8756 VPWR.n1293 VPWR.n1292 9.34497
R8757 VPWR.n1295 VPWR.n1294 9.34497
R8758 VPWR.n1298 VPWR.n1297 9.34497
R8759 VPWR.n1300 VPWR.n1299 9.34497
R8760 VPWR.n1302 VPWR.n1301 9.34497
R8761 VPWR.n1304 VPWR.n1303 9.34497
R8762 VPWR.n1306 VPWR.n1305 9.34497
R8763 VPWR.n1308 VPWR.n1307 9.34497
R8764 VPWR.n1281 VPWR.n1280 9.34497
R8765 VPWR.n934 VPWR.n933 9.34497
R8766 VPWR.n950 VPWR.n655 9.34497
R8767 VPWR.n947 VPWR.n726 9.34497
R8768 VPWR.n946 VPWR.n727 9.34497
R8769 VPWR.n945 VPWR.n728 9.34497
R8770 VPWR.n944 VPWR.n729 9.34497
R8771 VPWR.n943 VPWR.n730 9.34497
R8772 VPWR.n942 VPWR.n731 9.34497
R8773 VPWR.n941 VPWR.n732 9.34497
R8774 VPWR.n940 VPWR.n734 9.34497
R8775 VPWR.n939 VPWR.n735 9.34497
R8776 VPWR.n938 VPWR.n736 9.34497
R8777 VPWR.n937 VPWR.n737 9.34497
R8778 VPWR.n936 VPWR.n738 9.34497
R8779 VPWR.n935 VPWR.n739 9.34497
R8780 VPWR.n741 VPWR.n740 9.34497
R8781 VPWR.n949 VPWR.n948 9.34497
R8782 VPWR.n1777 VPWR.n1776 9.34497
R8783 VPWR.n1743 VPWR.n1741 9.34497
R8784 VPWR.n1748 VPWR.n1747 9.34497
R8785 VPWR.n1750 VPWR.n1749 9.34497
R8786 VPWR.n1752 VPWR.n1751 9.34497
R8787 VPWR.n1754 VPWR.n1753 9.34497
R8788 VPWR.n1756 VPWR.n1755 9.34497
R8789 VPWR.n1758 VPWR.n1757 9.34497
R8790 VPWR.n1760 VPWR.n1759 9.34497
R8791 VPWR.n1763 VPWR.n1762 9.34497
R8792 VPWR.n1765 VPWR.n1764 9.34497
R8793 VPWR.n1767 VPWR.n1766 9.34497
R8794 VPWR.n1769 VPWR.n1768 9.34497
R8795 VPWR.n1771 VPWR.n1770 9.34497
R8796 VPWR.n1773 VPWR.n1772 9.34497
R8797 VPWR.n1746 VPWR.n1745 9.34497
R8798 VPWR.n604 VPWR.n603 9.34497
R8799 VPWR.n620 VPWR.n343 9.34497
R8800 VPWR.n617 VPWR.n396 9.34497
R8801 VPWR.n616 VPWR.n397 9.34497
R8802 VPWR.n615 VPWR.n398 9.34497
R8803 VPWR.n614 VPWR.n399 9.34497
R8804 VPWR.n613 VPWR.n400 9.34497
R8805 VPWR.n612 VPWR.n401 9.34497
R8806 VPWR.n611 VPWR.n402 9.34497
R8807 VPWR.n610 VPWR.n404 9.34497
R8808 VPWR.n609 VPWR.n405 9.34497
R8809 VPWR.n608 VPWR.n406 9.34497
R8810 VPWR.n607 VPWR.n407 9.34497
R8811 VPWR.n606 VPWR.n408 9.34497
R8812 VPWR.n605 VPWR.n409 9.34497
R8813 VPWR.n411 VPWR.n410 9.34497
R8814 VPWR.n619 VPWR.n618 9.34497
R8815 VPWR.n1014 VPWR.n1013 9.34497
R8816 VPWR.n984 VPWR.n983 9.34497
R8817 VPWR.n1012 VPWR.n1011 9.34497
R8818 VPWR.n1024 VPWR.n1015 9.34497
R8819 VPWR.n1023 VPWR.n1016 9.34497
R8820 VPWR.n1022 VPWR.n1019 9.34497
R8821 VPWR.n1021 VPWR.n1020 9.34497
R8822 VPWR.n1067 VPWR.n1066 9.34497
R8823 VPWR.n1026 VPWR.n1025 9.34497
R8824 VPWR.n1010 VPWR.n1009 9.34497
R8825 VPWR.n2278 VPWR.n2277 9.34497
R8826 VPWR.n52 VPWR.n51 9.34497
R8827 VPWR.n54 VPWR.n53 9.34497
R8828 VPWR.n56 VPWR.n55 9.34497
R8829 VPWR.n58 VPWR.n57 9.34497
R8830 VPWR.n60 VPWR.n59 9.34497
R8831 VPWR.n62 VPWR.n61 9.34497
R8832 VPWR.n64 VPWR.n63 9.34497
R8833 VPWR.n1736 VPWR.n338 9.3005
R8834 VPWR.n1736 VPWR.n340 9.3005
R8835 VPWR.n1736 VPWR.n337 9.3005
R8836 VPWR.n1736 VPWR.n651 9.3005
R8837 VPWR.n1736 VPWR.n336 9.3005
R8838 VPWR.n1736 VPWR.n652 9.3005
R8839 VPWR.n1736 VPWR.n335 9.3005
R8840 VPWR.n1736 VPWR.n972 9.3005
R8841 VPWR.n1736 VPWR.n334 9.3005
R8842 VPWR.n1736 VPWR.n977 9.3005
R8843 VPWR.n1736 VPWR.n333 9.3005
R8844 VPWR.n1736 VPWR.n978 9.3005
R8845 VPWR.n1737 VPWR.n1736 9.3005
R8846 VPWR.n1736 VPWR.n1735 9.3005
R8847 VPWR.n1736 VPWR.n332 9.3005
R8848 VPWR.n1451 VPWR.n338 9.3005
R8849 VPWR.n1451 VPWR.n340 9.3005
R8850 VPWR.n1451 VPWR.n337 9.3005
R8851 VPWR.n1451 VPWR.n652 9.3005
R8852 VPWR.n1451 VPWR.n335 9.3005
R8853 VPWR.n1735 VPWR.n1451 9.3005
R8854 VPWR.n1451 VPWR.n332 9.3005
R8855 VPWR.n1451 VPWR.n979 9.3005
R8856 VPWR.n1451 VPWR.n1450 9.3005
R8857 VPWR.n1254 VPWR.n1251 8.5126
R8858 VPWR.n1254 VPWR.n1250 8.5126
R8859 VPWR.n1259 VPWR.n1256 8.5126
R8860 VPWR.n1259 VPWR.n1255 8.5126
R8861 VPWR.n1264 VPWR.n1261 8.5126
R8862 VPWR.n1264 VPWR.n1260 8.5126
R8863 VPWR.n1269 VPWR.n1266 8.5126
R8864 VPWR.n1269 VPWR.n1265 8.5126
R8865 VPWR.n660 VPWR.n657 8.5126
R8866 VPWR.n660 VPWR.n656 8.5126
R8867 VPWR.n665 VPWR.n662 8.5126
R8868 VPWR.n665 VPWR.n661 8.5126
R8869 VPWR.n670 VPWR.n667 8.5126
R8870 VPWR.n670 VPWR.n666 8.5126
R8871 VPWR.n675 VPWR.n672 8.5126
R8872 VPWR.n675 VPWR.n671 8.5126
R8873 VPWR.n202 VPWR.n199 8.5126
R8874 VPWR.n202 VPWR.n198 8.5126
R8875 VPWR.n207 VPWR.n204 8.5126
R8876 VPWR.n207 VPWR.n203 8.5126
R8877 VPWR.n212 VPWR.n209 8.5126
R8878 VPWR.n212 VPWR.n208 8.5126
R8879 VPWR.n217 VPWR.n214 8.5126
R8880 VPWR.n217 VPWR.n213 8.5126
R8881 VPWR.n349 VPWR.n346 8.5126
R8882 VPWR.n349 VPWR.n345 8.5126
R8883 VPWR.n354 VPWR.n351 8.5126
R8884 VPWR.n354 VPWR.n350 8.5126
R8885 VPWR.n359 VPWR.n356 8.5126
R8886 VPWR.n359 VPWR.n355 8.5126
R8887 VPWR.n364 VPWR.n361 8.5126
R8888 VPWR.n364 VPWR.n360 8.5126
R8889 VPWR.n1552 VPWR.n1512 8.10069
R8890 VPWR.n1577 VPWR.n1511 8.10069
R8891 VPWR.n1122 VPWR.n1117 8.10069
R8892 VPWR.n1254 VPWR.n1253 7.99054
R8893 VPWR.n1259 VPWR.n1258 7.99054
R8894 VPWR.n1264 VPWR.n1263 7.99054
R8895 VPWR.n1269 VPWR.n1268 7.99054
R8896 VPWR.n660 VPWR.n659 7.99054
R8897 VPWR.n665 VPWR.n664 7.99054
R8898 VPWR.n670 VPWR.n669 7.99054
R8899 VPWR.n675 VPWR.n674 7.99054
R8900 VPWR.n202 VPWR.n201 7.99054
R8901 VPWR.n207 VPWR.n206 7.99054
R8902 VPWR.n212 VPWR.n211 7.99054
R8903 VPWR.n217 VPWR.n216 7.99054
R8904 VPWR.n349 VPWR.n348 7.99054
R8905 VPWR.n354 VPWR.n353 7.99054
R8906 VPWR.n359 VPWR.n358 7.99054
R8907 VPWR.n364 VPWR.n363 7.99054
R8908 VPWR VPWR.n1980 7.89251
R8909 VPWR VPWR.n156 7.89251
R8910 VPWR VPWR.n116 7.89251
R8911 VPWR VPWR.n76 7.89251
R8912 VPWR VPWR.n29 7.89251
R8913 VPWR.n1982 VPWR.n1981 7.87003
R8914 VPWR.n1984 VPWR.n1983 7.87003
R8915 VPWR.n1986 VPWR.n1985 7.87003
R8916 VPWR.n1988 VPWR.n1987 7.87003
R8917 VPWR.n1990 VPWR.n1989 7.87003
R8918 VPWR.n1992 VPWR.n1991 7.87003
R8919 VPWR.n1995 VPWR.n1994 7.87003
R8920 VPWR.n1997 VPWR.n1996 7.87003
R8921 VPWR.n1999 VPWR.n1998 7.87003
R8922 VPWR.n158 VPWR.n157 7.87003
R8923 VPWR.n160 VPWR.n159 7.87003
R8924 VPWR.n162 VPWR.n161 7.87003
R8925 VPWR.n164 VPWR.n163 7.87003
R8926 VPWR.n166 VPWR.n165 7.87003
R8927 VPWR.n168 VPWR.n167 7.87003
R8928 VPWR.n170 VPWR.n169 7.87003
R8929 VPWR.n118 VPWR.n117 7.87003
R8930 VPWR.n120 VPWR.n119 7.87003
R8931 VPWR.n122 VPWR.n121 7.87003
R8932 VPWR.n124 VPWR.n123 7.87003
R8933 VPWR.n126 VPWR.n125 7.87003
R8934 VPWR.n128 VPWR.n127 7.87003
R8935 VPWR.n130 VPWR.n129 7.87003
R8936 VPWR.n78 VPWR.n77 7.87003
R8937 VPWR.n80 VPWR.n79 7.87003
R8938 VPWR.n82 VPWR.n81 7.87003
R8939 VPWR.n84 VPWR.n83 7.87003
R8940 VPWR.n86 VPWR.n85 7.87003
R8941 VPWR.n88 VPWR.n87 7.87003
R8942 VPWR.n90 VPWR.n89 7.87003
R8943 VPWR.n1213 VPWR.n1212 7.87003
R8944 VPWR.n1215 VPWR.n1214 7.87003
R8945 VPWR.n1217 VPWR.n1216 7.87003
R8946 VPWR.n1219 VPWR.n1218 7.87003
R8947 VPWR.n1221 VPWR.n1220 7.87003
R8948 VPWR.n1223 VPWR.n1222 7.87003
R8949 VPWR.n1225 VPWR.n1224 7.87003
R8950 VPWR.n1228 VPWR.n1227 7.87003
R8951 VPWR.n1230 VPWR.n1229 7.87003
R8952 VPWR.n1232 VPWR.n1231 7.87003
R8953 VPWR.n1234 VPWR.n1233 7.87003
R8954 VPWR.n1236 VPWR.n1235 7.87003
R8955 VPWR.n1238 VPWR.n1237 7.87003
R8956 VPWR.n1514 VPWR.n1513 7.87003
R8957 VPWR.n1516 VPWR.n1515 7.87003
R8958 VPWR.n1518 VPWR.n1517 7.87003
R8959 VPWR.n1520 VPWR.n1519 7.87003
R8960 VPWR.n1522 VPWR.n1521 7.87003
R8961 VPWR.n1544 VPWR.n1543 7.87003
R8962 VPWR.n1546 VPWR.n1545 7.87003
R8963 VPWR.n1549 VPWR.n1548 7.87003
R8964 VPWR.n1552 VPWR.n1551 7.87003
R8965 VPWR.n1555 VPWR.n1554 7.87003
R8966 VPWR.n1557 VPWR.n1556 7.87003
R8967 VPWR.n1560 VPWR.n1559 7.87003
R8968 VPWR.n1562 VPWR.n1561 7.87003
R8969 VPWR.n1564 VPWR.n1563 7.87003
R8970 VPWR.n1567 VPWR.n1566 7.87003
R8971 VPWR.n1569 VPWR.n1568 7.87003
R8972 VPWR.n1571 VPWR.n1570 7.87003
R8973 VPWR.n1574 VPWR.n1573 7.87003
R8974 VPWR.n1577 VPWR.n1576 7.87003
R8975 VPWR.n1580 VPWR.n1579 7.87003
R8976 VPWR.n1602 VPWR.n1601 7.87003
R8977 VPWR.n746 VPWR.n745 7.87003
R8978 VPWR.n748 VPWR.n747 7.87003
R8979 VPWR.n750 VPWR.n749 7.87003
R8980 VPWR.n752 VPWR.n751 7.87003
R8981 VPWR.n754 VPWR.n753 7.87003
R8982 VPWR.n756 VPWR.n755 7.87003
R8983 VPWR.n758 VPWR.n757 7.87003
R8984 VPWR.n761 VPWR.n760 7.87003
R8985 VPWR.n763 VPWR.n762 7.87003
R8986 VPWR.n765 VPWR.n764 7.87003
R8987 VPWR.n767 VPWR.n766 7.87003
R8988 VPWR.n769 VPWR.n768 7.87003
R8989 VPWR.n771 VPWR.n770 7.87003
R8990 VPWR.n292 VPWR.n291 7.87003
R8991 VPWR.n294 VPWR.n293 7.87003
R8992 VPWR.n296 VPWR.n295 7.87003
R8993 VPWR.n298 VPWR.n297 7.87003
R8994 VPWR.n300 VPWR.n299 7.87003
R8995 VPWR.n302 VPWR.n301 7.87003
R8996 VPWR.n304 VPWR.n303 7.87003
R8997 VPWR.n307 VPWR.n306 7.87003
R8998 VPWR.n309 VPWR.n308 7.87003
R8999 VPWR.n311 VPWR.n310 7.87003
R9000 VPWR.n313 VPWR.n312 7.87003
R9001 VPWR.n315 VPWR.n314 7.87003
R9002 VPWR.n317 VPWR.n316 7.87003
R9003 VPWR.n416 VPWR.n415 7.87003
R9004 VPWR.n418 VPWR.n417 7.87003
R9005 VPWR.n420 VPWR.n419 7.87003
R9006 VPWR.n422 VPWR.n421 7.87003
R9007 VPWR.n424 VPWR.n423 7.87003
R9008 VPWR.n426 VPWR.n425 7.87003
R9009 VPWR.n428 VPWR.n427 7.87003
R9010 VPWR.n431 VPWR.n430 7.87003
R9011 VPWR.n433 VPWR.n432 7.87003
R9012 VPWR.n435 VPWR.n434 7.87003
R9013 VPWR.n437 VPWR.n436 7.87003
R9014 VPWR.n439 VPWR.n438 7.87003
R9015 VPWR.n441 VPWR.n440 7.87003
R9016 VPWR.n1110 VPWR.n1109 7.87003
R9017 VPWR.n1124 VPWR.n1115 7.87003
R9018 VPWR.n1123 VPWR.n1116 7.87003
R9019 VPWR.n1122 VPWR.n1119 7.87003
R9020 VPWR.n1121 VPWR.n1120 7.87003
R9021 VPWR.n31 VPWR.n30 7.87003
R9022 VPWR.n33 VPWR.n32 7.87003
R9023 VPWR.n35 VPWR.n34 7.87003
R9024 VPWR.n37 VPWR.n36 7.87003
R9025 VPWR.n39 VPWR.n38 7.87003
R9026 VPWR.n41 VPWR.n40 7.87003
R9027 VPWR.n43 VPWR.n42 7.87003
R9028 VPWR VPWR.n2025 7.82272
R9029 VPWR.n2028 VPWR 7.82272
R9030 VPWR.n2027 VPWR 7.82272
R9031 VPWR VPWR.n2036 7.82272
R9032 VPWR.n2037 VPWR 7.82272
R9033 VPWR VPWR.n2046 7.82272
R9034 VPWR.n2047 VPWR 7.82272
R9035 VPWR VPWR.n2054 7.82272
R9036 VPWR VPWR.n2055 7.82272
R9037 VPWR.n2056 VPWR 7.82272
R9038 VPWR VPWR.n2065 7.82272
R9039 VPWR.n2131 VPWR 7.82272
R9040 VPWR.n2128 VPWR 7.82272
R9041 VPWR.n2124 VPWR 7.82272
R9042 VPWR.n2123 VPWR 7.82272
R9043 VPWR.n2119 VPWR 7.82272
R9044 VPWR.n2115 VPWR 7.82272
R9045 VPWR.n2112 VPWR 7.82272
R9046 VPWR.n2108 VPWR 7.82272
R9047 VPWR.n2107 VPWR 7.82272
R9048 VPWR.n2103 VPWR 7.82272
R9049 VPWR.n2099 VPWR 7.82272
R9050 VPWR.n2197 VPWR 7.82272
R9051 VPWR.n2194 VPWR 7.82272
R9052 VPWR.n2190 VPWR 7.82272
R9053 VPWR.n2189 VPWR 7.82272
R9054 VPWR.n2185 VPWR 7.82272
R9055 VPWR.n2181 VPWR 7.82272
R9056 VPWR.n2178 VPWR 7.82272
R9057 VPWR.n2174 VPWR 7.82272
R9058 VPWR.n2173 VPWR 7.82272
R9059 VPWR.n2169 VPWR 7.82272
R9060 VPWR.n2165 VPWR 7.82272
R9061 VPWR.n2263 VPWR 7.82272
R9062 VPWR.n2260 VPWR 7.82272
R9063 VPWR.n2256 VPWR 7.82272
R9064 VPWR.n2255 VPWR 7.82272
R9065 VPWR.n2251 VPWR 7.82272
R9066 VPWR.n2247 VPWR 7.82272
R9067 VPWR.n2244 VPWR 7.82272
R9068 VPWR.n2240 VPWR 7.82272
R9069 VPWR.n2239 VPWR 7.82272
R9070 VPWR.n2235 VPWR 7.82272
R9071 VPWR.n2231 VPWR 7.82272
R9072 VPWR VPWR.n1179 7.82272
R9073 VPWR.n1317 VPWR 7.82272
R9074 VPWR VPWR.n1320 7.82272
R9075 VPWR VPWR.n1324 7.82272
R9076 VPWR VPWR.n1328 7.82272
R9077 VPWR.n1329 VPWR 7.82272
R9078 VPWR.n1333 VPWR 7.82272
R9079 VPWR.n1337 VPWR 7.82272
R9080 VPWR.n1341 VPWR 7.82272
R9081 VPWR VPWR.n1344 7.82272
R9082 VPWR.n1345 VPWR 7.82272
R9083 VPWR VPWR.n1348 7.82272
R9084 VPWR VPWR.n1352 7.82272
R9085 VPWR.n1353 VPWR 7.82272
R9086 VPWR VPWR.n1356 7.82272
R9087 VPWR.n1357 VPWR 7.82272
R9088 VPWR.n1361 VPWR 7.82272
R9089 VPWR VPWR.n1364 7.82272
R9090 VPWR.n1365 VPWR 7.82272
R9091 VPWR VPWR.n1368 7.82272
R9092 VPWR VPWR.n1372 7.82272
R9093 VPWR.n1373 VPWR 7.82272
R9094 VPWR VPWR.n1376 7.82272
R9095 VPWR.n1377 VPWR 7.82272
R9096 VPWR.n1381 VPWR 7.82272
R9097 VPWR VPWR.n1384 7.82272
R9098 VPWR.n1385 VPWR 7.82272
R9099 VPWR VPWR.n1388 7.82272
R9100 VPWR VPWR.n1392 7.82272
R9101 VPWR.n1393 VPWR 7.82272
R9102 VPWR VPWR.n1396 7.82272
R9103 VPWR VPWR.n1400 7.82272
R9104 VPWR.n1401 VPWR 7.82272
R9105 VPWR VPWR.n1404 7.82272
R9106 VPWR VPWR.n1408 7.82272
R9107 VPWR VPWR.n1412 7.82272
R9108 VPWR VPWR.n1416 7.82272
R9109 VPWR VPWR.n1420 7.82272
R9110 VPWR VPWR.n1424 7.82272
R9111 VPWR VPWR.n1455 7.82272
R9112 VPWR.n1715 VPWR 7.82272
R9113 VPWR.n1714 VPWR 7.82272
R9114 VPWR.n1708 VPWR 7.82272
R9115 VPWR.n1707 VPWR 7.82272
R9116 VPWR VPWR.n1462 7.82272
R9117 VPWR.n1699 VPWR 7.82272
R9118 VPWR.n1698 VPWR 7.82272
R9119 VPWR VPWR.n1469 7.82272
R9120 VPWR.n1692 VPWR 7.82272
R9121 VPWR.n1691 VPWR 7.82272
R9122 VPWR.n1690 VPWR 7.82272
R9123 VPWR VPWR.n1474 7.82272
R9124 VPWR.n1683 VPWR 7.82272
R9125 VPWR.n1682 VPWR 7.82272
R9126 VPWR VPWR.n1477 7.82272
R9127 VPWR.n1676 VPWR 7.82272
R9128 VPWR.n1675 VPWR 7.82272
R9129 VPWR.n1674 VPWR 7.82272
R9130 VPWR VPWR.n1482 7.82272
R9131 VPWR.n1667 VPWR 7.82272
R9132 VPWR.n1666 VPWR 7.82272
R9133 VPWR VPWR.n1485 7.82272
R9134 VPWR.n1660 VPWR 7.82272
R9135 VPWR.n1658 VPWR 7.82272
R9136 VPWR VPWR.n1489 7.82272
R9137 VPWR.n1652 VPWR 7.82272
R9138 VPWR.n1651 VPWR 7.82272
R9139 VPWR VPWR.n1490 7.82272
R9140 VPWR.n1644 VPWR 7.82272
R9141 VPWR.n1643 VPWR 7.82272
R9142 VPWR.n1642 VPWR 7.82272
R9143 VPWR VPWR.n1497 7.82272
R9144 VPWR.n1636 VPWR 7.82272
R9145 VPWR.n1635 VPWR 7.82272
R9146 VPWR VPWR.n1498 7.82272
R9147 VPWR.n1628 VPWR 7.82272
R9148 VPWR.n1627 VPWR 7.82272
R9149 VPWR.n1626 VPWR 7.82272
R9150 VPWR VPWR.n1505 7.82272
R9151 VPWR.n1620 VPWR 7.82272
R9152 VPWR.n1619 VPWR 7.82272
R9153 VPWR.n814 VPWR 7.82272
R9154 VPWR.n818 VPWR 7.82272
R9155 VPWR VPWR.n821 7.82272
R9156 VPWR VPWR.n825 7.82272
R9157 VPWR VPWR.n829 7.82272
R9158 VPWR.n830 VPWR 7.82272
R9159 VPWR.n834 VPWR 7.82272
R9160 VPWR.n838 VPWR 7.82272
R9161 VPWR.n842 VPWR 7.82272
R9162 VPWR VPWR.n845 7.82272
R9163 VPWR.n846 VPWR 7.82272
R9164 VPWR VPWR.n849 7.82272
R9165 VPWR VPWR.n853 7.82272
R9166 VPWR.n854 VPWR 7.82272
R9167 VPWR VPWR.n857 7.82272
R9168 VPWR.n858 VPWR 7.82272
R9169 VPWR.n862 VPWR 7.82272
R9170 VPWR VPWR.n865 7.82272
R9171 VPWR.n866 VPWR 7.82272
R9172 VPWR VPWR.n869 7.82272
R9173 VPWR VPWR.n873 7.82272
R9174 VPWR.n874 VPWR 7.82272
R9175 VPWR VPWR.n877 7.82272
R9176 VPWR.n878 VPWR 7.82272
R9177 VPWR.n882 VPWR 7.82272
R9178 VPWR VPWR.n885 7.82272
R9179 VPWR.n886 VPWR 7.82272
R9180 VPWR VPWR.n889 7.82272
R9181 VPWR VPWR.n893 7.82272
R9182 VPWR.n894 VPWR 7.82272
R9183 VPWR VPWR.n897 7.82272
R9184 VPWR VPWR.n901 7.82272
R9185 VPWR.n902 VPWR 7.82272
R9186 VPWR VPWR.n905 7.82272
R9187 VPWR VPWR.n909 7.82272
R9188 VPWR VPWR.n913 7.82272
R9189 VPWR VPWR.n917 7.82272
R9190 VPWR VPWR.n921 7.82272
R9191 VPWR VPWR.n924 7.82272
R9192 VPWR VPWR.n258 7.82272
R9193 VPWR.n1782 VPWR 7.82272
R9194 VPWR VPWR.n1785 7.82272
R9195 VPWR VPWR.n1789 7.82272
R9196 VPWR VPWR.n1793 7.82272
R9197 VPWR.n1794 VPWR 7.82272
R9198 VPWR.n1798 VPWR 7.82272
R9199 VPWR.n1802 VPWR 7.82272
R9200 VPWR.n1806 VPWR 7.82272
R9201 VPWR VPWR.n1809 7.82272
R9202 VPWR.n1810 VPWR 7.82272
R9203 VPWR VPWR.n1813 7.82272
R9204 VPWR VPWR.n1817 7.82272
R9205 VPWR.n1818 VPWR 7.82272
R9206 VPWR VPWR.n1821 7.82272
R9207 VPWR.n1822 VPWR 7.82272
R9208 VPWR.n1826 VPWR 7.82272
R9209 VPWR VPWR.n1829 7.82272
R9210 VPWR.n1830 VPWR 7.82272
R9211 VPWR VPWR.n1833 7.82272
R9212 VPWR VPWR.n1837 7.82272
R9213 VPWR.n1838 VPWR 7.82272
R9214 VPWR VPWR.n1841 7.82272
R9215 VPWR.n1842 VPWR 7.82272
R9216 VPWR.n1846 VPWR 7.82272
R9217 VPWR VPWR.n1849 7.82272
R9218 VPWR.n1850 VPWR 7.82272
R9219 VPWR VPWR.n1853 7.82272
R9220 VPWR VPWR.n1857 7.82272
R9221 VPWR.n1858 VPWR 7.82272
R9222 VPWR VPWR.n1861 7.82272
R9223 VPWR VPWR.n1865 7.82272
R9224 VPWR.n1866 VPWR 7.82272
R9225 VPWR VPWR.n1869 7.82272
R9226 VPWR VPWR.n1873 7.82272
R9227 VPWR VPWR.n1877 7.82272
R9228 VPWR VPWR.n1881 7.82272
R9229 VPWR VPWR.n1885 7.82272
R9230 VPWR VPWR.n1889 7.82272
R9231 VPWR VPWR.n1920 7.82272
R9232 VPWR.n1931 VPWR 7.82272
R9233 VPWR VPWR.n1924 7.82272
R9234 VPWR.n484 VPWR 7.82272
R9235 VPWR.n488 VPWR 7.82272
R9236 VPWR VPWR.n491 7.82272
R9237 VPWR VPWR.n495 7.82272
R9238 VPWR VPWR.n499 7.82272
R9239 VPWR.n500 VPWR 7.82272
R9240 VPWR.n504 VPWR 7.82272
R9241 VPWR.n508 VPWR 7.82272
R9242 VPWR.n512 VPWR 7.82272
R9243 VPWR VPWR.n515 7.82272
R9244 VPWR.n516 VPWR 7.82272
R9245 VPWR VPWR.n519 7.82272
R9246 VPWR VPWR.n523 7.82272
R9247 VPWR.n524 VPWR 7.82272
R9248 VPWR VPWR.n527 7.82272
R9249 VPWR.n528 VPWR 7.82272
R9250 VPWR.n532 VPWR 7.82272
R9251 VPWR VPWR.n535 7.82272
R9252 VPWR.n536 VPWR 7.82272
R9253 VPWR VPWR.n539 7.82272
R9254 VPWR VPWR.n543 7.82272
R9255 VPWR.n544 VPWR 7.82272
R9256 VPWR VPWR.n547 7.82272
R9257 VPWR.n548 VPWR 7.82272
R9258 VPWR.n552 VPWR 7.82272
R9259 VPWR VPWR.n555 7.82272
R9260 VPWR.n556 VPWR 7.82272
R9261 VPWR VPWR.n559 7.82272
R9262 VPWR VPWR.n563 7.82272
R9263 VPWR.n564 VPWR 7.82272
R9264 VPWR VPWR.n567 7.82272
R9265 VPWR VPWR.n571 7.82272
R9266 VPWR.n572 VPWR 7.82272
R9267 VPWR VPWR.n575 7.82272
R9268 VPWR VPWR.n579 7.82272
R9269 VPWR VPWR.n583 7.82272
R9270 VPWR VPWR.n587 7.82272
R9271 VPWR VPWR.n591 7.82272
R9272 VPWR VPWR.n594 7.82272
R9273 VPWR.n1096 VPWR 7.82272
R9274 VPWR VPWR.n1138 7.82272
R9275 VPWR.n1141 VPWR 7.82272
R9276 VPWR.n1140 VPWR 7.82272
R9277 VPWR VPWR.n1149 7.82272
R9278 VPWR.n1151 VPWR 7.82272
R9279 VPWR.n1150 VPWR 7.82272
R9280 VPWR VPWR.n1159 7.82272
R9281 VPWR.n1000 VPWR 7.82272
R9282 VPWR VPWR.n1036 7.82272
R9283 VPWR.n1039 VPWR 7.82272
R9284 VPWR.n1038 VPWR 7.82272
R9285 VPWR VPWR.n1047 7.82272
R9286 VPWR.n1049 VPWR 7.82272
R9287 VPWR.n1048 VPWR 7.82272
R9288 VPWR VPWR.n1057 7.82272
R9289 VPWR.n2329 VPWR 7.82272
R9290 VPWR.n2326 VPWR 7.82272
R9291 VPWR.n2322 VPWR 7.82272
R9292 VPWR.n2321 VPWR 7.82272
R9293 VPWR.n2317 VPWR 7.82272
R9294 VPWR.n2313 VPWR 7.82272
R9295 VPWR.n2310 VPWR 7.82272
R9296 VPWR.n2306 VPWR 7.82272
R9297 VPWR.n2305 VPWR 7.82272
R9298 VPWR.n2301 VPWR 7.82272
R9299 VPWR.n2297 VPWR 7.82272
R9300 VPWR.n2003 VPWR 7.52991
R9301 VPWR.n2001 VPWR 7.52991
R9302 VPWR.n174 VPWR 7.52991
R9303 VPWR.n172 VPWR 7.52991
R9304 VPWR.n134 VPWR 7.52991
R9305 VPWR.n132 VPWR 7.52991
R9306 VPWR.n94 VPWR 7.52991
R9307 VPWR.n92 VPWR 7.52991
R9308 VPWR.n1177 VPWR 7.52991
R9309 VPWR.n1244 VPWR 7.52991
R9310 VPWR.n1240 VPWR 7.52991
R9311 VPWR.n1437 VPWR 7.52991
R9312 VPWR.n1453 VPWR 7.52991
R9313 VPWR.n1608 VPWR 7.52991
R9314 VPWR.n1604 VPWR 7.52991
R9315 VPWR.n1726 VPWR 7.52991
R9316 VPWR.n744 VPWR 7.52991
R9317 VPWR.n724 VPWR 7.52991
R9318 VPWR.n956 VPWR 7.52991
R9319 VPWR.n773 VPWR 7.52991
R9320 VPWR.n256 VPWR 7.52991
R9321 VPWR.n323 VPWR 7.52991
R9322 VPWR.n319 VPWR 7.52991
R9323 VPWR.n1902 VPWR 7.52991
R9324 VPWR.n1918 VPWR.n1917 7.52991
R9325 VPWR.n1915 VPWR 7.52991
R9326 VPWR.n1944 VPWR.n1942 7.52991
R9327 VPWR.n1914 VPWR 7.52991
R9328 VPWR.n1947 VPWR 7.52991
R9329 VPWR.n1952 VPWR 7.52991
R9330 VPWR.n1957 VPWR 7.52991
R9331 VPWR.n414 VPWR 7.52991
R9332 VPWR.n394 VPWR 7.52991
R9333 VPWR.n626 VPWR 7.52991
R9334 VPWR.n443 VPWR 7.52991
R9335 VPWR.n1092 VPWR 7.52991
R9336 VPWR.n1070 VPWR 7.52991
R9337 VPWR.n1072 VPWR 7.52991
R9338 VPWR.n1126 VPWR 7.52991
R9339 VPWR.n1112 VPWR 7.52991
R9340 VPWR.n1091 VPWR 7.52991
R9341 VPWR.n47 VPWR 7.52991
R9342 VPWR.n45 VPWR 7.52991
R9343 VPWR.n1979 VPWR.n1978 7.23528
R9344 VPWR.n195 VPWR.n155 7.23528
R9345 VPWR.n690 VPWR.n154 7.23528
R9346 VPWR.n691 VPWR.n115 7.23528
R9347 VPWR.n638 VPWR.n75 7.23528
R9348 VPWR.n74 VPWR.n28 7.23528
R9349 VPWR.n373 VPWR.n370 7.03865
R9350 VPWR.n373 VPWR.n369 7.03865
R9351 VPWR.n378 VPWR.n375 7.03865
R9352 VPWR.n378 VPWR.n374 7.03865
R9353 VPWR.n383 VPWR.n380 7.03865
R9354 VPWR.n383 VPWR.n379 7.03865
R9355 VPWR.n388 VPWR.n385 7.03865
R9356 VPWR.n388 VPWR.n384 7.03865
R9357 VPWR.n7 VPWR.n4 7.03865
R9358 VPWR.n7 VPWR.n3 7.03865
R9359 VPWR.n12 VPWR.n9 7.03865
R9360 VPWR.n12 VPWR.n8 7.03865
R9361 VPWR.n17 VPWR.n14 7.03865
R9362 VPWR.n17 VPWR.n13 7.03865
R9363 VPWR.n22 VPWR.n19 7.03865
R9364 VPWR.n22 VPWR.n18 7.03865
R9365 VPWR.n703 VPWR.n700 7.03865
R9366 VPWR.n703 VPWR.n699 7.03865
R9367 VPWR.n708 VPWR.n705 7.03865
R9368 VPWR.n708 VPWR.n704 7.03865
R9369 VPWR.n713 VPWR.n710 7.03865
R9370 VPWR.n713 VPWR.n709 7.03865
R9371 VPWR.n718 VPWR.n715 7.03865
R9372 VPWR.n718 VPWR.n714 7.03865
R9373 VPWR.n234 VPWR.n231 7.03865
R9374 VPWR.n234 VPWR.n230 7.03865
R9375 VPWR.n239 VPWR.n236 7.03865
R9376 VPWR.n239 VPWR.n235 7.03865
R9377 VPWR.n244 VPWR.n241 7.03865
R9378 VPWR.n244 VPWR.n240 7.03865
R9379 VPWR.n249 VPWR.n246 7.03865
R9380 VPWR.n249 VPWR.n245 7.03865
R9381 VPWR.n2005 VPWR.n2002 6.77697
R9382 VPWR.n2075 VPWR.n2074 6.77697
R9383 VPWR.n176 VPWR.n173 6.77697
R9384 VPWR.n2140 VPWR.n2139 6.77697
R9385 VPWR.n136 VPWR.n133 6.77697
R9386 VPWR.n2206 VPWR.n2205 6.77697
R9387 VPWR.n96 VPWR.n93 6.77697
R9388 VPWR.n2272 VPWR.n2271 6.77697
R9389 VPWR.n1442 VPWR.n1441 6.77697
R9390 VPWR.n1246 VPWR.n1211 6.77697
R9391 VPWR.n1239 VPWR.n1210 6.77697
R9392 VPWR.n1439 VPWR.n1436 6.77697
R9393 VPWR.n1731 VPWR.n1730 6.77697
R9394 VPWR.n1610 VPWR.n1510 6.77697
R9395 VPWR.n1603 VPWR.n1509 6.77697
R9396 VPWR.n1728 VPWR.n1725 6.77697
R9397 VPWR.n778 VPWR.n743 6.77697
R9398 VPWR.n961 VPWR.n960 6.77697
R9399 VPWR.n958 VPWR.n955 6.77697
R9400 VPWR.n772 VPWR.n742 6.77697
R9401 VPWR.n1907 VPWR.n1906 6.77697
R9402 VPWR.n325 VPWR.n290 6.77697
R9403 VPWR.n318 VPWR.n289 6.77697
R9404 VPWR.n1904 VPWR.n1901 6.77697
R9405 VPWR.n1917 VPWR.n1916 6.77697
R9406 VPWR.n1944 VPWR.n1943 6.77697
R9407 VPWR.n1949 VPWR.n1948 6.77697
R9408 VPWR.n1954 VPWR.n1953 6.77697
R9409 VPWR.n1959 VPWR.n1958 6.77697
R9410 VPWR.n448 VPWR.n413 6.77697
R9411 VPWR.n631 VPWR.n630 6.77697
R9412 VPWR.n628 VPWR.n625 6.77697
R9413 VPWR.n442 VPWR.n412 6.77697
R9414 VPWR.n1094 VPWR.n1093 6.77697
R9415 VPWR.n1169 VPWR.n1168 6.77697
R9416 VPWR.n1074 VPWR.n1071 6.77697
R9417 VPWR.n1128 VPWR.n1089 6.77697
R9418 VPWR.n1111 VPWR.n1088 6.77697
R9419 VPWR.n1106 VPWR.n1105 6.77697
R9420 VPWR.n49 VPWR.n46 6.77697
R9421 VPWR.n2338 VPWR.n2337 6.77697
R9422 VPWR.n373 VPWR.n372 6.51659
R9423 VPWR.n378 VPWR.n377 6.51659
R9424 VPWR.n383 VPWR.n382 6.51659
R9425 VPWR.n388 VPWR.n387 6.51659
R9426 VPWR.n7 VPWR.n6 6.51659
R9427 VPWR.n12 VPWR.n11 6.51659
R9428 VPWR.n17 VPWR.n16 6.51659
R9429 VPWR.n22 VPWR.n21 6.51659
R9430 VPWR.n703 VPWR.n702 6.51659
R9431 VPWR.n708 VPWR.n707 6.51659
R9432 VPWR.n713 VPWR.n712 6.51659
R9433 VPWR.n718 VPWR.n717 6.51659
R9434 VPWR.n234 VPWR.n233 6.51659
R9435 VPWR.n239 VPWR.n238 6.51659
R9436 VPWR.n244 VPWR.n243 6.51659
R9437 VPWR.n249 VPWR.n248 6.51659
R9438 VPWR.n1173 VPWR 6.4005
R9439 VPWR.n2345 VPWR 6.02075
R9440 VPWR.n2346 VPWR 5.97326
R9441 VPWR.n1543 VPWR.n1542 5.39616
R9442 VPWR.n1601 VPWR.n1600 5.39616
R9443 VPWR.n2071 VPWR.n2006 5.21532
R9444 VPWR.n2136 VPWR.n2083 5.21532
R9445 VPWR.n2202 VPWR.n2149 5.21532
R9446 VPWR.n2268 VPWR.n2215 5.21532
R9447 VPWR.n1428 VPWR.n1427 5.21532
R9448 VPWR.n1613 VPWR.n1506 5.21532
R9449 VPWR.n930 VPWR.n781 5.21532
R9450 VPWR.n1893 VPWR.n1892 5.21532
R9451 VPWR.n600 VPWR.n451 5.21532
R9452 VPWR.n1132 VPWR.n1131 5.21532
R9453 VPWR.n1165 VPWR.n1075 5.21532
R9454 VPWR.n1030 VPWR.n1029 5.21532
R9455 VPWR.n1063 VPWR.n985 5.21532
R9456 VPWR.n2334 VPWR.n2281 5.21532
R9457 VPWR.n1249 VPWR.n339 4.67341
R9458 VPWR.n74 VPWR.n73 4.6505
R9459 VPWR.n693 VPWR.n691 4.6505
R9460 VPWR.n683 VPWR.n154 4.6505
R9461 VPWR.n226 VPWR.n195 4.6505
R9462 VPWR.n1979 VPWR.n194 4.6505
R9463 VPWR.n67 VPWR.n28 4.6505
R9464 VPWR.n692 VPWR.n115 4.6505
R9465 VPWR.n690 VPWR.n689 4.6505
R9466 VPWR.n225 VPWR.n155 4.6505
R9467 VPWR.n1978 VPWR.n1977 4.6505
R9468 VPWR.n639 VPWR.n75 4.6505
R9469 VPWR.n640 VPWR.n638 4.6505
R9470 VPWR.n1451 VPWR.n982 4.6334
R9471 VPWR.n1451 VPWR.n981 4.6334
R9472 VPWR.n1451 VPWR.n980 4.6334
R9473 VPWR.n1451 VPWR.n330 4.6334
R9474 VPWR.n1736 VPWR.n331 4.6334
R9475 VPWR.n1946 VPWR.n1913 3.95786
R9476 VPWR.n1108 VPWR.n1090 3.95489
R9477 VPWR.n1961 VPWR.n1960 3.9165
R9478 VPWR.n1956 VPWR.n1955 3.9165
R9479 VPWR.n1951 VPWR.n1950 3.9165
R9480 VPWR.n1946 VPWR.n1945 3.9165
R9481 VPWR.n2077 VPWR.n2076 3.90993
R9482 VPWR.n2004 VPWR.n2000 3.90993
R9483 VPWR.n2142 VPWR.n2141 3.90993
R9484 VPWR.n175 VPWR.n171 3.90993
R9485 VPWR.n2208 VPWR.n2207 3.90993
R9486 VPWR.n135 VPWR.n131 3.90993
R9487 VPWR.n2274 VPWR.n2273 3.90993
R9488 VPWR.n95 VPWR.n91 3.90993
R9489 VPWR.n1438 VPWR.n1176 3.90993
R9490 VPWR.n1727 VPWR.n1452 3.90993
R9491 VPWR.n1606 VPWR.n1605 3.90993
R9492 VPWR.n1609 VPWR.n1607 3.90993
R9493 VPWR.n1733 VPWR.n1732 3.90993
R9494 VPWR.n777 VPWR.n776 3.90993
R9495 VPWR.n957 VPWR.n723 3.90993
R9496 VPWR.n963 VPWR.n962 3.90993
R9497 VPWR.n775 VPWR.n774 3.90993
R9498 VPWR.n1903 VPWR.n255 3.90993
R9499 VPWR.n321 VPWR.n320 3.90993
R9500 VPWR.n324 VPWR.n322 3.90993
R9501 VPWR.n1909 VPWR.n1908 3.90993
R9502 VPWR.n447 VPWR.n446 3.90993
R9503 VPWR.n627 VPWR.n393 3.90993
R9504 VPWR.n633 VPWR.n632 3.90993
R9505 VPWR.n445 VPWR.n444 3.90993
R9506 VPWR.n1108 VPWR.n1107 3.90993
R9507 VPWR.n1114 VPWR.n1113 3.90993
R9508 VPWR.n1127 VPWR.n1125 3.90993
R9509 VPWR.n1073 VPWR.n1069 3.90993
R9510 VPWR.n1171 VPWR.n1170 3.90993
R9511 VPWR.n1242 VPWR.n1241 3.90993
R9512 VPWR.n1245 VPWR.n1243 3.90993
R9513 VPWR.n1444 VPWR.n1443 3.90993
R9514 VPWR.n2340 VPWR.n2339 3.90993
R9515 VPWR.n48 VPWR.n44 3.90993
R9516 VPWR.n1172 VPWR 3.62284
R9517 VPWR.n1068 VPWR 3.62284
R9518 VPWR.n2143 VPWR 3.45629
R9519 VPWR.n2209 VPWR 3.45629
R9520 VPWR.n2275 VPWR 3.45629
R9521 VPWR.n2341 VPWR 3.45629
R9522 VPWR VPWR.n2078 3.45604
R9523 VPWR VPWR.n2144 3.45604
R9524 VPWR VPWR.n2210 3.45604
R9525 VPWR VPWR.n2276 3.45604
R9526 VPWR.n970 VPWR.n654 3.4105
R9527 VPWR.n971 VPWR.n970 3.4105
R9528 VPWR.n694 VPWR.n681 3.4105
R9529 VPWR.n682 VPWR.n681 3.4105
R9530 VPWR.n1975 VPWR.n197 3.4105
R9531 VPWR.n1976 VPWR.n1975 3.4105
R9532 VPWR.n1738 VPWR.n328 3.4105
R9533 VPWR.n329 VPWR.n328 3.4105
R9534 VPWR.n975 VPWR.n974 3.4105
R9535 VPWR.n976 VPWR.n975 3.4105
R9536 VPWR.n227 VPWR.n223 3.4105
R9537 VPWR.n224 VPWR.n223 3.4105
R9538 VPWR.n687 VPWR.n685 3.4105
R9539 VPWR.n688 VPWR.n687 3.4105
R9540 VPWR.n649 VPWR.n342 3.4105
R9541 VPWR.n650 VPWR.n649 3.4105
R9542 VPWR.n1449 VPWR.n1448 3.4105
R9543 VPWR.n1448 VPWR.n1447 3.4105
R9544 VPWR.n72 VPWR.n71 3.4105
R9545 VPWR.n71 VPWR.n70 3.4105
R9546 VPWR.n641 VPWR.n636 3.4105
R9547 VPWR.n637 VPWR.n636 3.4105
R9548 VPWR.n344 VPWR.n114 3.32807
R9549 VPWR.n2343 VPWR.n2342 3.31376
R9550 VPWR VPWR.n2019 2.60791
R9551 VPWR.n2026 VPWR 2.60791
R9552 VPWR VPWR.n2027 2.60791
R9553 VPWR.n2035 VPWR 2.60791
R9554 VPWR.n2038 VPWR 2.60791
R9555 VPWR.n2045 VPWR 2.60791
R9556 VPWR.n2047 VPWR 2.60791
R9557 VPWR VPWR.n2011 2.60791
R9558 VPWR.n2055 VPWR 2.60791
R9559 VPWR.n2057 VPWR 2.60791
R9560 VPWR.n2064 VPWR 2.60791
R9561 VPWR.n2066 VPWR 2.60791
R9562 VPWR.n2071 VPWR 2.60791
R9563 VPWR VPWR.n2132 2.60791
R9564 VPWR.n2128 VPWR 2.60791
R9565 VPWR VPWR.n2127 2.60791
R9566 VPWR VPWR.n2123 2.60791
R9567 VPWR.n2120 VPWR 2.60791
R9568 VPWR.n2116 VPWR 2.60791
R9569 VPWR.n2112 VPWR 2.60791
R9570 VPWR VPWR.n2111 2.60791
R9571 VPWR VPWR.n2107 2.60791
R9572 VPWR.n2104 VPWR 2.60791
R9573 VPWR.n2100 VPWR 2.60791
R9574 VPWR.n2096 VPWR 2.60791
R9575 VPWR.n2136 VPWR 2.60791
R9576 VPWR VPWR.n2198 2.60791
R9577 VPWR.n2194 VPWR 2.60791
R9578 VPWR VPWR.n2193 2.60791
R9579 VPWR VPWR.n2189 2.60791
R9580 VPWR.n2186 VPWR 2.60791
R9581 VPWR.n2182 VPWR 2.60791
R9582 VPWR.n2178 VPWR 2.60791
R9583 VPWR VPWR.n2177 2.60791
R9584 VPWR VPWR.n2173 2.60791
R9585 VPWR.n2170 VPWR 2.60791
R9586 VPWR.n2166 VPWR 2.60791
R9587 VPWR.n2162 VPWR 2.60791
R9588 VPWR.n2202 VPWR 2.60791
R9589 VPWR VPWR.n2264 2.60791
R9590 VPWR.n2260 VPWR 2.60791
R9591 VPWR VPWR.n2259 2.60791
R9592 VPWR VPWR.n2255 2.60791
R9593 VPWR.n2252 VPWR 2.60791
R9594 VPWR.n2248 VPWR 2.60791
R9595 VPWR.n2244 VPWR 2.60791
R9596 VPWR VPWR.n2243 2.60791
R9597 VPWR VPWR.n2239 2.60791
R9598 VPWR.n2236 VPWR 2.60791
R9599 VPWR.n2232 VPWR 2.60791
R9600 VPWR.n2228 VPWR 2.60791
R9601 VPWR.n2268 VPWR 2.60791
R9602 VPWR.n1434 VPWR 2.60791
R9603 VPWR VPWR.n1433 2.60791
R9604 VPWR.n1316 VPWR 2.60791
R9605 VPWR.n1320 VPWR 2.60791
R9606 VPWR.n1321 VPWR 2.60791
R9607 VPWR.n1325 VPWR 2.60791
R9608 VPWR.n1329 VPWR 2.60791
R9609 VPWR.n1332 VPWR 2.60791
R9610 VPWR.n1336 VPWR 2.60791
R9611 VPWR.n1340 VPWR 2.60791
R9612 VPWR.n1344 VPWR 2.60791
R9613 VPWR.n1345 VPWR 2.60791
R9614 VPWR.n1348 VPWR 2.60791
R9615 VPWR.n1349 VPWR 2.60791
R9616 VPWR.n1353 VPWR 2.60791
R9617 VPWR.n1356 VPWR 2.60791
R9618 VPWR.n1357 VPWR 2.60791
R9619 VPWR.n1360 VPWR 2.60791
R9620 VPWR.n1364 VPWR 2.60791
R9621 VPWR.n1365 VPWR 2.60791
R9622 VPWR.n1368 VPWR 2.60791
R9623 VPWR.n1369 VPWR 2.60791
R9624 VPWR.n1373 VPWR 2.60791
R9625 VPWR.n1376 VPWR 2.60791
R9626 VPWR.n1377 VPWR 2.60791
R9627 VPWR.n1380 VPWR 2.60791
R9628 VPWR.n1384 VPWR 2.60791
R9629 VPWR.n1385 VPWR 2.60791
R9630 VPWR.n1388 VPWR 2.60791
R9631 VPWR.n1389 VPWR 2.60791
R9632 VPWR.n1393 VPWR 2.60791
R9633 VPWR.n1396 VPWR 2.60791
R9634 VPWR.n1397 VPWR 2.60791
R9635 VPWR.n1401 VPWR 2.60791
R9636 VPWR.n1404 VPWR 2.60791
R9637 VPWR.n1405 VPWR 2.60791
R9638 VPWR.n1409 VPWR 2.60791
R9639 VPWR.n1413 VPWR 2.60791
R9640 VPWR.n1417 VPWR 2.60791
R9641 VPWR.n1421 VPWR 2.60791
R9642 VPWR.n1426 VPWR 2.60791
R9643 VPWR VPWR.n1428 2.60791
R9644 VPWR.n1723 VPWR 2.60791
R9645 VPWR VPWR.n1722 2.60791
R9646 VPWR.n1716 VPWR 2.60791
R9647 VPWR VPWR.n1714 2.60791
R9648 VPWR.n1461 VPWR 2.60791
R9649 VPWR VPWR.n1707 2.60791
R9650 VPWR VPWR.n1706 2.60791
R9651 VPWR.n1700 VPWR 2.60791
R9652 VPWR VPWR.n1698 2.60791
R9653 VPWR.n1469 VPWR 2.60791
R9654 VPWR.n1692 VPWR 2.60791
R9655 VPWR VPWR.n1691 2.60791
R9656 VPWR VPWR.n1690 2.60791
R9657 VPWR.n1474 VPWR 2.60791
R9658 VPWR.n1684 VPWR 2.60791
R9659 VPWR VPWR.n1682 2.60791
R9660 VPWR.n1477 VPWR 2.60791
R9661 VPWR.n1676 VPWR 2.60791
R9662 VPWR VPWR.n1675 2.60791
R9663 VPWR VPWR.n1674 2.60791
R9664 VPWR.n1482 VPWR 2.60791
R9665 VPWR.n1668 VPWR 2.60791
R9666 VPWR VPWR.n1666 2.60791
R9667 VPWR.n1485 VPWR 2.60791
R9668 VPWR.n1660 VPWR 2.60791
R9669 VPWR VPWR.n1659 2.60791
R9670 VPWR.n1489 VPWR 2.60791
R9671 VPWR.n1652 VPWR 2.60791
R9672 VPWR VPWR.n1651 2.60791
R9673 VPWR VPWR.n1650 2.60791
R9674 VPWR.n1644 VPWR 2.60791
R9675 VPWR VPWR.n1643 2.60791
R9676 VPWR VPWR.n1642 2.60791
R9677 VPWR.n1497 VPWR 2.60791
R9678 VPWR.n1636 VPWR 2.60791
R9679 VPWR VPWR.n1635 2.60791
R9680 VPWR VPWR.n1634 2.60791
R9681 VPWR.n1628 VPWR 2.60791
R9682 VPWR VPWR.n1627 2.60791
R9683 VPWR VPWR.n1626 2.60791
R9684 VPWR.n1505 VPWR 2.60791
R9685 VPWR.n1620 VPWR 2.60791
R9686 VPWR VPWR.n1619 2.60791
R9687 VPWR VPWR.n1618 2.60791
R9688 VPWR VPWR.n1613 2.60791
R9689 VPWR.n953 VPWR 2.60791
R9690 VPWR.n813 VPWR 2.60791
R9691 VPWR.n817 VPWR 2.60791
R9692 VPWR.n821 VPWR 2.60791
R9693 VPWR.n822 VPWR 2.60791
R9694 VPWR.n826 VPWR 2.60791
R9695 VPWR.n830 VPWR 2.60791
R9696 VPWR.n833 VPWR 2.60791
R9697 VPWR.n837 VPWR 2.60791
R9698 VPWR.n841 VPWR 2.60791
R9699 VPWR.n845 VPWR 2.60791
R9700 VPWR.n846 VPWR 2.60791
R9701 VPWR.n849 VPWR 2.60791
R9702 VPWR.n850 VPWR 2.60791
R9703 VPWR.n854 VPWR 2.60791
R9704 VPWR.n857 VPWR 2.60791
R9705 VPWR.n858 VPWR 2.60791
R9706 VPWR.n861 VPWR 2.60791
R9707 VPWR.n865 VPWR 2.60791
R9708 VPWR.n866 VPWR 2.60791
R9709 VPWR.n869 VPWR 2.60791
R9710 VPWR.n870 VPWR 2.60791
R9711 VPWR.n874 VPWR 2.60791
R9712 VPWR.n877 VPWR 2.60791
R9713 VPWR.n878 VPWR 2.60791
R9714 VPWR.n881 VPWR 2.60791
R9715 VPWR.n885 VPWR 2.60791
R9716 VPWR.n886 VPWR 2.60791
R9717 VPWR.n889 VPWR 2.60791
R9718 VPWR.n890 VPWR 2.60791
R9719 VPWR.n894 VPWR 2.60791
R9720 VPWR.n897 VPWR 2.60791
R9721 VPWR.n898 VPWR 2.60791
R9722 VPWR.n902 VPWR 2.60791
R9723 VPWR.n905 VPWR 2.60791
R9724 VPWR.n906 VPWR 2.60791
R9725 VPWR.n910 VPWR 2.60791
R9726 VPWR.n914 VPWR 2.60791
R9727 VPWR.n918 VPWR 2.60791
R9728 VPWR.n923 VPWR 2.60791
R9729 VPWR.n925 VPWR 2.60791
R9730 VPWR.n930 VPWR 2.60791
R9731 VPWR.n1899 VPWR 2.60791
R9732 VPWR VPWR.n1898 2.60791
R9733 VPWR.n1781 VPWR 2.60791
R9734 VPWR.n1785 VPWR 2.60791
R9735 VPWR.n1786 VPWR 2.60791
R9736 VPWR.n1790 VPWR 2.60791
R9737 VPWR.n1794 VPWR 2.60791
R9738 VPWR.n1797 VPWR 2.60791
R9739 VPWR.n1801 VPWR 2.60791
R9740 VPWR.n1805 VPWR 2.60791
R9741 VPWR.n1809 VPWR 2.60791
R9742 VPWR.n1810 VPWR 2.60791
R9743 VPWR.n1813 VPWR 2.60791
R9744 VPWR.n1814 VPWR 2.60791
R9745 VPWR.n1818 VPWR 2.60791
R9746 VPWR.n1821 VPWR 2.60791
R9747 VPWR.n1822 VPWR 2.60791
R9748 VPWR.n1825 VPWR 2.60791
R9749 VPWR.n1829 VPWR 2.60791
R9750 VPWR.n1830 VPWR 2.60791
R9751 VPWR.n1833 VPWR 2.60791
R9752 VPWR.n1834 VPWR 2.60791
R9753 VPWR.n1838 VPWR 2.60791
R9754 VPWR.n1841 VPWR 2.60791
R9755 VPWR.n1842 VPWR 2.60791
R9756 VPWR.n1845 VPWR 2.60791
R9757 VPWR.n1849 VPWR 2.60791
R9758 VPWR.n1850 VPWR 2.60791
R9759 VPWR.n1853 VPWR 2.60791
R9760 VPWR.n1854 VPWR 2.60791
R9761 VPWR.n1858 VPWR 2.60791
R9762 VPWR.n1861 VPWR 2.60791
R9763 VPWR.n1862 VPWR 2.60791
R9764 VPWR.n1866 VPWR 2.60791
R9765 VPWR.n1869 VPWR 2.60791
R9766 VPWR.n1870 VPWR 2.60791
R9767 VPWR.n1874 VPWR 2.60791
R9768 VPWR.n1878 VPWR 2.60791
R9769 VPWR.n1882 VPWR 2.60791
R9770 VPWR.n1886 VPWR 2.60791
R9771 VPWR.n1891 VPWR 2.60791
R9772 VPWR VPWR.n1893 2.60791
R9773 VPWR.n1939 VPWR 2.60791
R9774 VPWR VPWR.n1938 2.60791
R9775 VPWR.n1932 VPWR 2.60791
R9776 VPWR VPWR.n1930 2.60791
R9777 VPWR.n623 VPWR 2.60791
R9778 VPWR.n483 VPWR 2.60791
R9779 VPWR.n487 VPWR 2.60791
R9780 VPWR.n491 VPWR 2.60791
R9781 VPWR.n492 VPWR 2.60791
R9782 VPWR.n496 VPWR 2.60791
R9783 VPWR.n500 VPWR 2.60791
R9784 VPWR.n503 VPWR 2.60791
R9785 VPWR.n507 VPWR 2.60791
R9786 VPWR.n511 VPWR 2.60791
R9787 VPWR.n515 VPWR 2.60791
R9788 VPWR.n516 VPWR 2.60791
R9789 VPWR.n519 VPWR 2.60791
R9790 VPWR.n520 VPWR 2.60791
R9791 VPWR.n524 VPWR 2.60791
R9792 VPWR.n527 VPWR 2.60791
R9793 VPWR.n528 VPWR 2.60791
R9794 VPWR.n531 VPWR 2.60791
R9795 VPWR.n535 VPWR 2.60791
R9796 VPWR.n536 VPWR 2.60791
R9797 VPWR.n539 VPWR 2.60791
R9798 VPWR.n540 VPWR 2.60791
R9799 VPWR.n544 VPWR 2.60791
R9800 VPWR.n547 VPWR 2.60791
R9801 VPWR.n548 VPWR 2.60791
R9802 VPWR.n551 VPWR 2.60791
R9803 VPWR.n555 VPWR 2.60791
R9804 VPWR.n556 VPWR 2.60791
R9805 VPWR.n559 VPWR 2.60791
R9806 VPWR.n560 VPWR 2.60791
R9807 VPWR.n564 VPWR 2.60791
R9808 VPWR.n567 VPWR 2.60791
R9809 VPWR.n568 VPWR 2.60791
R9810 VPWR.n572 VPWR 2.60791
R9811 VPWR.n575 VPWR 2.60791
R9812 VPWR.n576 VPWR 2.60791
R9813 VPWR.n580 VPWR 2.60791
R9814 VPWR.n584 VPWR 2.60791
R9815 VPWR.n588 VPWR 2.60791
R9816 VPWR.n593 VPWR 2.60791
R9817 VPWR.n595 VPWR 2.60791
R9818 VPWR.n600 VPWR 2.60791
R9819 VPWR.n1102 VPWR 2.60791
R9820 VPWR VPWR.n1101 2.60791
R9821 VPWR VPWR.n1087 2.60791
R9822 VPWR.n1131 VPWR 2.60791
R9823 VPWR VPWR.n1083 2.60791
R9824 VPWR.n1139 VPWR 2.60791
R9825 VPWR VPWR.n1140 2.60791
R9826 VPWR.n1148 VPWR 2.60791
R9827 VPWR.n1151 VPWR 2.60791
R9828 VPWR VPWR.n1150 2.60791
R9829 VPWR.n1158 VPWR 2.60791
R9830 VPWR.n1160 VPWR 2.60791
R9831 VPWR.n1165 VPWR 2.60791
R9832 VPWR.n1006 VPWR 2.60791
R9833 VPWR VPWR.n1005 2.60791
R9834 VPWR VPWR.n997 2.60791
R9835 VPWR.n1029 VPWR 2.60791
R9836 VPWR VPWR.n993 2.60791
R9837 VPWR.n1037 VPWR 2.60791
R9838 VPWR VPWR.n1038 2.60791
R9839 VPWR.n1046 VPWR 2.60791
R9840 VPWR.n1049 VPWR 2.60791
R9841 VPWR VPWR.n1048 2.60791
R9842 VPWR.n1056 VPWR 2.60791
R9843 VPWR.n1058 VPWR 2.60791
R9844 VPWR.n1063 VPWR 2.60791
R9845 VPWR VPWR.n2330 2.60791
R9846 VPWR.n2326 VPWR 2.60791
R9847 VPWR VPWR.n2325 2.60791
R9848 VPWR VPWR.n2321 2.60791
R9849 VPWR.n2318 VPWR 2.60791
R9850 VPWR.n2314 VPWR 2.60791
R9851 VPWR.n2310 VPWR 2.60791
R9852 VPWR VPWR.n2309 2.60791
R9853 VPWR VPWR.n2305 2.60791
R9854 VPWR.n2302 VPWR 2.60791
R9855 VPWR.n2298 VPWR 2.60791
R9856 VPWR.n2294 VPWR 2.60791
R9857 VPWR.n2334 VPWR 2.60791
R9858 VPWR.n1734 VPWR.n1733 2.54762
R9859 VPWR.n654 VPWR.n334 2.2505
R9860 VPWR.n972 VPWR.n971 2.2505
R9861 VPWR.n694 VPWR.n693 2.2505
R9862 VPWR.n692 VPWR.n682 2.2505
R9863 VPWR.n197 VPWR.n194 2.2505
R9864 VPWR.n1977 VPWR.n1976 2.2505
R9865 VPWR.n1738 VPWR.n1737 2.2505
R9866 VPWR.n978 VPWR.n329 2.2505
R9867 VPWR.n974 VPWR.n333 2.2505
R9868 VPWR.n977 VPWR.n976 2.2505
R9869 VPWR.n227 VPWR.n226 2.2505
R9870 VPWR.n225 VPWR.n224 2.2505
R9871 VPWR.n685 VPWR.n683 2.2505
R9872 VPWR.n689 VPWR.n688 2.2505
R9873 VPWR.n342 VPWR.n336 2.2505
R9874 VPWR.n651 VPWR.n650 2.2505
R9875 VPWR.n1450 VPWR.n1449 2.2505
R9876 VPWR.n1447 VPWR.n979 2.2505
R9877 VPWR.n73 VPWR.n72 2.2505
R9878 VPWR.n70 VPWR.n67 2.2505
R9879 VPWR.n641 VPWR.n640 2.2505
R9880 VPWR.n639 VPWR.n637 2.2505
R9881 VPWR.n635 VPWR.n634 2.02909
R9882 VPWR.n1275 VPWR.n1249 2.02398
R9883 VPWR.n965 VPWR.n964 2.01887
R9884 VPWR.n1971 VPWR.n1970 1.82542
R9885 VPWR.n969 VPWR.n653 1.68852
R9886 VPWR.n696 VPWR.n695 1.68852
R9887 VPWR.n1974 VPWR.n196 1.68852
R9888 VPWR.n1740 VPWR.n1739 1.68852
R9889 VPWR.n973 VPWR.n254 1.68852
R9890 VPWR.n229 VPWR.n228 1.68852
R9891 VPWR.n686 VPWR.n684 1.68852
R9892 VPWR.n648 VPWR.n341 1.68852
R9893 VPWR.n1446 VPWR.n1175 1.68852
R9894 VPWR.n69 VPWR.n68 1.68852
R9895 VPWR.n643 VPWR.n642 1.68852
R9896 VPWR.n389 VPWR.n388 1.38097
R9897 VPWR.n390 VPWR.n383 1.38097
R9898 VPWR.n391 VPWR.n378 1.38097
R9899 VPWR.n392 VPWR.n373 1.38097
R9900 VPWR.n1273 VPWR.n1254 1.38097
R9901 VPWR.n1272 VPWR.n1259 1.38097
R9902 VPWR.n1271 VPWR.n1264 1.38097
R9903 VPWR.n1270 VPWR.n1269 1.38097
R9904 VPWR.n23 VPWR.n22 1.38097
R9905 VPWR.n24 VPWR.n17 1.38097
R9906 VPWR.n25 VPWR.n12 1.38097
R9907 VPWR.n26 VPWR.n7 1.38097
R9908 VPWR.n679 VPWR.n660 1.38097
R9909 VPWR.n678 VPWR.n665 1.38097
R9910 VPWR.n677 VPWR.n670 1.38097
R9911 VPWR.n676 VPWR.n675 1.38097
R9912 VPWR.n250 VPWR.n249 1.38097
R9913 VPWR.n251 VPWR.n244 1.38097
R9914 VPWR.n252 VPWR.n239 1.38097
R9915 VPWR.n253 VPWR.n234 1.38097
R9916 VPWR.n221 VPWR.n202 1.38097
R9917 VPWR.n220 VPWR.n207 1.38097
R9918 VPWR.n219 VPWR.n212 1.38097
R9919 VPWR.n218 VPWR.n217 1.38097
R9920 VPWR.n719 VPWR.n718 1.38097
R9921 VPWR.n720 VPWR.n713 1.38097
R9922 VPWR.n721 VPWR.n708 1.38097
R9923 VPWR.n722 VPWR.n703 1.38097
R9924 VPWR.n368 VPWR.n349 1.38097
R9925 VPWR.n367 VPWR.n354 1.38097
R9926 VPWR.n366 VPWR.n359 1.38097
R9927 VPWR.n365 VPWR.n364 1.38097
R9928 VPWR.n1911 VPWR.n253 1.28252
R9929 VPWR.n222 VPWR.n221 1.28252
R9930 VPWR.n967 VPWR.n679 1.27742
R9931 VPWR.n966 VPWR.n722 1.27742
R9932 VPWR.n1274 VPWR.n1273 1.27231
R9933 VPWR.n27 VPWR.n26 1.27231
R9934 VPWR.n645 VPWR.n392 1.2672
R9935 VPWR.n646 VPWR.n368 1.2672
R9936 VPWR.n1970 VPWR.n1969 1.10509
R9937 VPWR.n1300 VPWR 1.05698
R9938 VPWR.n763 VPWR 1.05698
R9939 VPWR VPWR.n939 1.05698
R9940 VPWR.n1765 VPWR 1.05698
R9941 VPWR.n309 VPWR 1.05698
R9942 VPWR.n433 VPWR 1.05698
R9943 VPWR VPWR.n609 1.05698
R9944 VPWR.n1230 VPWR 1.05698
R9945 VPWR.n1971 VPWR.n0 0.78681
R9946 VPWR.n1972 VPWR.n1971 0.379389
R9947 VPWR.n697 VPWR.n0 0.379389
R9948 VPWR.n2345 VPWR.n1 0.379389
R9949 VPWR.n2345 VPWR.n2344 0.379389
R9950 VPWR.n1741 VPWR.n1740 0.354022
R9951 VPWR.n1544 VPWR 0.292717
R9952 VPWR.n1602 VPWR 0.292717
R9953 VPWR.n1308 VPWR.n1306 0.270239
R9954 VPWR.n771 VPWR.n769 0.270239
R9955 VPWR.n936 VPWR.n935 0.270239
R9956 VPWR.n1773 VPWR.n1771 0.270239
R9957 VPWR.n317 VPWR.n315 0.270239
R9958 VPWR.n441 VPWR.n439 0.270239
R9959 VPWR.n606 VPWR.n605 0.270239
R9960 VPWR.n1238 VPWR.n1236 0.270239
R9961 VPWR.n1910 VPWR.n1909 0.262576
R9962 VPWR.n965 VPWR.n963 0.257467
R9963 VPWR.n968 VPWR.n655 0.257467
R9964 VPWR.n1276 VPWR.n1275 0.252359
R9965 VPWR.n1445 VPWR.n1444 0.252359
R9966 VPWR.n635 VPWR.n633 0.24725
R9967 VPWR.n647 VPWR.n343 0.24725
R9968 VPWR.n1962 VPWR.t604 0.22969
R9969 VPWR.n1963 VPWR.n1962 0.227365
R9970 VPWR.n1964 VPWR.n1963 0.227365
R9971 VPWR.n1965 VPWR.n1964 0.227365
R9972 VPWR.n1966 VPWR.n1965 0.227365
R9973 VPWR.n1967 VPWR.n1966 0.227365
R9974 VPWR.n1968 VPWR.n1967 0.227365
R9975 VPWR.n1969 VPWR.n1968 0.227365
R9976 VPWR.n1970 VPWR 0.220388
R9977 VPWR VPWR.n391 0.202546
R9978 VPWR VPWR.n390 0.202546
R9979 VPWR VPWR.n389 0.202546
R9980 VPWR VPWR.n1272 0.202546
R9981 VPWR VPWR.n1271 0.202546
R9982 VPWR VPWR.n1270 0.202546
R9983 VPWR VPWR.n25 0.202546
R9984 VPWR VPWR.n24 0.202546
R9985 VPWR VPWR.n23 0.202546
R9986 VPWR VPWR.n678 0.202546
R9987 VPWR VPWR.n677 0.202546
R9988 VPWR VPWR.n676 0.202546
R9989 VPWR VPWR.n252 0.202546
R9990 VPWR VPWR.n251 0.202546
R9991 VPWR VPWR.n250 0.202546
R9992 VPWR VPWR.n220 0.202546
R9993 VPWR VPWR.n219 0.202546
R9994 VPWR VPWR.n218 0.202546
R9995 VPWR VPWR.n721 0.202546
R9996 VPWR VPWR.n720 0.202546
R9997 VPWR VPWR.n719 0.202546
R9998 VPWR VPWR.n367 0.202546
R9999 VPWR VPWR.n366 0.202546
R10000 VPWR VPWR.n365 0.202546
R10001 VPWR.n1302 VPWR 0.157848
R10002 VPWR.n765 VPWR 0.157848
R10003 VPWR VPWR.n938 0.157848
R10004 VPWR.n1767 VPWR 0.157848
R10005 VPWR.n311 VPWR 0.157848
R10006 VPWR.n435 VPWR 0.157848
R10007 VPWR VPWR.n608 0.157848
R10008 VPWR.n1232 VPWR 0.157848
R10009 VPWR.n1911 VPWR.n222 0.155804
R10010 VPWR.n967 VPWR.n966 0.155804
R10011 VPWR.n646 VPWR.n645 0.155804
R10012 VPWR.n1274 VPWR.n27 0.155804
R10013 VPWR.n1911 VPWR.n1910 0.14763
R10014 VPWR.n968 VPWR.n967 0.14763
R10015 VPWR.n966 VPWR.n965 0.14763
R10016 VPWR.n647 VPWR.n646 0.14763
R10017 VPWR.n645 VPWR.n635 0.14763
R10018 VPWR.n1275 VPWR.n1274 0.14763
R10019 VPWR.n1445 VPWR.n27 0.14763
R10020 VPWR.n646 VPWR.n344 0.131283
R10021 VPWR.n645 VPWR.n644 0.131283
R10022 VPWR VPWR.n2346 0.123828
R10023 VPWR.n2343 VPWR.n27 0.120043
R10024 VPWR.n1274 VPWR.n2 0.120043
R10025 VPWR.n1973 VPWR.n222 0.115957
R10026 VPWR.n1912 VPWR.n1911 0.115957
R10027 VPWR.n967 VPWR.n680 0.114935
R10028 VPWR.n966 VPWR.n698 0.114935
R10029 VPWR.n1992 VPWR 0.112891
R10030 VPWR.n179 VPWR 0.112891
R10031 VPWR.n181 VPWR 0.112891
R10032 VPWR.n185 VPWR 0.112891
R10033 VPWR.n187 VPWR 0.112891
R10034 VPWR.n158 VPWR 0.112891
R10035 VPWR.n160 VPWR 0.112891
R10036 VPWR.n164 VPWR 0.112891
R10037 VPWR.n166 VPWR 0.112891
R10038 VPWR.n139 VPWR 0.112891
R10039 VPWR.n141 VPWR 0.112891
R10040 VPWR.n145 VPWR 0.112891
R10041 VPWR.n147 VPWR 0.112891
R10042 VPWR.n118 VPWR 0.112891
R10043 VPWR.n120 VPWR 0.112891
R10044 VPWR.n124 VPWR 0.112891
R10045 VPWR.n126 VPWR 0.112891
R10046 VPWR.n99 VPWR 0.112891
R10047 VPWR.n101 VPWR 0.112891
R10048 VPWR.n105 VPWR 0.112891
R10049 VPWR.n107 VPWR 0.112891
R10050 VPWR.n78 VPWR 0.112891
R10051 VPWR.n80 VPWR 0.112891
R10052 VPWR.n84 VPWR 0.112891
R10053 VPWR.n86 VPWR 0.112891
R10054 VPWR.n1285 VPWR 0.112891
R10055 VPWR.n1298 VPWR 0.112891
R10056 VPWR VPWR.n1298 0.112891
R10057 VPWR.n1516 VPWR 0.112891
R10058 VPWR.n748 VPWR 0.112891
R10059 VPWR.n761 VPWR 0.112891
R10060 VPWR VPWR.n761 0.112891
R10061 VPWR VPWR.n946 0.112891
R10062 VPWR VPWR.n940 0.112891
R10063 VPWR.n940 VPWR 0.112891
R10064 VPWR.n1750 VPWR 0.112891
R10065 VPWR.n1763 VPWR 0.112891
R10066 VPWR VPWR.n1763 0.112891
R10067 VPWR.n294 VPWR 0.112891
R10068 VPWR.n307 VPWR 0.112891
R10069 VPWR VPWR.n307 0.112891
R10070 VPWR.n418 VPWR 0.112891
R10071 VPWR.n431 VPWR 0.112891
R10072 VPWR VPWR.n431 0.112891
R10073 VPWR VPWR.n616 0.112891
R10074 VPWR VPWR.n610 0.112891
R10075 VPWR.n610 VPWR 0.112891
R10076 VPWR.n1123 VPWR 0.112891
R10077 VPWR VPWR.n1122 0.112891
R10078 VPWR.n1023 VPWR 0.112891
R10079 VPWR VPWR.n1022 0.112891
R10080 VPWR.n1215 VPWR 0.112891
R10081 VPWR.n1228 VPWR 0.112891
R10082 VPWR VPWR.n1228 0.112891
R10083 VPWR.n52 VPWR 0.112891
R10084 VPWR.n54 VPWR 0.112891
R10085 VPWR.n58 VPWR 0.112891
R10086 VPWR.n60 VPWR 0.112891
R10087 VPWR.n31 VPWR 0.112891
R10088 VPWR.n33 VPWR 0.112891
R10089 VPWR.n37 VPWR 0.112891
R10090 VPWR.n39 VPWR 0.112891
R10091 VPWR.n1986 VPWR.n1984 0.090413
R10092 VPWR.n1291 VPWR.n1289 0.090413
R10093 VPWR.n1520 VPWR.n1518 0.090413
R10094 VPWR.n1549 VPWR.n1546 0.090413
R10095 VPWR.n1552 VPWR.n1549 0.090413
R10096 VPWR.n1555 VPWR.n1552 0.090413
R10097 VPWR.n1560 VPWR.n1557 0.090413
R10098 VPWR.n1562 VPWR.n1560 0.090413
R10099 VPWR.n1567 VPWR.n1564 0.090413
R10100 VPWR.n1569 VPWR.n1567 0.090413
R10101 VPWR.n1574 VPWR.n1571 0.090413
R10102 VPWR.n1577 VPWR.n1574 0.090413
R10103 VPWR.n1580 VPWR.n1577 0.090413
R10104 VPWR.n754 VPWR.n752 0.090413
R10105 VPWR.n944 VPWR.n943 0.090413
R10106 VPWR.n1756 VPWR.n1754 0.090413
R10107 VPWR.n300 VPWR.n298 0.090413
R10108 VPWR.n424 VPWR.n422 0.090413
R10109 VPWR.n614 VPWR.n613 0.090413
R10110 VPWR.n1221 VPWR.n1219 0.090413
R10111 VPWR.n693 VPWR.n692 0.0711522
R10112 VPWR.n1977 VPWR.n194 0.0711522
R10113 VPWR.n226 VPWR.n225 0.0711522
R10114 VPWR.n689 VPWR.n683 0.0711522
R10115 VPWR.n73 VPWR.n67 0.0711522
R10116 VPWR.n640 VPWR.n639 0.0711522
R10117 VPWR.n1982 VPWR 0.0679348
R10118 VPWR.n1988 VPWR 0.0679348
R10119 VPWR.n1990 VPWR 0.0679348
R10120 VPWR.n1995 VPWR 0.0679348
R10121 VPWR VPWR.n1995 0.0679348
R10122 VPWR.n1997 VPWR 0.0679348
R10123 VPWR.n1999 VPWR 0.0679348
R10124 VPWR.n183 VPWR 0.0679348
R10125 VPWR.n189 VPWR 0.0679348
R10126 VPWR.n191 VPWR 0.0679348
R10127 VPWR.n162 VPWR 0.0679348
R10128 VPWR.n168 VPWR 0.0679348
R10129 VPWR.n170 VPWR 0.0679348
R10130 VPWR.n143 VPWR 0.0679348
R10131 VPWR.n149 VPWR 0.0679348
R10132 VPWR.n151 VPWR 0.0679348
R10133 VPWR.n122 VPWR 0.0679348
R10134 VPWR.n128 VPWR 0.0679348
R10135 VPWR.n130 VPWR 0.0679348
R10136 VPWR.n103 VPWR 0.0679348
R10137 VPWR.n109 VPWR 0.0679348
R10138 VPWR.n111 VPWR 0.0679348
R10139 VPWR.n82 VPWR 0.0679348
R10140 VPWR.n88 VPWR 0.0679348
R10141 VPWR.n90 VPWR 0.0679348
R10142 VPWR.n1283 VPWR 0.0679348
R10143 VPWR.n1287 VPWR 0.0679348
R10144 VPWR.n1293 VPWR 0.0679348
R10145 VPWR.n1295 VPWR 0.0679348
R10146 VPWR.n1304 VPWR 0.0679348
R10147 VPWR VPWR.n1308 0.0679348
R10148 VPWR.n1514 VPWR 0.0679348
R10149 VPWR.n1522 VPWR 0.0679348
R10150 VPWR VPWR.n1544 0.0679348
R10151 VPWR VPWR.n1555 0.0679348
R10152 VPWR VPWR.n1580 0.0679348
R10153 VPWR VPWR.n1602 0.0679348
R10154 VPWR.n746 VPWR 0.0679348
R10155 VPWR.n750 VPWR 0.0679348
R10156 VPWR.n756 VPWR 0.0679348
R10157 VPWR.n758 VPWR 0.0679348
R10158 VPWR.n767 VPWR 0.0679348
R10159 VPWR VPWR.n771 0.0679348
R10160 VPWR VPWR.n947 0.0679348
R10161 VPWR VPWR.n945 0.0679348
R10162 VPWR VPWR.n942 0.0679348
R10163 VPWR VPWR.n941 0.0679348
R10164 VPWR VPWR.n937 0.0679348
R10165 VPWR.n935 VPWR 0.0679348
R10166 VPWR.n1748 VPWR 0.0679348
R10167 VPWR.n1752 VPWR 0.0679348
R10168 VPWR.n1758 VPWR 0.0679348
R10169 VPWR.n1760 VPWR 0.0679348
R10170 VPWR.n1769 VPWR 0.0679348
R10171 VPWR VPWR.n1773 0.0679348
R10172 VPWR.n292 VPWR 0.0679348
R10173 VPWR.n296 VPWR 0.0679348
R10174 VPWR.n302 VPWR 0.0679348
R10175 VPWR.n304 VPWR 0.0679348
R10176 VPWR.n313 VPWR 0.0679348
R10177 VPWR VPWR.n317 0.0679348
R10178 VPWR.n416 VPWR 0.0679348
R10179 VPWR.n420 VPWR 0.0679348
R10180 VPWR.n426 VPWR 0.0679348
R10181 VPWR.n428 VPWR 0.0679348
R10182 VPWR.n437 VPWR 0.0679348
R10183 VPWR VPWR.n441 0.0679348
R10184 VPWR VPWR.n617 0.0679348
R10185 VPWR VPWR.n615 0.0679348
R10186 VPWR VPWR.n612 0.0679348
R10187 VPWR VPWR.n611 0.0679348
R10188 VPWR VPWR.n607 0.0679348
R10189 VPWR.n605 VPWR 0.0679348
R10190 VPWR.n1110 VPWR 0.0679348
R10191 VPWR VPWR.n1124 0.0679348
R10192 VPWR.n1122 VPWR 0.0679348
R10193 VPWR VPWR.n1121 0.0679348
R10194 VPWR.n1012 VPWR 0.0679348
R10195 VPWR VPWR.n1024 0.0679348
R10196 VPWR.n1022 VPWR 0.0679348
R10197 VPWR VPWR.n1021 0.0679348
R10198 VPWR.n1213 VPWR 0.0679348
R10199 VPWR.n1217 VPWR 0.0679348
R10200 VPWR.n1223 VPWR 0.0679348
R10201 VPWR.n1225 VPWR 0.0679348
R10202 VPWR.n1234 VPWR 0.0679348
R10203 VPWR VPWR.n1238 0.0679348
R10204 VPWR.n56 VPWR 0.0679348
R10205 VPWR.n62 VPWR 0.0679348
R10206 VPWR.n64 VPWR 0.0679348
R10207 VPWR.n35 VPWR 0.0679348
R10208 VPWR.n41 VPWR 0.0679348
R10209 VPWR.n43 VPWR 0.0679348
R10210 VPWR VPWR.n1961 0.06442
R10211 VPWR.n1951 VPWR 0.06066
R10212 VPWR.n1956 VPWR 0.06066
R10213 VPWR.n648 VPWR.n647 0.0602717
R10214 VPWR.n1446 VPWR.n1445 0.055163
R10215 VPWR.n1973 VPWR.n1972 0.0522
R10216 VPWR.n969 VPWR.n968 0.0500543
R10217 VPWR.n344 VPWR.n1 0.0490667
R10218 VPWR.n644 VPWR.n1 0.0471867
R10219 VPWR.n2077 VPWR.n2000 0.0454565
R10220 VPWR.n2079 VPWR.n193 0.0454565
R10221 VPWR.n2142 VPWR.n171 0.0454565
R10222 VPWR.n2145 VPWR.n153 0.0454565
R10223 VPWR.n2208 VPWR.n131 0.0454565
R10224 VPWR.n2211 VPWR.n113 0.0454565
R10225 VPWR.n2274 VPWR.n91 0.0454565
R10226 VPWR.n1281 VPWR.n1276 0.0454565
R10227 VPWR.n1311 VPWR.n1310 0.0454565
R10228 VPWR.n1733 VPWR.n1452 0.0454565
R10229 VPWR.n1607 VPWR.n1606 0.0454565
R10230 VPWR.n963 VPWR.n723 0.0454565
R10231 VPWR.n776 VPWR.n775 0.0454565
R10232 VPWR.n948 VPWR.n655 0.0454565
R10233 VPWR.n934 VPWR.n740 0.0454565
R10234 VPWR.n1746 VPWR.n1741 0.0454565
R10235 VPWR.n1776 VPWR.n1775 0.0454565
R10236 VPWR.n1909 VPWR.n255 0.0454565
R10237 VPWR.n322 VPWR.n321 0.0454565
R10238 VPWR.n633 VPWR.n393 0.0454565
R10239 VPWR.n446 VPWR.n445 0.0454565
R10240 VPWR.n618 VPWR.n343 0.0454565
R10241 VPWR.n604 VPWR.n410 0.0454565
R10242 VPWR.n1125 VPWR.n1114 0.0454565
R10243 VPWR.n1171 VPWR.n1069 0.0454565
R10244 VPWR.n1025 VPWR.n1014 0.0454565
R10245 VPWR.n1067 VPWR.n983 0.0454565
R10246 VPWR.n1444 VPWR.n1176 0.0454565
R10247 VPWR.n1243 VPWR.n1242 0.0454565
R10248 VPWR.n2277 VPWR.n66 0.0454565
R10249 VPWR.n2340 VPWR.n44 0.0454565
R10250 VPWR.n1910 VPWR.n254 0.0449457
R10251 VPWR.n1972 VPWR.n1912 0.0440533
R10252 VPWR.n1961 VPWR.n1956 0.04186
R10253 VPWR.n697 VPWR.n680 0.0409722
R10254 VPWR.n698 VPWR.n697 0.0394056
R10255 VPWR.n2344 VPWR.n2 0.0388421
R10256 VPWR.n2344 VPWR.n2343 0.0373579
R10257 VPWR.n1974 VPWR.n1973 0.0367717
R10258 VPWR.n1912 VPWR.n229 0.0367717
R10259 VPWR.n644 VPWR.n643 0.0367717
R10260 VPWR.n981 VPWR.n972 0.0361924
R10261 VPWR.n978 VPWR.n330 0.0361924
R10262 VPWR.n980 VPWR.n977 0.0361924
R10263 VPWR.n982 VPWR.n651 0.0361924
R10264 VPWR.n982 VPWR.n336 0.0361924
R10265 VPWR.n981 VPWR.n334 0.0361924
R10266 VPWR.n980 VPWR.n333 0.0361924
R10267 VPWR.n1737 VPWR.n330 0.0361924
R10268 VPWR.n1450 VPWR.n331 0.0361924
R10269 VPWR.n979 VPWR.n331 0.0361924
R10270 VPWR.n971 VPWR.n653 0.0359639
R10271 VPWR.n654 VPWR.n653 0.0359639
R10272 VPWR.n695 VPWR.n682 0.0359639
R10273 VPWR.n695 VPWR.n694 0.0359639
R10274 VPWR.n1976 VPWR.n196 0.0359639
R10275 VPWR.n197 VPWR.n196 0.0359639
R10276 VPWR.n1739 VPWR.n329 0.0359639
R10277 VPWR.n1739 VPWR.n1738 0.0359639
R10278 VPWR.n976 VPWR.n973 0.0359639
R10279 VPWR.n974 VPWR.n973 0.0359639
R10280 VPWR.n228 VPWR.n224 0.0359639
R10281 VPWR.n228 VPWR.n227 0.0359639
R10282 VPWR.n688 VPWR.n684 0.0359639
R10283 VPWR.n685 VPWR.n684 0.0359639
R10284 VPWR.n650 VPWR.n341 0.0359639
R10285 VPWR.n342 VPWR.n341 0.0359639
R10286 VPWR.n1447 VPWR.n1175 0.0359639
R10287 VPWR.n1449 VPWR.n1175 0.0359639
R10288 VPWR.n70 VPWR.n68 0.0359639
R10289 VPWR.n72 VPWR.n68 0.0359639
R10290 VPWR.n642 VPWR.n637 0.0359639
R10291 VPWR.n642 VPWR.n641 0.0359639
R10292 VPWR.n1735 VPWR.n1734 0.0357905
R10293 VPWR.n964 VPWR.n652 0.0357905
R10294 VPWR.n634 VPWR.n340 0.0357905
R10295 VPWR.n1734 VPWR.n332 0.0357863
R10296 VPWR.n964 VPWR.n335 0.0357863
R10297 VPWR.n634 VPWR.n337 0.0357863
R10298 VPWR.n1249 VPWR.n338 0.0357863
R10299 VPWR.n698 VPWR.n696 0.0275761
R10300 VPWR.n686 VPWR.n680 0.0275761
R10301 VPWR.n970 VPWR.n969 0.0270652
R10302 VPWR.n696 VPWR.n681 0.0270652
R10303 VPWR.n1975 VPWR.n1974 0.0270652
R10304 VPWR.n1740 VPWR.n328 0.0270652
R10305 VPWR.n975 VPWR.n254 0.0270652
R10306 VPWR.n229 VPWR.n223 0.0270652
R10307 VPWR.n687 VPWR.n686 0.0270652
R10308 VPWR.n649 VPWR.n648 0.0270652
R10309 VPWR.n1448 VPWR.n1446 0.0270652
R10310 VPWR.n71 VPWR.n69 0.0270652
R10311 VPWR.n643 VPWR.n636 0.0270652
R10312 VPWR.n1451 VPWR.n339 0.026751
R10313 VPWR.n1736 VPWR.n339 0.026751
R10314 VPWR.n392 VPWR 0.0250279
R10315 VPWR.n391 VPWR 0.0250279
R10316 VPWR.n390 VPWR 0.0250279
R10317 VPWR.n389 VPWR 0.0250279
R10318 VPWR.n1273 VPWR 0.0250279
R10319 VPWR.n1272 VPWR 0.0250279
R10320 VPWR.n1271 VPWR 0.0250279
R10321 VPWR.n1270 VPWR 0.0250279
R10322 VPWR.n26 VPWR 0.0250279
R10323 VPWR.n25 VPWR 0.0250279
R10324 VPWR.n24 VPWR 0.0250279
R10325 VPWR.n23 VPWR 0.0250279
R10326 VPWR.n679 VPWR 0.0250279
R10327 VPWR.n678 VPWR 0.0250279
R10328 VPWR.n677 VPWR 0.0250279
R10329 VPWR.n676 VPWR 0.0250279
R10330 VPWR.n253 VPWR 0.0250279
R10331 VPWR.n252 VPWR 0.0250279
R10332 VPWR.n251 VPWR 0.0250279
R10333 VPWR.n250 VPWR 0.0250279
R10334 VPWR.n221 VPWR 0.0250279
R10335 VPWR.n220 VPWR 0.0250279
R10336 VPWR.n219 VPWR 0.0250279
R10337 VPWR.n218 VPWR 0.0250279
R10338 VPWR.n722 VPWR 0.0250279
R10339 VPWR.n721 VPWR 0.0250279
R10340 VPWR.n720 VPWR 0.0250279
R10341 VPWR.n719 VPWR 0.0250279
R10342 VPWR.n368 VPWR 0.0250279
R10343 VPWR.n367 VPWR 0.0250279
R10344 VPWR.n366 VPWR 0.0250279
R10345 VPWR.n365 VPWR 0.0250279
R10346 VPWR.n2345 VPWR.n0 0.024
R10347 VPWR VPWR.n1946 0.02306
R10348 VPWR VPWR.n1951 0.02306
R10349 VPWR VPWR.n1982 0.0229783
R10350 VPWR.n1984 VPWR 0.0229783
R10351 VPWR VPWR.n1986 0.0229783
R10352 VPWR VPWR.n1988 0.0229783
R10353 VPWR VPWR.n1990 0.0229783
R10354 VPWR VPWR.n1992 0.0229783
R10355 VPWR VPWR.n1997 0.0229783
R10356 VPWR VPWR.n1999 0.0229783
R10357 VPWR.n2000 VPWR 0.0229783
R10358 VPWR VPWR.n2077 0.0229783
R10359 VPWR VPWR.n179 0.0229783
R10360 VPWR VPWR.n181 0.0229783
R10361 VPWR VPWR.n183 0.0229783
R10362 VPWR VPWR.n185 0.0229783
R10363 VPWR VPWR.n187 0.0229783
R10364 VPWR VPWR.n189 0.0229783
R10365 VPWR VPWR.n191 0.0229783
R10366 VPWR.n193 VPWR 0.0229783
R10367 VPWR.n2079 VPWR 0.0229783
R10368 VPWR VPWR.n158 0.0229783
R10369 VPWR VPWR.n160 0.0229783
R10370 VPWR VPWR.n162 0.0229783
R10371 VPWR VPWR.n164 0.0229783
R10372 VPWR VPWR.n166 0.0229783
R10373 VPWR VPWR.n168 0.0229783
R10374 VPWR VPWR.n170 0.0229783
R10375 VPWR.n171 VPWR 0.0229783
R10376 VPWR VPWR.n2142 0.0229783
R10377 VPWR VPWR.n139 0.0229783
R10378 VPWR VPWR.n141 0.0229783
R10379 VPWR VPWR.n143 0.0229783
R10380 VPWR VPWR.n145 0.0229783
R10381 VPWR VPWR.n147 0.0229783
R10382 VPWR VPWR.n149 0.0229783
R10383 VPWR VPWR.n151 0.0229783
R10384 VPWR.n153 VPWR 0.0229783
R10385 VPWR.n2145 VPWR 0.0229783
R10386 VPWR VPWR.n118 0.0229783
R10387 VPWR VPWR.n120 0.0229783
R10388 VPWR VPWR.n122 0.0229783
R10389 VPWR VPWR.n124 0.0229783
R10390 VPWR VPWR.n126 0.0229783
R10391 VPWR VPWR.n128 0.0229783
R10392 VPWR VPWR.n130 0.0229783
R10393 VPWR.n131 VPWR 0.0229783
R10394 VPWR VPWR.n2208 0.0229783
R10395 VPWR VPWR.n99 0.0229783
R10396 VPWR VPWR.n101 0.0229783
R10397 VPWR VPWR.n103 0.0229783
R10398 VPWR VPWR.n105 0.0229783
R10399 VPWR VPWR.n107 0.0229783
R10400 VPWR VPWR.n109 0.0229783
R10401 VPWR VPWR.n111 0.0229783
R10402 VPWR.n113 VPWR 0.0229783
R10403 VPWR.n2211 VPWR 0.0229783
R10404 VPWR VPWR.n78 0.0229783
R10405 VPWR VPWR.n80 0.0229783
R10406 VPWR VPWR.n82 0.0229783
R10407 VPWR VPWR.n84 0.0229783
R10408 VPWR VPWR.n86 0.0229783
R10409 VPWR VPWR.n88 0.0229783
R10410 VPWR VPWR.n90 0.0229783
R10411 VPWR.n91 VPWR 0.0229783
R10412 VPWR VPWR.n2274 0.0229783
R10413 VPWR VPWR.n1281 0.0229783
R10414 VPWR VPWR.n1283 0.0229783
R10415 VPWR VPWR.n1285 0.0229783
R10416 VPWR VPWR.n1287 0.0229783
R10417 VPWR.n1289 VPWR 0.0229783
R10418 VPWR VPWR.n1291 0.0229783
R10419 VPWR VPWR.n1293 0.0229783
R10420 VPWR VPWR.n1295 0.0229783
R10421 VPWR VPWR.n1300 0.0229783
R10422 VPWR VPWR.n1302 0.0229783
R10423 VPWR VPWR.n1304 0.0229783
R10424 VPWR.n1306 VPWR 0.0229783
R10425 VPWR.n1310 VPWR 0.0229783
R10426 VPWR.n1311 VPWR 0.0229783
R10427 VPWR VPWR.n1452 0.0229783
R10428 VPWR VPWR.n1514 0.0229783
R10429 VPWR VPWR.n1516 0.0229783
R10430 VPWR.n1518 VPWR 0.0229783
R10431 VPWR VPWR.n1520 0.0229783
R10432 VPWR VPWR.n1522 0.0229783
R10433 VPWR.n1546 VPWR 0.0229783
R10434 VPWR.n1557 VPWR 0.0229783
R10435 VPWR VPWR.n1562 0.0229783
R10436 VPWR.n1564 VPWR 0.0229783
R10437 VPWR VPWR.n1569 0.0229783
R10438 VPWR.n1571 VPWR 0.0229783
R10439 VPWR.n1606 VPWR 0.0229783
R10440 VPWR.n1607 VPWR 0.0229783
R10441 VPWR VPWR.n723 0.0229783
R10442 VPWR VPWR.n746 0.0229783
R10443 VPWR VPWR.n748 0.0229783
R10444 VPWR VPWR.n750 0.0229783
R10445 VPWR.n752 VPWR 0.0229783
R10446 VPWR VPWR.n754 0.0229783
R10447 VPWR VPWR.n756 0.0229783
R10448 VPWR VPWR.n758 0.0229783
R10449 VPWR VPWR.n763 0.0229783
R10450 VPWR VPWR.n765 0.0229783
R10451 VPWR VPWR.n767 0.0229783
R10452 VPWR.n769 VPWR 0.0229783
R10453 VPWR.n775 VPWR 0.0229783
R10454 VPWR.n776 VPWR 0.0229783
R10455 VPWR.n948 VPWR 0.0229783
R10456 VPWR.n947 VPWR 0.0229783
R10457 VPWR.n946 VPWR 0.0229783
R10458 VPWR.n945 VPWR 0.0229783
R10459 VPWR VPWR.n944 0.0229783
R10460 VPWR.n943 VPWR 0.0229783
R10461 VPWR.n942 VPWR 0.0229783
R10462 VPWR.n941 VPWR 0.0229783
R10463 VPWR.n939 VPWR 0.0229783
R10464 VPWR.n938 VPWR 0.0229783
R10465 VPWR.n937 VPWR 0.0229783
R10466 VPWR VPWR.n936 0.0229783
R10467 VPWR VPWR.n934 0.0229783
R10468 VPWR.n740 VPWR 0.0229783
R10469 VPWR VPWR.n1746 0.0229783
R10470 VPWR VPWR.n1748 0.0229783
R10471 VPWR VPWR.n1750 0.0229783
R10472 VPWR VPWR.n1752 0.0229783
R10473 VPWR.n1754 VPWR 0.0229783
R10474 VPWR VPWR.n1756 0.0229783
R10475 VPWR VPWR.n1758 0.0229783
R10476 VPWR VPWR.n1760 0.0229783
R10477 VPWR VPWR.n1765 0.0229783
R10478 VPWR VPWR.n1767 0.0229783
R10479 VPWR VPWR.n1769 0.0229783
R10480 VPWR.n1771 VPWR 0.0229783
R10481 VPWR.n1775 VPWR 0.0229783
R10482 VPWR.n1776 VPWR 0.0229783
R10483 VPWR VPWR.n255 0.0229783
R10484 VPWR VPWR.n292 0.0229783
R10485 VPWR VPWR.n294 0.0229783
R10486 VPWR VPWR.n296 0.0229783
R10487 VPWR.n298 VPWR 0.0229783
R10488 VPWR VPWR.n300 0.0229783
R10489 VPWR VPWR.n302 0.0229783
R10490 VPWR VPWR.n304 0.0229783
R10491 VPWR VPWR.n309 0.0229783
R10492 VPWR VPWR.n311 0.0229783
R10493 VPWR VPWR.n313 0.0229783
R10494 VPWR.n315 VPWR 0.0229783
R10495 VPWR.n321 VPWR 0.0229783
R10496 VPWR.n322 VPWR 0.0229783
R10497 VPWR VPWR.n393 0.0229783
R10498 VPWR VPWR.n416 0.0229783
R10499 VPWR VPWR.n418 0.0229783
R10500 VPWR VPWR.n420 0.0229783
R10501 VPWR.n422 VPWR 0.0229783
R10502 VPWR VPWR.n424 0.0229783
R10503 VPWR VPWR.n426 0.0229783
R10504 VPWR VPWR.n428 0.0229783
R10505 VPWR VPWR.n433 0.0229783
R10506 VPWR VPWR.n435 0.0229783
R10507 VPWR VPWR.n437 0.0229783
R10508 VPWR.n439 VPWR 0.0229783
R10509 VPWR.n445 VPWR 0.0229783
R10510 VPWR.n446 VPWR 0.0229783
R10511 VPWR.n618 VPWR 0.0229783
R10512 VPWR.n617 VPWR 0.0229783
R10513 VPWR.n616 VPWR 0.0229783
R10514 VPWR.n615 VPWR 0.0229783
R10515 VPWR VPWR.n614 0.0229783
R10516 VPWR.n613 VPWR 0.0229783
R10517 VPWR.n612 VPWR 0.0229783
R10518 VPWR.n611 VPWR 0.0229783
R10519 VPWR.n609 VPWR 0.0229783
R10520 VPWR.n608 VPWR 0.0229783
R10521 VPWR.n607 VPWR 0.0229783
R10522 VPWR VPWR.n606 0.0229783
R10523 VPWR VPWR.n604 0.0229783
R10524 VPWR.n410 VPWR 0.0229783
R10525 VPWR VPWR.n1108 0.0229783
R10526 VPWR VPWR.n1110 0.0229783
R10527 VPWR.n1114 VPWR 0.0229783
R10528 VPWR.n1125 VPWR 0.0229783
R10529 VPWR.n1124 VPWR 0.0229783
R10530 VPWR VPWR.n1123 0.0229783
R10531 VPWR.n1121 VPWR 0.0229783
R10532 VPWR VPWR.n1069 0.0229783
R10533 VPWR VPWR.n1171 0.0229783
R10534 VPWR VPWR.n1010 0.0229783
R10535 VPWR VPWR.n1012 0.0229783
R10536 VPWR.n1014 VPWR 0.0229783
R10537 VPWR.n1025 VPWR 0.0229783
R10538 VPWR.n1024 VPWR 0.0229783
R10539 VPWR VPWR.n1023 0.0229783
R10540 VPWR.n1021 VPWR 0.0229783
R10541 VPWR VPWR.n983 0.0229783
R10542 VPWR VPWR.n1067 0.0229783
R10543 VPWR VPWR.n1176 0.0229783
R10544 VPWR VPWR.n1213 0.0229783
R10545 VPWR VPWR.n1215 0.0229783
R10546 VPWR VPWR.n1217 0.0229783
R10547 VPWR.n1219 VPWR 0.0229783
R10548 VPWR VPWR.n1221 0.0229783
R10549 VPWR VPWR.n1223 0.0229783
R10550 VPWR VPWR.n1225 0.0229783
R10551 VPWR VPWR.n1230 0.0229783
R10552 VPWR VPWR.n1232 0.0229783
R10553 VPWR VPWR.n1234 0.0229783
R10554 VPWR.n1236 VPWR 0.0229783
R10555 VPWR.n1242 VPWR 0.0229783
R10556 VPWR.n1243 VPWR 0.0229783
R10557 VPWR VPWR.n52 0.0229783
R10558 VPWR VPWR.n54 0.0229783
R10559 VPWR VPWR.n56 0.0229783
R10560 VPWR VPWR.n58 0.0229783
R10561 VPWR VPWR.n60 0.0229783
R10562 VPWR VPWR.n62 0.0229783
R10563 VPWR VPWR.n64 0.0229783
R10564 VPWR.n66 VPWR 0.0229783
R10565 VPWR.n2277 VPWR 0.0229783
R10566 VPWR VPWR.n31 0.0229783
R10567 VPWR VPWR.n33 0.0229783
R10568 VPWR VPWR.n35 0.0229783
R10569 VPWR VPWR.n37 0.0229783
R10570 VPWR VPWR.n39 0.0229783
R10571 VPWR VPWR.n41 0.0229783
R10572 VPWR VPWR.n43 0.0229783
R10573 VPWR.n44 VPWR 0.0229783
R10574 VPWR VPWR.n2340 0.0229783
R10575 VPWR.n69 VPWR.n2 0.0224674
R10576 VPWR.n1451 VPWR.n1174 0.0203634
R10577 VPWR.n1962 VPWR.t602 0.00282438
R10578 VPWR.n1963 VPWR.t607 0.00282438
R10579 VPWR.n1964 VPWR.t608 0.00282438
R10580 VPWR.n1965 VPWR.t606 0.00282438
R10581 VPWR.n1966 VPWR.t603 0.00282438
R10582 VPWR.n1967 VPWR.t605 0.00282438
R10583 VPWR.n1968 VPWR.t610 0.00282438
R10584 VPWR.n1969 VPWR.t609 0.00282438
R10585 VPWR.n2346 VPWR.n2345 0.000985236
R10586 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t4 1060.4
R10587 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t9 1060.4
R10588 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t2 1060.4
R10589 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t3 1060.4
R10590 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n3 568.956
R10591 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t8 568.956
R10592 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n5 568.956
R10593 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t6 568.956
R10594 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t5 568.956
R10595 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n8 568.956
R10596 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t7 568.956
R10597 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n2 568.956
R10598 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.D SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t1 376.673
R10599 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.t0 131.389
R10600 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.D 121.977
R10601 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n3 20.3299
R10602 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA4.XA4.MP3.G 20.3299
R10603 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA4.XA4.MN3.G 20.3299
R10604 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n2 20.3299
R10605 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n4 20.3299
R10606 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA4.XA4.MN2.G 20.3299
R10607 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA4.XA4.MP2.G 20.3299
R10608 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA4.XA4.MP0.G 20.3299
R10609 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n7 20.3299
R10610 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n6 20.3299
R10611 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA4.XA4.MP1.G 20.3299
R10612 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA4.XA4.MN1.G 20.3299
R10613 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n2 20.3299
R10614 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n0 12.8005
R10615 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA4.XA4.MN0.G 10.6968
R10616 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n1 9.49168
R10617 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n10 9.47055
R10618 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n11 9.3005
R10619 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n12 7.52991
R10620 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n0 6.77697
R10621 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n9 5.36434
R10622 SUNSAR_SAR8B_CV_0.XA4.CP0.t15 SUNSAR_SAR8B_CV_0.XA4.CP0.t10 1060.4
R10623 SUNSAR_SAR8B_CV_0.XA4.CP0.t8 SUNSAR_SAR8B_CV_0.XA4.CP0.t9 1060.4
R10624 SUNSAR_SAR8B_CV_0.XA4.CP0.t13 SUNSAR_SAR8B_CV_0.XA4.CP0.t12 1060.4
R10625 SUNSAR_SAR8B_CV_0.XA4.CP0.t11 SUNSAR_SAR8B_CV_0.XA4.CP0.t14 1060.4
R10626 SUNSAR_SAR8B_CV_0.XA4.CP0.t10 SUNSAR_SAR8B_CV_0.XA4.CP0.n4 568.956
R10627 SUNSAR_SAR8B_CV_0.XA4.CP0.n5 SUNSAR_SAR8B_CV_0.XA4.CP0.t15 568.956
R10628 SUNSAR_SAR8B_CV_0.XA4.CP0.t9 SUNSAR_SAR8B_CV_0.XA4.CP0.n6 568.956
R10629 SUNSAR_SAR8B_CV_0.XA4.CP0.n7 SUNSAR_SAR8B_CV_0.XA4.CP0.t8 568.956
R10630 SUNSAR_SAR8B_CV_0.XA4.CP0.n10 SUNSAR_SAR8B_CV_0.XA4.CP0.t13 568.956
R10631 SUNSAR_SAR8B_CV_0.XA4.CP0.t12 SUNSAR_SAR8B_CV_0.XA4.CP0.n9 568.956
R10632 SUNSAR_SAR8B_CV_0.XA4.CP0.n8 SUNSAR_SAR8B_CV_0.XA4.CP0.t11 568.956
R10633 SUNSAR_SAR8B_CV_0.XA4.CP0.t14 SUNSAR_SAR8B_CV_0.XA4.CP0.n3 568.956
R10634 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.CP0.n1 312.829
R10635 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.CP0.n0 312.829
R10636 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.CP0.n10 197.272
R10637 SUNSAR_SAR8B_CV_0.XA4.CP0.n12 SUNSAR_SAR8B_CV_0.XA4.CP0.n11 92.5005
R10638 SUNSAR_SAR8B_CV_0.XA4.CP0.n15 SUNSAR_SAR8B_CV_0.XA4.CP0.n14 92.5005
R10639 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.CP0.n16 90.7299
R10640 SUNSAR_SAR8B_CV_0.XA4.CP0.n0 SUNSAR_SAR8B_CV_0.XA4.CP0.t5 63.8431
R10641 SUNSAR_SAR8B_CV_0.XA4.CP0.n0 SUNSAR_SAR8B_CV_0.XA4.CP0.t6 63.8431
R10642 SUNSAR_SAR8B_CV_0.XA4.CP0.n1 SUNSAR_SAR8B_CV_0.XA4.CP0.t4 63.8431
R10643 SUNSAR_SAR8B_CV_0.XA4.CP0.n1 SUNSAR_SAR8B_CV_0.XA4.CP0.t7 63.8431
R10644 SUNSAR_SAR8B_CV_0.XA4.CP0.n2 SUNSAR_SAR8B_CV_0.XA4.CP0 61.177
R10645 SUNSAR_SAR8B_CV_0.XA4.CP0.n16 SUNSAR_SAR8B_CV_0.XA4.CP0.n13 53.4593
R10646 SUNSAR_SAR8B_CV_0.XA4.CP0.n11 SUNSAR_SAR8B_CV_0.XA4.CP0.t1 38.8894
R10647 SUNSAR_SAR8B_CV_0.XA4.CP0.n11 SUNSAR_SAR8B_CV_0.XA4.CP0.t0 38.8894
R10648 SUNSAR_SAR8B_CV_0.XA4.CP0.n14 SUNSAR_SAR8B_CV_0.XA4.CP0.t3 38.8894
R10649 SUNSAR_SAR8B_CV_0.XA4.CP0.n14 SUNSAR_SAR8B_CV_0.XA4.CP0.t2 38.8894
R10650 SUNSAR_SAR8B_CV_0.XA4.CP0.n13 SUNSAR_SAR8B_CV_0.XA4.CP0.n12 38.024
R10651 SUNSAR_SAR8B_CV_0.XA4.CP0.n16 SUNSAR_SAR8B_CV_0.XA4.CP0.n15 38.024
R10652 SUNSAR_SAR8B_CV_0.XA4.CP0.n13 SUNSAR_SAR8B_CV_0.XA4.CP0.n2 29.5534
R10653 SUNSAR_SAR8B_CV_0.XA4.CP0.n7 SUNSAR_SAR8B_CV_0.XA4.CP0.n4 20.3299
R10654 SUNSAR_SAR8B_CV_0.XA4.CP0.n4 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10655 SUNSAR_SAR8B_CV_0.XA4.CP0.n5 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10656 SUNSAR_SAR8B_CV_0.XA4.CP0.n6 SUNSAR_SAR8B_CV_0.XA4.CP0.n3 20.3299
R10657 SUNSAR_SAR8B_CV_0.XA4.CP0.n6 SUNSAR_SAR8B_CV_0.XA4.CP0.n5 20.3299
R10658 SUNSAR_SAR8B_CV_0.XA4.CP0.n6 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10659 SUNSAR_SAR8B_CV_0.XA4.CP0.n7 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10660 SUNSAR_SAR8B_CV_0.XA4.CP0.n9 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10661 SUNSAR_SAR8B_CV_0.XA4.CP0.n9 SUNSAR_SAR8B_CV_0.XA4.CP0.n8 20.3299
R10662 SUNSAR_SAR8B_CV_0.XA4.CP0.n8 SUNSAR_SAR8B_CV_0.XA4.CP0.n7 20.3299
R10663 SUNSAR_SAR8B_CV_0.XA4.CP0.n8 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10664 SUNSAR_SAR8B_CV_0.XA4.CP0.n3 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10665 SUNSAR_SAR8B_CV_0.XA4.CP0.n10 SUNSAR_SAR8B_CV_0.XA4.CP0.n3 20.3299
R10666 SUNSAR_SAR8B_CV_0.XA4.CP0.n10 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10667 SUNSAR_SAR8B_CV_0.XA4.CP0.n12 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10668 SUNSAR_SAR8B_CV_0.XA4.CP0.n15 SUNSAR_SAR8B_CV_0.XA4.CP0 20.3299
R10669 SUNSAR_SAR8B_CV_0.XA4.CP0.n2 SUNSAR_SAR8B_CV_0.XA4.CP0 10.3476
R10670 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t10 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t4 1060.4
R10671 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t11 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t2 1060.4
R10672 SUNSAR_SAR8B_CV_0.XA20.XA1.MN6.G SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t3 589.284
R10673 SUNSAR_SAR8B_CV_0.XA20.XA2.MN0.G SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t10 589.284
R10674 SUNSAR_SAR8B_CV_0.XA20.XA3.MN0.G SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t11 589.284
R10675 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n9 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n4 583.529
R10676 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n10 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t9 568.956
R10677 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n0 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t6 568.956
R10678 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n1 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t8 568.956
R10679 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t4 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n3 568.956
R10680 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n5 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t7 568.956
R10681 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n6 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t5 568.956
R10682 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n8 568.956
R10683 SUNSAR_SAR8B_CV_0.XA20.XA4.MN6.G SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n9 468.707
R10684 SUNSAR_SAR8B_CV_0.XA20.XA9.MP0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t1 376.673
R10685 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n11 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.t0 131.389
R10686 SUNSAR_SAR8B_CV_0.XA20.XA9.MN0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n10 131.012
R10687 SUNSAR_SAR8B_CV_0.XA20.XA9.MP0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n11 128.754
R10688 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n0 91.4829
R10689 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n7 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n5 91.4829
R10690 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n4 SUNSAR_SAR8B_CV_0.XA20.XA1.MN6.G 71.1534
R10691 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n3 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n2 58.3534
R10692 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n8 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n7 58.3534
R10693 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n2 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n1 38.024
R10694 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n7 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n6 38.024
R10695 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n0 SUNSAR_SAR8B_CV_0.XA20.XA2.MP3.G 20.3299
R10696 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n1 SUNSAR_SAR8B_CV_0.XA20.XA2.MP1.G 20.3299
R10697 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.MP0.G 20.3299
R10698 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n5 SUNSAR_SAR8B_CV_0.XA20.XA3.MP3.G 20.3299
R10699 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n6 SUNSAR_SAR8B_CV_0.XA20.XA3.MP1.G 20.3299
R10700 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n8 SUNSAR_SAR8B_CV_0.XA20.XA3.MP0.G 20.3299
R10701 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n10 SUNSAR_SAR8B_CV_0.XA20.XA4.MN6.G 20.3299
R10702 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n11 SUNSAR_SAR8B_CV_0.XA20.XA9.MN0.D 20.3299
R10703 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n4 SUNSAR_SAR8B_CV_0.XA20.XA2.MN0.G 17.6946
R10704 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n9 SUNSAR_SAR8B_CV_0.XA20.XA3.MN0.G 17.6946
R10705 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t8 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t29 1060.4
R10706 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t30 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t31 1060.4
R10707 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t11 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t10 1060.4
R10708 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t16 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t27 1060.4
R10709 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t15 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t22 1060.4
R10710 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t23 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t9 1060.4
R10711 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t24 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t20 1060.4
R10712 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t13 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t26 1060.4
R10713 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t29 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10714 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t31 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10715 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t10 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10716 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t27 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10717 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t22 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10718 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t9 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10719 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t20 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10720 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t26 SUNSAR_SAR8B_CV_0.XA20.CPO 589.284
R10721 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n53 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t8 574.383
R10722 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n34 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t11 574.383
R10723 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n24 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t15 574.383
R10724 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n14 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t24 574.383
R10725 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n39 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t30 572.859
R10726 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n29 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t16 572.859
R10727 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n19 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t23 572.859
R10728 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n9 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t13 572.859
R10729 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n51 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t17 568.956
R10730 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n41 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t28 568.956
R10731 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n37 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t19 568.956
R10732 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n31 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t21 568.956
R10733 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n27 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t25 568.956
R10734 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n21 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t12 568.956
R10735 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n17 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t14 568.956
R10736 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n11 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t18 568.956
R10737 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n2 312.829
R10738 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n6 312.829
R10739 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n4 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n3 92.5005
R10740 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n1 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n0 92.5005
R10741 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n5 SUNSAR_SAR8B_CV_0.XA20.CPO 90.7299
R10742 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n7 SUNSAR_SAR8B_CV_0.XA20.CPO 90.7299
R10743 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n6 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t1 63.8431
R10744 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n6 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t7 63.8431
R10745 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n2 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t4 63.8431
R10746 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n2 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t3 63.8431
R10747 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n7 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n5 53.4593
R10748 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n3 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t6 38.8894
R10749 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n3 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t2 38.8894
R10750 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n0 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t0 38.8894
R10751 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n0 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.t5 38.8894
R10752 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n5 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n4 38.024
R10753 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n8 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n7 22.7142
R10754 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n41 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n40 22.1005
R10755 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n31 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n30 22.1005
R10756 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n21 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n20 22.1005
R10757 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n11 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n10 22.1005
R10758 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n4 SUNSAR_SAR8B_CV_0.XA20.CPO 20.3299
R10759 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n38 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n37 16.1731
R10760 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n28 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n27 16.1731
R10761 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n18 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n17 16.1731
R10762 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n55 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n51 16.077
R10763 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n39 SUNSAR_SAR8B_CV_0.XA20.CPO 15.2303
R10764 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n29 SUNSAR_SAR8B_CV_0.XA20.CPO 15.2303
R10765 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n19 SUNSAR_SAR8B_CV_0.XA20.CPO 15.2303
R10766 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n9 SUNSAR_SAR8B_CV_0.XA20.CPO 15.2303
R10767 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n59 SUNSAR_SAR8B_CV_0.XA20.CPO 13.6005
R10768 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n42 SUNSAR_SAR8B_CV_0.XA20.CPO 13.5534
R10769 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n32 SUNSAR_SAR8B_CV_0.XA20.CPO 13.5534
R10770 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n22 SUNSAR_SAR8B_CV_0.XA20.CPO 13.5534
R10771 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n12 SUNSAR_SAR8B_CV_0.XA20.CPO 13.5534
R10772 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n52 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n51 12.8005
R10773 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n37 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n36 12.8005
R10774 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n27 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n26 12.8005
R10775 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n17 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n16 12.8005
R10776 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n53 SUNSAR_SAR8B_CV_0.XA20.CPO 10.633
R10777 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n34 SUNSAR_SAR8B_CV_0.XA20.CPO 10.633
R10778 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n24 SUNSAR_SAR8B_CV_0.XA20.CPO 10.633
R10779 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n14 SUNSAR_SAR8B_CV_0.XA20.CPO 10.633
R10780 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n57 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n8 9.39659
R10781 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n43 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n42 9.39269
R10782 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n33 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n32 9.39269
R10783 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n23 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n22 9.39269
R10784 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n13 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n12 9.39269
R10785 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n58 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n57 9.39269
R10786 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n54 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n52 9.3005
R10787 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n36 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n35 9.3005
R10788 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n26 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n25 9.3005
R10789 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n16 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n15 9.3005
R10790 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n8 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n1 8.53383
R10791 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n44 SUNSAR_SAR8B_CV_0.XA20.CPO 8.063
R10792 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n49 8.063
R10793 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n40 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n39 7.7768
R10794 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n30 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n29 7.7768
R10795 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n20 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n19 7.7768
R10796 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n10 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n9 7.7768
R10797 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n48 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n47 7.61815
R10798 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n46 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n45 7.61815
R10799 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n52 SUNSAR_SAR8B_CV_0.XA20.CPO 7.52991
R10800 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n36 SUNSAR_SAR8B_CV_0.XA20.CPO 7.52991
R10801 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n26 SUNSAR_SAR8B_CV_0.XA20.CPO 7.52991
R10802 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n16 SUNSAR_SAR8B_CV_0.XA20.CPO 7.52991
R10803 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n42 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n41 6.77697
R10804 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n32 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n31 6.77697
R10805 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n22 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n21 6.77697
R10806 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n12 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n11 6.77697
R10807 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n57 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n56 6.41644
R10808 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n54 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n53 6.25297
R10809 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n35 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n34 6.25297
R10810 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n25 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n24 6.25297
R10811 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n15 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n14 6.25297
R10812 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n59 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n58 5.02011
R10813 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n58 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n1 4.51815
R10814 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n56 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n55 4.5005
R10815 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n54 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n50 4.5005
R10816 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n59 4.01619
R10817 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n43 2.32453
R10818 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n38 2.32453
R10819 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n33 2.32453
R10820 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n28 2.32453
R10821 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n23 2.32453
R10822 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n18 2.32453
R10823 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n13 2.32453
R10824 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n49 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n48 1.64756
R10825 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n47 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n46 1.64756
R10826 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n45 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n44 1.64756
R10827 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n44 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10828 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n45 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10829 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n46 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10830 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n47 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10831 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n48 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10832 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n49 SUNSAR_SAR8B_CV_0.XA20.CPO 0.445353
R10833 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n55 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n54 0.191676
R10834 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n56 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n50 0.191676
R10835 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n43 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n40 0.0965882
R10836 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n33 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n30 0.0965882
R10837 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n23 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n20 0.0965882
R10838 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n13 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n10 0.0965882
R10839 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n38 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n35 0.0926928
R10840 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n28 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n25 0.0926928
R10841 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n18 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n15 0.0926928
R10842 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n50 SUNSAR_SAR8B_CV_0.XA20.CPO 0.0740294
R10843 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t3 1060.4
R10844 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t8 1060.4
R10845 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t9 1060.4
R10846 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t7 1060.4
R10847 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n2 568.956
R10848 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t4 568.956
R10849 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n4 568.956
R10850 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t2 568.956
R10851 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t6 568.956
R10852 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n7 568.956
R10853 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t5 568.956
R10854 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n1 568.956
R10855 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t1 356.344
R10856 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.D SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.t0 151.719
R10857 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.D 128.754
R10858 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n8 97.8829
R10859 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n2 20.3299
R10860 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA1.XA2.MN3.G 20.3299
R10861 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA1.XA2.MP3.G 20.3299
R10862 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n1 20.3299
R10863 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n3 20.3299
R10864 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA1.XA2.MP2.G 20.3299
R10865 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA1.XA2.MN2.G 20.3299
R10866 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA1.XA2.MN0.G 20.3299
R10867 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n6 20.3299
R10868 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n5 20.3299
R10869 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA1.XA2.MN1.G 20.3299
R10870 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA1.XA2.MP1.G 20.3299
R10871 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n1 20.3299
R10872 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA1.XA2.MP0.G 20.3299
R10873 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n0 20.3299
R10874 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t12 1060.4
R10875 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t11 1060.4
R10876 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t14 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t8 1060.4
R10877 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t15 1060.4
R10878 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t12 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n1 568.956
R10879 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t9 568.956
R10880 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t11 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n3 568.956
R10881 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t13 568.956
R10882 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t14 568.956
R10883 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n6 568.956
R10884 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t10 568.956
R10885 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n0 568.956
R10886 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n14 292.5
R10887 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n19 292.5
R10888 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 197.272
R10889 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n17 112.829
R10890 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n15 111.059
R10891 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n18 111.059
R10892 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n12 92.5005
R10893 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t5 63.8431
R10894 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t7 63.8431
R10895 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t4 63.8431
R10896 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t6 63.8431
R10897 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n16 53.4593
R10898 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n9 45.4094
R10899 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t2 38.8894
R10900 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t0 38.8894
R10901 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t1 38.8894
R10902 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t3 38.8894
R10903 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n1 20.3299
R10904 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10905 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10906 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n0 20.3299
R10907 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n2 20.3299
R10908 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10909 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10910 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10911 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n5 20.3299
R10912 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n4 20.3299
R10913 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10914 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10915 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n0 20.3299
R10916 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n13 20.3299
R10917 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 20.3299
R10918 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n20 20.3299
R10919 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 17.6946
R10920 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 17.6946
R10921 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 12.325
R10922 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 12.323
R10923 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n11 10.6647
R10924 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n8 7.91541
R10925 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n10 7.89196
R10926 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n7 5.39616
R10927 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.168144
R10928 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.024
R10929 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t8 568.956
R10930 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t9 568.956
R10931 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n0 312.829
R10932 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n3 297.865
R10933 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n1 92.5005
R10934 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n16 92.5005
R10935 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n18 90.7299
R10936 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 81.6946
R10937 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t7 63.8431
R10938 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t3 63.8431
R10939 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t1 63.8431
R10940 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t5 63.8431
R10941 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n15 50.928
R10942 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t2 38.8894
R10943 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t6 38.8894
R10944 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t0 38.8894
R10945 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.t4 38.8894
R10946 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n17 38.024
R10947 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n2 31.624
R10948 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n14 28.5591
R10949 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 20.3299
R10950 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n4 20.3299
R10951 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 20.3299
R10952 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 20.3299
R10953 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10954 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10955 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10956 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10957 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10958 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 19.5486
R10959 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n6 13.7377
R10960 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n7 10.6968
R10961 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 10.633
R10962 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 8.72926
R10963 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n5 5.42812
R10964 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n8 4.12548
R10965 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n13 1.10785
R10966 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n12 1.10785
R10967 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n11 1.10785
R10968 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n10 1.10785
R10969 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n9 1.10785
R10970 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.168144
R10971 SUNSAR_SAR8B_CV_0.D<3>.t11 SUNSAR_SAR8B_CV_0.D<3>.t9 1060.4
R10972 SUNSAR_SAR8B_CV_0.D<3>.t9 SUNSAR_SAR8B_CV_0.D<3> 589.284
R10973 SUNSAR_SAR8B_CV_0.D<3>.n10 SUNSAR_SAR8B_CV_0.D<3>.t11 573.85
R10974 SUNSAR_SAR8B_CV_0.D<3>.n5 SUNSAR_SAR8B_CV_0.D<3>.t10 568.956
R10975 SUNSAR_SAR8B_CV_0.D<3>.n4 SUNSAR_SAR8B_CV_0.D<3>.t8 568.956
R10976 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<3>.n0 312.829
R10977 SUNSAR_SAR8B_CV_0.D<3>.n7 SUNSAR_SAR8B_CV_0.D<3>.n3 297.865
R10978 SUNSAR_SAR8B_CV_0.D<3>.n2 SUNSAR_SAR8B_CV_0.D<3>.n1 92.5005
R10979 SUNSAR_SAR8B_CV_0.D<3>.n23 SUNSAR_SAR8B_CV_0.D<3>.n22 92.5005
R10980 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<3>.n24 90.7299
R10981 SUNSAR_SAR8B_CV_0.D<3>.n8 SUNSAR_SAR8B_CV_0.D<3> 81.6946
R10982 SUNSAR_SAR8B_CV_0.D<3>.n3 SUNSAR_SAR8B_CV_0.D<3>.t4 63.8431
R10983 SUNSAR_SAR8B_CV_0.D<3>.n3 SUNSAR_SAR8B_CV_0.D<3>.t7 63.8431
R10984 SUNSAR_SAR8B_CV_0.D<3>.n0 SUNSAR_SAR8B_CV_0.D<3>.t0 63.8431
R10985 SUNSAR_SAR8B_CV_0.D<3>.n0 SUNSAR_SAR8B_CV_0.D<3>.t6 63.8431
R10986 SUNSAR_SAR8B_CV_0.D<3>.n24 SUNSAR_SAR8B_CV_0.D<3>.n21 48.7856
R10987 SUNSAR_SAR8B_CV_0.D<3>.n22 SUNSAR_SAR8B_CV_0.D<3>.t5 38.8894
R10988 SUNSAR_SAR8B_CV_0.D<3>.n22 SUNSAR_SAR8B_CV_0.D<3>.t1 38.8894
R10989 SUNSAR_SAR8B_CV_0.D<3>.n1 SUNSAR_SAR8B_CV_0.D<3>.t2 38.8894
R10990 SUNSAR_SAR8B_CV_0.D<3>.n1 SUNSAR_SAR8B_CV_0.D<3>.t3 38.8894
R10991 SUNSAR_SAR8B_CV_0.D<3>.n24 SUNSAR_SAR8B_CV_0.D<3>.n23 38.024
R10992 SUNSAR_SAR8B_CV_0.D<3>.n8 SUNSAR_SAR8B_CV_0.D<3>.n2 31.624
R10993 SUNSAR_SAR8B_CV_0.D<3>.n16 SUNSAR_SAR8B_CV_0.D<3>.n15 23.6453
R10994 SUNSAR_SAR8B_CV_0.D<3>.n15 SUNSAR_SAR8B_CV_0.D<3> 21.9678
R10995 SUNSAR_SAR8B_CV_0.D<3>.n4 SUNSAR_SAR8B_CV_0.D<3> 20.3299
R10996 SUNSAR_SAR8B_CV_0.D<3>.n5 SUNSAR_SAR8B_CV_0.D<3>.n4 20.3299
R10997 SUNSAR_SAR8B_CV_0.D<3>.n2 SUNSAR_SAR8B_CV_0.D<3> 20.3299
R10998 SUNSAR_SAR8B_CV_0.D<3>.n23 SUNSAR_SAR8B_CV_0.D<3> 20.3299
R10999 SUNSAR_SAR8B_CV_0.D<3>.n19 SUNSAR_SAR8B_CV_0.D<3>.n8 17.9961
R11000 SUNSAR_SAR8B_CV_0.D<3>.n14 SUNSAR_SAR8B_CV_0.D<3>.n13 16.9417
R11001 SUNSAR_SAR8B_CV_0.D<3>.n7 SUNSAR_SAR8B_CV_0.D<3>.n6 13.7377
R11002 SUNSAR_SAR8B_CV_0.D<3>.n10 SUNSAR_SAR8B_CV_0.D<3> 12.939
R11003 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<3>.n7 10.6968
R11004 SUNSAR_SAR8B_CV_0.D<3>.n6 SUNSAR_SAR8B_CV_0.D<3> 10.633
R11005 SUNSAR_SAR8B_CV_0.D<3>.n12 SUNSAR_SAR8B_CV_0.D<3>.n10 10.4477
R11006 SUNSAR_SAR8B_CV_0.D<3>.n21 SUNSAR_SAR8B_CV_0.D<3>.n20 9.3005
R11007 SUNSAR_SAR8B_CV_0.D<3>.n21 SUNSAR_SAR8B_CV_0.D<3>.n8 8.11757
R11008 SUNSAR_SAR8B_CV_0.D<3>.n6 SUNSAR_SAR8B_CV_0.D<3>.n5 5.42812
R11009 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<3>.n16 5.16471
R11010 SUNSAR_SAR8B_CV_0.D<3>.n20 SUNSAR_SAR8B_CV_0.D<3>.n9 4.5005
R11011 SUNSAR_SAR8B_CV_0.D<3>.n19 SUNSAR_SAR8B_CV_0.D<3>.n18 4.5005
R11012 SUNSAR_SAR8B_CV_0.D<3>.n14 SUNSAR_SAR8B_CV_0.D<3>.n9 3.4105
R11013 SUNSAR_SAR8B_CV_0.D<3>.n18 SUNSAR_SAR8B_CV_0.D<3>.n17 3.4105
R11014 SUNSAR_SAR8B_CV_0.D<3>.n13 SUNSAR_SAR8B_CV_0.D<3> 0.329788
R11015 SUNSAR_SAR8B_CV_0.D<3>.n18 SUNSAR_SAR8B_CV_0.D<3>.n9 0.191676
R11016 SUNSAR_SAR8B_CV_0.D<3>.n20 SUNSAR_SAR8B_CV_0.D<3>.n19 0.191676
R11017 SUNSAR_SAR8B_CV_0.D<3>.n15 SUNSAR_SAR8B_CV_0.D<3> 0.168144
R11018 SUNSAR_SAR8B_CV_0.D<3>.n11 SUNSAR_SAR8B_CV_0.D<3> 0.132853
R11019 SUNSAR_SAR8B_CV_0.D<3>.n11 SUNSAR_SAR8B_CV_0.D<3> 0.108934
R11020 SUNSAR_SAR8B_CV_0.D<3>.n17 SUNSAR_SAR8B_CV_0.D<3>.n14 0.0723824
R11021 SUNSAR_SAR8B_CV_0.D<3>.n12 SUNSAR_SAR8B_CV_0.D<3>.n11 0.0547169
R11022 SUNSAR_SAR8B_CV_0.D<3>.n17 SUNSAR_SAR8B_CV_0.D<3> 0.0281471
R11023 SUNSAR_SAR8B_CV_0.D<3>.n16 SUNSAR_SAR8B_CV_0.D<3> 0.00726261
R11024 SUNSAR_SAR8B_CV_0.D<3>.n13 SUNSAR_SAR8B_CV_0.D<3>.n12 0.00351205
R11025 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t16 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t17 1060.4
R11026 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t6 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t11 1060.4
R11027 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t17 SUNSAR_SAR8B_CV_0.XA20.XA11.MN0.G 589.284
R11028 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t11 SUNSAR_CAPT8B_CV_0.XA5a.MP0.G 589.284
R11029 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n4 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t16 574.351
R11030 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n8 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t21 568.956
R11031 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n6 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t8 568.956
R11032 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n7 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t4 568.956
R11033 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n3 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t18 568.956
R11034 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n13 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t5 568.956
R11035 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n11 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t15 568.956
R11036 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n12 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t22 568.956
R11037 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n10 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t25 568.956
R11038 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n18 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t3 568.956
R11039 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n16 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t33 568.956
R11040 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n17 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t2 568.956
R11041 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n15 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t19 568.956
R11042 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n23 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t23 568.956
R11043 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n21 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t37 568.956
R11044 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n22 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t14 568.956
R11045 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n20 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t7 568.956
R11046 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n28 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t30 568.956
R11047 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n26 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t26 568.956
R11048 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n27 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t29 568.956
R11049 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n25 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t12 568.956
R11050 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n33 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t24 568.956
R11051 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n31 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t32 568.956
R11052 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n32 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t31 568.956
R11053 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n30 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t9 568.956
R11054 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n38 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t20 568.956
R11055 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n36 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t10 568.956
R11056 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n37 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t13 568.956
R11057 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n35 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t34 568.956
R11058 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n43 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t36 568.956
R11059 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n41 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t28 568.956
R11060 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n42 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t27 568.956
R11061 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n40 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t35 568.956
R11062 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n0 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t6 568.956
R11063 SUNSAR_CAPT8B_CV_0.XA5.XA2.MP0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE.t1 376.673
R11064 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n1 SUNSAR_SAR8B_CV_0.CK_SAMPLE.t0 131.389
R11065 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n2 SUNSAR_CAPT8B_CV_0.XA5.XA2.MP0.D 121.977
R11066 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n55 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n0 90.7299
R11067 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n52 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n51 32.1954
R11068 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n7 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n6 20.3299
R11069 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n7 SUNSAR_SAR8B_CV_0.XA7.XA6.MN2.G 20.3299
R11070 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n3 SUNSAR_SAR8B_CV_0.XA7.XA6.MN0.G 20.3299
R11071 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n8 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n3 20.3299
R11072 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n8 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n7 20.3299
R11073 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n11 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.G 20.3299
R11074 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n12 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n11 20.3299
R11075 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n12 SUNSAR_SAR8B_CV_0.XA6.XA6.MN2.G 20.3299
R11076 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n10 SUNSAR_SAR8B_CV_0.XA6.XA6.MN0.G 20.3299
R11077 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n13 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n10 20.3299
R11078 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n13 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n12 20.3299
R11079 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n16 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.G 20.3299
R11080 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n17 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n16 20.3299
R11081 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n17 SUNSAR_SAR8B_CV_0.XA5.XA6.MN2.G 20.3299
R11082 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n15 SUNSAR_SAR8B_CV_0.XA5.XA6.MN0.G 20.3299
R11083 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n18 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n15 20.3299
R11084 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n18 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n17 20.3299
R11085 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n21 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.G 20.3299
R11086 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n22 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n21 20.3299
R11087 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n22 SUNSAR_SAR8B_CV_0.XA4.XA6.MN2.G 20.3299
R11088 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n20 SUNSAR_SAR8B_CV_0.XA4.XA6.MN0.G 20.3299
R11089 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n23 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n20 20.3299
R11090 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n23 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n22 20.3299
R11091 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n26 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.G 20.3299
R11092 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n27 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n26 20.3299
R11093 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n27 SUNSAR_SAR8B_CV_0.XA3.XA6.MN2.G 20.3299
R11094 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n25 SUNSAR_SAR8B_CV_0.XA3.XA6.MN0.G 20.3299
R11095 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n28 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n25 20.3299
R11096 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n28 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n27 20.3299
R11097 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n31 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.G 20.3299
R11098 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n32 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n31 20.3299
R11099 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n32 SUNSAR_SAR8B_CV_0.XA2.XA6.MN2.G 20.3299
R11100 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n30 SUNSAR_SAR8B_CV_0.XA2.XA6.MN0.G 20.3299
R11101 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n33 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n30 20.3299
R11102 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n33 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n32 20.3299
R11103 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n36 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.G 20.3299
R11104 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n37 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n36 20.3299
R11105 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n37 SUNSAR_SAR8B_CV_0.XA1.XA6.MN2.G 20.3299
R11106 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n35 SUNSAR_SAR8B_CV_0.XA1.XA6.MN0.G 20.3299
R11107 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n38 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n35 20.3299
R11108 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n38 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n37 20.3299
R11109 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n41 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.G 20.3299
R11110 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n42 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n41 20.3299
R11111 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n42 SUNSAR_SAR8B_CV_0.XA0.XA6.MN2.G 20.3299
R11112 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n40 SUNSAR_SAR8B_CV_0.XA0.XA6.MN0.G 20.3299
R11113 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n43 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n40 20.3299
R11114 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n43 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n42 20.3299
R11115 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n0 SUNSAR_CAPT8B_CV_0.XA5a.MN0.G 20.3299
R11116 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n5 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n4 19.6062
R11117 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n45 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n44 14.1335
R11118 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n54 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n1 12.8005
R11119 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n4 SUNSAR_SAR8B_CV_0.XA20.XA11.MP0.G 10.6653
R11120 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n5 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.G 10.6653
R11121 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n9 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.G 10.664
R11122 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n14 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.G 10.664
R11123 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n19 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.G 10.664
R11124 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n24 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.G 10.664
R11125 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n29 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.G 10.664
R11126 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n34 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.G 10.664
R11127 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n39 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.G 10.664
R11128 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n44 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.G 10.664
R11129 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n54 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n53 9.39659
R11130 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n53 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n2 9.39269
R11131 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n51 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n50 7.67697
R11132 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n49 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n48 7.67697
R11133 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n47 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n46 7.67697
R11134 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n2 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n1 6.77697
R11135 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n51 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n9 6.45708
R11136 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n50 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n14 6.45708
R11137 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n49 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n19 6.45708
R11138 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n48 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n24 6.45708
R11139 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n47 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n29 6.45708
R11140 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n46 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n34 6.45708
R11141 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n45 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n39 6.45708
R11142 SUNSAR_CAPT8B_CV_0.XA5.XA2.MN0.D SUNSAR_SAR8B_CV_0.CK_SAMPLE.n55 5.64756
R11143 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n9 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n8 5.39681
R11144 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n14 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n13 5.39681
R11145 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n19 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n18 5.39681
R11146 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n24 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n23 5.39681
R11147 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n29 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n28 5.39681
R11148 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n34 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n33 5.39681
R11149 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n39 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n38 5.39681
R11150 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n44 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n43 5.39681
R11151 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n6 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n5 5.39551
R11152 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n53 SUNSAR_CAPT8B_CV_0.CK_SAMPLE 4.83188
R11153 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n55 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n54 1.88285
R11154 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n50 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n49 1.58874
R11155 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n48 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n47 1.58874
R11156 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n46 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n45 1.58874
R11157 SUNSAR_CAPT8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.CK_SAMPLE.n52 0.140206
R11158 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n52 SUNSAR_CAPT8B_CV_0.CK_SAMPLE 0.122295
R11159 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t5 1060.4
R11160 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t6 1060.4
R11161 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t3 1060.4
R11162 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t9 1060.4
R11163 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n3 568.956
R11164 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t4 568.956
R11165 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n5 568.956
R11166 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t7 568.956
R11167 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t2 568.956
R11168 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n8 568.956
R11169 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t8 568.956
R11170 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n2 568.956
R11171 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.D SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t0 376.673
R11172 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.t1 131.389
R11173 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.D 121.977
R11174 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n3 20.3299
R11175 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA0.XA4.MP3.G 20.3299
R11176 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA0.XA4.MN3.G 20.3299
R11177 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n2 20.3299
R11178 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n4 20.3299
R11179 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA0.XA4.MN2.G 20.3299
R11180 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA0.XA4.MP2.G 20.3299
R11181 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA0.XA4.MP0.G 20.3299
R11182 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n7 20.3299
R11183 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n6 20.3299
R11184 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA0.XA4.MP1.G 20.3299
R11185 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA0.XA4.MN1.G 20.3299
R11186 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n2 20.3299
R11187 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n0 12.8005
R11188 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA0.XA4.MN0.G 10.6968
R11189 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n1 9.49168
R11190 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n10 9.47055
R11191 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n11 9.3005
R11192 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n12 7.52991
R11193 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n0 6.77697
R11194 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n9 5.36434
R11195 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t10 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t13 1060.4
R11196 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t11 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t12 1060.4
R11197 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t14 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t9 1060.4
R11198 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t15 1060.4
R11199 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t13 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n16 568.956
R11200 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t10 568.956
R11201 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t12 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n18 568.956
R11202 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n19 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t11 568.956
R11203 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n22 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t14 568.956
R11204 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n21 568.956
R11205 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n20 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t8 568.956
R11206 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t15 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n15 568.956
R11207 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n0 312.829
R11208 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n10 312.829
R11209 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n22 197.272
R11210 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n1 92.5005
R11211 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n13 92.5005
R11212 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 90.7299
R11213 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t4 63.8431
R11214 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t5 63.8431
R11215 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t6 63.8431
R11216 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t7 63.8431
R11217 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 61.177
R11218 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n3 53.4593
R11219 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n9 49.4935
R11220 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t0 38.8894
R11221 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t2 38.8894
R11222 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t1 38.8894
R11223 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t3 38.8894
R11224 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n2 38.024
R11225 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n12 38.024
R11226 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n11 29.5534
R11227 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11228 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n19 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n16 20.3299
R11229 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11230 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11231 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n15 20.3299
R11232 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n17 20.3299
R11233 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n18 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11234 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n19 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11235 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11236 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n20 20.3299
R11237 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n20 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n19 20.3299
R11238 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n20 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11239 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11240 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n22 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n15 20.3299
R11241 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n22 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 20.3299
R11242 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n14 20.3299
R11243 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11244 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11245 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11246 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11247 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11248 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 19.8942
R11249 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 10.3476
R11250 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n8 1.10785
R11251 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n7 1.10785
R11252 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n6 1.10785
R11253 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n5 1.10785
R11254 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n4 1.10785
R11255 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.168144
R11256 clk.t0 clk.t1 1060.4
R11257 clk.t1 clk 589.284
R11258 clk.n0 clk.t0 574.351
R11259 clk.n0 clk 10.6647
R11260 clk.n1 clk.n0 9.99729
R11261 clk.n1 clk 9.98704
R11262 clk clk.n1 0.0958824
R11263 SUNSAR_SAR8B_CV_0.XA3.CN1.t9 SUNSAR_SAR8B_CV_0.XA3.CN1.t12 1060.4
R11264 SUNSAR_SAR8B_CV_0.XA3.CN1.t15 SUNSAR_SAR8B_CV_0.XA3.CN1.t13 1060.4
R11265 SUNSAR_SAR8B_CV_0.XA3.CN1.t14 SUNSAR_SAR8B_CV_0.XA3.CN1.t10 1060.4
R11266 SUNSAR_SAR8B_CV_0.XA3.CN1.t8 SUNSAR_SAR8B_CV_0.XA3.CN1.t11 1060.4
R11267 SUNSAR_SAR8B_CV_0.XA3.CN1.t12 SUNSAR_SAR8B_CV_0.XA3.CN1.n5 568.956
R11268 SUNSAR_SAR8B_CV_0.XA3.CN1.n6 SUNSAR_SAR8B_CV_0.XA3.CN1.t9 568.956
R11269 SUNSAR_SAR8B_CV_0.XA3.CN1.t13 SUNSAR_SAR8B_CV_0.XA3.CN1.n7 568.956
R11270 SUNSAR_SAR8B_CV_0.XA3.CN1.n8 SUNSAR_SAR8B_CV_0.XA3.CN1.t15 568.956
R11271 SUNSAR_SAR8B_CV_0.XA3.CN1.n11 SUNSAR_SAR8B_CV_0.XA3.CN1.t14 568.956
R11272 SUNSAR_SAR8B_CV_0.XA3.CN1.t10 SUNSAR_SAR8B_CV_0.XA3.CN1.n10 568.956
R11273 SUNSAR_SAR8B_CV_0.XA3.CN1.n9 SUNSAR_SAR8B_CV_0.XA3.CN1.t8 568.956
R11274 SUNSAR_SAR8B_CV_0.XA3.CN1.t11 SUNSAR_SAR8B_CV_0.XA3.CN1.n4 568.956
R11275 SUNSAR_SAR8B_CV_0.XA3.CN1.n2 SUNSAR_SAR8B_CV_0.XA3.CN1.n1 292.5
R11276 SUNSAR_SAR8B_CV_0.XA3.CN1.n17 SUNSAR_SAR8B_CV_0.XA3.CN1.n16 292.5
R11277 SUNSAR_SAR8B_CV_0.XA3.CN1.n14 SUNSAR_SAR8B_CV_0.XA3.CN1 197.272
R11278 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.CN1.n0 112.829
R11279 SUNSAR_SAR8B_CV_0.XA3.CN1.n3 SUNSAR_SAR8B_CV_0.XA3.CN1.n2 111.059
R11280 SUNSAR_SAR8B_CV_0.XA3.CN1.n17 SUNSAR_SAR8B_CV_0.XA3.CN1.n15 111.059
R11281 SUNSAR_SAR8B_CV_0.XA3.CN1.n14 SUNSAR_SAR8B_CV_0.XA3.CN1.n13 92.5005
R11282 SUNSAR_SAR8B_CV_0.XA3.CN1.n16 SUNSAR_SAR8B_CV_0.XA3.CN1.t2 63.8431
R11283 SUNSAR_SAR8B_CV_0.XA3.CN1.n16 SUNSAR_SAR8B_CV_0.XA3.CN1.t5 63.8431
R11284 SUNSAR_SAR8B_CV_0.XA3.CN1.n1 SUNSAR_SAR8B_CV_0.XA3.CN1.t6 63.8431
R11285 SUNSAR_SAR8B_CV_0.XA3.CN1.n1 SUNSAR_SAR8B_CV_0.XA3.CN1.t7 63.8431
R11286 SUNSAR_SAR8B_CV_0.XA3.CN1.n15 SUNSAR_SAR8B_CV_0.XA3.CN1.n3 53.4593
R11287 SUNSAR_SAR8B_CV_0.XA3.CN1.n0 SUNSAR_SAR8B_CV_0.XA3.CN1.t1 38.8894
R11288 SUNSAR_SAR8B_CV_0.XA3.CN1.n0 SUNSAR_SAR8B_CV_0.XA3.CN1.t4 38.8894
R11289 SUNSAR_SAR8B_CV_0.XA3.CN1.n13 SUNSAR_SAR8B_CV_0.XA3.CN1.t3 38.8894
R11290 SUNSAR_SAR8B_CV_0.XA3.CN1.n13 SUNSAR_SAR8B_CV_0.XA3.CN1.t0 38.8894
R11291 SUNSAR_SAR8B_CV_0.XA3.CN1.n8 SUNSAR_SAR8B_CV_0.XA3.CN1.n5 20.3299
R11292 SUNSAR_SAR8B_CV_0.XA3.CN1.n5 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11293 SUNSAR_SAR8B_CV_0.XA3.CN1.n6 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11294 SUNSAR_SAR8B_CV_0.XA3.CN1.n7 SUNSAR_SAR8B_CV_0.XA3.CN1.n4 20.3299
R11295 SUNSAR_SAR8B_CV_0.XA3.CN1.n7 SUNSAR_SAR8B_CV_0.XA3.CN1.n6 20.3299
R11296 SUNSAR_SAR8B_CV_0.XA3.CN1.n7 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11297 SUNSAR_SAR8B_CV_0.XA3.CN1.n8 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11298 SUNSAR_SAR8B_CV_0.XA3.CN1.n10 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11299 SUNSAR_SAR8B_CV_0.XA3.CN1.n10 SUNSAR_SAR8B_CV_0.XA3.CN1.n9 20.3299
R11300 SUNSAR_SAR8B_CV_0.XA3.CN1.n9 SUNSAR_SAR8B_CV_0.XA3.CN1.n8 20.3299
R11301 SUNSAR_SAR8B_CV_0.XA3.CN1.n9 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11302 SUNSAR_SAR8B_CV_0.XA3.CN1.n4 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11303 SUNSAR_SAR8B_CV_0.XA3.CN1.n11 SUNSAR_SAR8B_CV_0.XA3.CN1.n4 20.3299
R11304 SUNSAR_SAR8B_CV_0.XA3.CN1.n2 SUNSAR_SAR8B_CV_0.XA3.CN1 20.3299
R11305 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.CN1.n14 20.3299
R11306 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.CN1.n17 20.3299
R11307 SUNSAR_SAR8B_CV_0.XA3.CN1.n3 SUNSAR_SAR8B_CV_0.XA3.CN1 17.6946
R11308 SUNSAR_SAR8B_CV_0.XA3.CN1.n15 SUNSAR_SAR8B_CV_0.XA3.CN1 17.6946
R11309 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.CN1.n12 10.6647
R11310 SUNSAR_SAR8B_CV_0.XA3.CN1.n12 SUNSAR_SAR8B_CV_0.XA3.CN1 7.91546
R11311 SUNSAR_SAR8B_CV_0.XA3.CN1.n12 SUNSAR_SAR8B_CV_0.XA3.CN1.n11 5.39616
R11312 SUNSAR_SAR8B_CV_0.D<4>.t11 SUNSAR_SAR8B_CV_0.D<4>.t10 1060.4
R11313 SUNSAR_SAR8B_CV_0.D<4>.t10 SUNSAR_SAR8B_CV_0.D<4> 589.284
R11314 SUNSAR_SAR8B_CV_0.D<4>.n16 SUNSAR_SAR8B_CV_0.D<4>.t11 573.85
R11315 SUNSAR_SAR8B_CV_0.D<4>.n4 SUNSAR_SAR8B_CV_0.D<4>.t8 568.956
R11316 SUNSAR_SAR8B_CV_0.D<4>.n3 SUNSAR_SAR8B_CV_0.D<4>.t9 568.956
R11317 SUNSAR_SAR8B_CV_0.D<4>.n2 SUNSAR_SAR8B_CV_0.D<4>.n1 292.5
R11318 SUNSAR_SAR8B_CV_0.D<4>.n11 SUNSAR_SAR8B_CV_0.D<4>.n10 292.5
R11319 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<4>.n9 112.829
R11320 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<4>.n0 112.829
R11321 SUNSAR_SAR8B_CV_0.D<4>.n12 SUNSAR_SAR8B_CV_0.D<4>.n11 111.059
R11322 SUNSAR_SAR8B_CV_0.D<4>.n26 SUNSAR_SAR8B_CV_0.D<4>.n8 89.224
R11323 SUNSAR_SAR8B_CV_0.D<4>.n1 SUNSAR_SAR8B_CV_0.D<4>.t7 63.8431
R11324 SUNSAR_SAR8B_CV_0.D<4>.n1 SUNSAR_SAR8B_CV_0.D<4>.t4 63.8431
R11325 SUNSAR_SAR8B_CV_0.D<4>.n10 SUNSAR_SAR8B_CV_0.D<4>.t6 63.8431
R11326 SUNSAR_SAR8B_CV_0.D<4>.n10 SUNSAR_SAR8B_CV_0.D<4>.t5 63.8431
R11327 SUNSAR_SAR8B_CV_0.D<4>.n13 SUNSAR_SAR8B_CV_0.D<4>.n12 48.7856
R11328 SUNSAR_SAR8B_CV_0.D<4>.n9 SUNSAR_SAR8B_CV_0.D<4>.t2 38.8894
R11329 SUNSAR_SAR8B_CV_0.D<4>.n9 SUNSAR_SAR8B_CV_0.D<4>.t0 38.8894
R11330 SUNSAR_SAR8B_CV_0.D<4>.n0 SUNSAR_SAR8B_CV_0.D<4>.t1 38.8894
R11331 SUNSAR_SAR8B_CV_0.D<4>.n0 SUNSAR_SAR8B_CV_0.D<4>.t3 38.8894
R11332 SUNSAR_SAR8B_CV_0.D<4>.n22 SUNSAR_SAR8B_CV_0.D<4>.n21 26.1435
R11333 SUNSAR_SAR8B_CV_0.D<4>.n21 SUNSAR_SAR8B_CV_0.D<4> 21.6222
R11334 SUNSAR_SAR8B_CV_0.D<4>.n3 SUNSAR_SAR8B_CV_0.D<4> 20.3299
R11335 SUNSAR_SAR8B_CV_0.D<4>.n4 SUNSAR_SAR8B_CV_0.D<4>.n3 20.3299
R11336 SUNSAR_SAR8B_CV_0.D<4>.n11 SUNSAR_SAR8B_CV_0.D<4> 20.3299
R11337 SUNSAR_SAR8B_CV_0.D<4>.n26 SUNSAR_SAR8B_CV_0.D<4>.n25 17.9961
R11338 SUNSAR_SAR8B_CV_0.D<4>.n12 SUNSAR_SAR8B_CV_0.D<4> 17.6946
R11339 SUNSAR_SAR8B_CV_0.D<4>.n20 SUNSAR_SAR8B_CV_0.D<4>.n19 17.0314
R11340 SUNSAR_SAR8B_CV_0.D<4>.n5 SUNSAR_SAR8B_CV_0.D<4> 15.2303
R11341 SUNSAR_SAR8B_CV_0.D<4>.n6 SUNSAR_SAR8B_CV_0.D<4> 13.5534
R11342 SUNSAR_SAR8B_CV_0.D<4>.n16 SUNSAR_SAR8B_CV_0.D<4> 12.939
R11343 SUNSAR_SAR8B_CV_0.D<4>.n8 SUNSAR_SAR8B_CV_0.D<4>.n2 12.8005
R11344 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<4>.n26 11.2946
R11345 SUNSAR_SAR8B_CV_0.D<4>.n7 SUNSAR_SAR8B_CV_0.D<4>.n5 11.2842
R11346 SUNSAR_SAR8B_CV_0.D<4>.n18 SUNSAR_SAR8B_CV_0.D<4>.n16 10.4477
R11347 SUNSAR_SAR8B_CV_0.D<4>.n8 SUNSAR_SAR8B_CV_0.D<4>.n7 9.49168
R11348 SUNSAR_SAR8B_CV_0.D<4>.n7 SUNSAR_SAR8B_CV_0.D<4>.n6 9.3005
R11349 SUNSAR_SAR8B_CV_0.D<4>.n14 SUNSAR_SAR8B_CV_0.D<4>.n13 9.3005
R11350 SUNSAR_SAR8B_CV_0.D<4>.n26 SUNSAR_SAR8B_CV_0.D<4>.n13 8.11757
R11351 SUNSAR_SAR8B_CV_0.D<4>.n6 SUNSAR_SAR8B_CV_0.D<4>.n2 6.77697
R11352 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<4>.n22 5.29327
R11353 SUNSAR_SAR8B_CV_0.D<4>.n15 SUNSAR_SAR8B_CV_0.D<4>.n14 4.5005
R11354 SUNSAR_SAR8B_CV_0.D<4>.n25 SUNSAR_SAR8B_CV_0.D<4>.n24 4.5005
R11355 SUNSAR_SAR8B_CV_0.D<4>.n5 SUNSAR_SAR8B_CV_0.D<4>.n4 3.90429
R11356 SUNSAR_SAR8B_CV_0.D<4>.n20 SUNSAR_SAR8B_CV_0.D<4>.n15 3.4105
R11357 SUNSAR_SAR8B_CV_0.D<4>.n24 SUNSAR_SAR8B_CV_0.D<4>.n23 3.4105
R11358 SUNSAR_SAR8B_CV_0.D<4>.n19 SUNSAR_SAR8B_CV_0.D<4> 0.337141
R11359 SUNSAR_SAR8B_CV_0.D<4>.n24 SUNSAR_SAR8B_CV_0.D<4>.n15 0.191676
R11360 SUNSAR_SAR8B_CV_0.D<4>.n25 SUNSAR_SAR8B_CV_0.D<4>.n14 0.191676
R11361 SUNSAR_SAR8B_CV_0.D<4>.n21 SUNSAR_SAR8B_CV_0.D<4> 0.168144
R11362 SUNSAR_SAR8B_CV_0.D<4>.n17 SUNSAR_SAR8B_CV_0.D<4> 0.136529
R11363 SUNSAR_SAR8B_CV_0.D<4>.n17 SUNSAR_SAR8B_CV_0.D<4> 0.111946
R11364 SUNSAR_SAR8B_CV_0.D<4>.n23 SUNSAR_SAR8B_CV_0.D<4>.n20 0.0713406
R11365 SUNSAR_SAR8B_CV_0.D<4>.n18 SUNSAR_SAR8B_CV_0.D<4>.n17 0.0517048
R11366 SUNSAR_SAR8B_CV_0.D<4>.n23 SUNSAR_SAR8B_CV_0.D<4> 0.0277464
R11367 SUNSAR_SAR8B_CV_0.D<4>.n19 SUNSAR_SAR8B_CV_0.D<4>.n18 0.00953614
R11368 SUNSAR_SAR8B_CV_0.D<4>.n22 SUNSAR_SAR8B_CV_0.D<4> 0.00726261
R11369 SUNSAR_SAR8B_CV_0.D<7>.t8 SUNSAR_SAR8B_CV_0.D<7>.t17 1060.4
R11370 SUNSAR_SAR8B_CV_0.D<7>.t13 SUNSAR_SAR8B_CV_0.D<7>.t14 1060.4
R11371 SUNSAR_SAR8B_CV_0.D<7>.t16 SUNSAR_SAR8B_CV_0.D<7>.t15 1060.4
R11372 SUNSAR_SAR8B_CV_0.D<7>.t9 SUNSAR_SAR8B_CV_0.D<7>.t10 1060.4
R11373 SUNSAR_SAR8B_CV_0.D<7>.t12 SUNSAR_SAR8B_CV_0.D<7>.t11 1060.4
R11374 SUNSAR_SAR8B_CV_0.D<7>.t11 SUNSAR_SAR8B_CV_0.D<7> 589.284
R11375 SUNSAR_SAR8B_CV_0.D<7>.n11 SUNSAR_SAR8B_CV_0.D<7>.t12 573.85
R11376 SUNSAR_SAR8B_CV_0.D<7>.t17 SUNSAR_SAR8B_CV_0.D<7>.n3 568.956
R11377 SUNSAR_SAR8B_CV_0.D<7>.n4 SUNSAR_SAR8B_CV_0.D<7>.t8 568.956
R11378 SUNSAR_SAR8B_CV_0.D<7>.t14 SUNSAR_SAR8B_CV_0.D<7>.n5 568.956
R11379 SUNSAR_SAR8B_CV_0.D<7>.n6 SUNSAR_SAR8B_CV_0.D<7>.t13 568.956
R11380 SUNSAR_SAR8B_CV_0.D<7>.n9 SUNSAR_SAR8B_CV_0.D<7>.t16 568.956
R11381 SUNSAR_SAR8B_CV_0.D<7>.t15 SUNSAR_SAR8B_CV_0.D<7>.n8 568.956
R11382 SUNSAR_SAR8B_CV_0.D<7>.n7 SUNSAR_SAR8B_CV_0.D<7>.t9 568.956
R11383 SUNSAR_SAR8B_CV_0.D<7>.t10 SUNSAR_SAR8B_CV_0.D<7>.n2 568.956
R11384 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<7>.n1 312.829
R11385 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<7>.n0 312.829
R11386 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<7>.n32 184.471
R11387 SUNSAR_SAR8B_CV_0.D<7>.n34 SUNSAR_SAR8B_CV_0.D<7>.n33 92.5005
R11388 SUNSAR_SAR8B_CV_0.D<7>.n37 SUNSAR_SAR8B_CV_0.D<7>.n36 92.5005
R11389 SUNSAR_SAR8B_CV_0.D<7>.n35 SUNSAR_SAR8B_CV_0.D<7> 90.7299
R11390 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<7>.n38 90.7299
R11391 SUNSAR_SAR8B_CV_0.D<7>.n0 SUNSAR_SAR8B_CV_0.D<7>.t6 63.8431
R11392 SUNSAR_SAR8B_CV_0.D<7>.n0 SUNSAR_SAR8B_CV_0.D<7>.t3 63.8431
R11393 SUNSAR_SAR8B_CV_0.D<7>.n1 SUNSAR_SAR8B_CV_0.D<7>.t4 63.8431
R11394 SUNSAR_SAR8B_CV_0.D<7>.n1 SUNSAR_SAR8B_CV_0.D<7>.t5 63.8431
R11395 SUNSAR_SAR8B_CV_0.D<7>.n38 SUNSAR_SAR8B_CV_0.D<7>.n35 53.4593
R11396 SUNSAR_SAR8B_CV_0.D<7>.n33 SUNSAR_SAR8B_CV_0.D<7>.t1 38.8894
R11397 SUNSAR_SAR8B_CV_0.D<7>.n33 SUNSAR_SAR8B_CV_0.D<7>.t7 38.8894
R11398 SUNSAR_SAR8B_CV_0.D<7>.n36 SUNSAR_SAR8B_CV_0.D<7>.t2 38.8894
R11399 SUNSAR_SAR8B_CV_0.D<7>.n36 SUNSAR_SAR8B_CV_0.D<7>.t0 38.8894
R11400 SUNSAR_SAR8B_CV_0.D<7>.n35 SUNSAR_SAR8B_CV_0.D<7>.n34 38.024
R11401 SUNSAR_SAR8B_CV_0.D<7>.n38 SUNSAR_SAR8B_CV_0.D<7>.n37 38.024
R11402 SUNSAR_SAR8B_CV_0.D<7>.n28 SUNSAR_SAR8B_CV_0.D<7>.n27 30.5203
R11403 SUNSAR_SAR8B_CV_0.D<7>.n6 SUNSAR_SAR8B_CV_0.D<7>.n3 20.3299
R11404 SUNSAR_SAR8B_CV_0.D<7>.n3 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11405 SUNSAR_SAR8B_CV_0.D<7>.n4 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11406 SUNSAR_SAR8B_CV_0.D<7>.n5 SUNSAR_SAR8B_CV_0.D<7>.n2 20.3299
R11407 SUNSAR_SAR8B_CV_0.D<7>.n5 SUNSAR_SAR8B_CV_0.D<7>.n4 20.3299
R11408 SUNSAR_SAR8B_CV_0.D<7>.n5 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11409 SUNSAR_SAR8B_CV_0.D<7>.n6 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11410 SUNSAR_SAR8B_CV_0.D<7>.n8 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11411 SUNSAR_SAR8B_CV_0.D<7>.n8 SUNSAR_SAR8B_CV_0.D<7>.n7 20.3299
R11412 SUNSAR_SAR8B_CV_0.D<7>.n7 SUNSAR_SAR8B_CV_0.D<7>.n6 20.3299
R11413 SUNSAR_SAR8B_CV_0.D<7>.n7 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11414 SUNSAR_SAR8B_CV_0.D<7>.n2 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11415 SUNSAR_SAR8B_CV_0.D<7>.n9 SUNSAR_SAR8B_CV_0.D<7>.n2 20.3299
R11416 SUNSAR_SAR8B_CV_0.D<7>.n34 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11417 SUNSAR_SAR8B_CV_0.D<7>.n37 SUNSAR_SAR8B_CV_0.D<7> 20.3299
R11418 SUNSAR_SAR8B_CV_0.D<7>.n10 SUNSAR_SAR8B_CV_0.D<7> 13.5534
R11419 SUNSAR_SAR8B_CV_0.D<7>.n11 SUNSAR_SAR8B_CV_0.D<7> 12.939
R11420 SUNSAR_SAR8B_CV_0.D<7>.n32 SUNSAR_SAR8B_CV_0.D<7>.n9 12.8005
R11421 SUNSAR_SAR8B_CV_0.D<7>.n16 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11422 SUNSAR_SAR8B_CV_0.D<7>.n18 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11423 SUNSAR_SAR8B_CV_0.D<7>.n20 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11424 SUNSAR_SAR8B_CV_0.D<7>.n22 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11425 SUNSAR_SAR8B_CV_0.D<7>.n24 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11426 SUNSAR_SAR8B_CV_0.D<7>.n26 SUNSAR_SAR8B_CV_0.D<7> 12.325
R11427 SUNSAR_SAR8B_CV_0.D<7>.n16 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11428 SUNSAR_SAR8B_CV_0.D<7>.n18 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11429 SUNSAR_SAR8B_CV_0.D<7>.n20 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11430 SUNSAR_SAR8B_CV_0.D<7>.n22 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11431 SUNSAR_SAR8B_CV_0.D<7>.n24 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11432 SUNSAR_SAR8B_CV_0.D<7>.n26 SUNSAR_SAR8B_CV_0.D<7> 12.323
R11433 SUNSAR_SAR8B_CV_0.D<7>.n13 SUNSAR_SAR8B_CV_0.D<7>.n11 10.4661
R11434 SUNSAR_SAR8B_CV_0.D<7>.n32 SUNSAR_SAR8B_CV_0.D<7>.n31 9.39465
R11435 SUNSAR_SAR8B_CV_0.D<7>.n31 SUNSAR_SAR8B_CV_0.D<7>.n10 9.39462
R11436 SUNSAR_SAR8B_CV_0.D<7>.n30 SUNSAR_SAR8B_CV_0.D<7>.n15 8.89607
R11437 SUNSAR_SAR8B_CV_0.D<7>.n17 SUNSAR_SAR8B_CV_0.D<7>.n16 7.22423
R11438 SUNSAR_SAR8B_CV_0.D<7>.n19 SUNSAR_SAR8B_CV_0.D<7>.n18 7.22423
R11439 SUNSAR_SAR8B_CV_0.D<7>.n21 SUNSAR_SAR8B_CV_0.D<7>.n20 7.22423
R11440 SUNSAR_SAR8B_CV_0.D<7>.n23 SUNSAR_SAR8B_CV_0.D<7>.n22 7.22423
R11441 SUNSAR_SAR8B_CV_0.D<7>.n25 SUNSAR_SAR8B_CV_0.D<7>.n24 7.22423
R11442 SUNSAR_SAR8B_CV_0.D<7>.n27 SUNSAR_SAR8B_CV_0.D<7>.n26 7.22423
R11443 SUNSAR_SAR8B_CV_0.D<7>.n10 SUNSAR_SAR8B_CV_0.D<7>.n9 6.77697
R11444 SUNSAR_SAR8B_CV_0.D<7>.n29 SUNSAR_SAR8B_CV_0.D<7>.n28 4.60555
R11445 SUNSAR_SAR8B_CV_0.D<7>.n29 SUNSAR_SAR8B_CV_0.D<7> 4.4796
R11446 SUNSAR_SAR8B_CV_0.D<7>.n31 SUNSAR_SAR8B_CV_0.D<7>.n30 3.92279
R11447 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<7>.n29 1.39774
R11448 SUNSAR_SAR8B_CV_0.D<7>.n27 SUNSAR_SAR8B_CV_0.D<7>.n25 1.10785
R11449 SUNSAR_SAR8B_CV_0.D<7>.n25 SUNSAR_SAR8B_CV_0.D<7>.n23 1.10785
R11450 SUNSAR_SAR8B_CV_0.D<7>.n23 SUNSAR_SAR8B_CV_0.D<7>.n21 1.10785
R11451 SUNSAR_SAR8B_CV_0.D<7>.n21 SUNSAR_SAR8B_CV_0.D<7>.n19 1.10785
R11452 SUNSAR_SAR8B_CV_0.D<7>.n19 SUNSAR_SAR8B_CV_0.D<7>.n17 1.10785
R11453 SUNSAR_SAR8B_CV_0.D<7>.n14 SUNSAR_SAR8B_CV_0.D<7> 0.8505
R11454 SUNSAR_SAR8B_CV_0.D<7>.n14 SUNSAR_SAR8B_CV_0.D<7> 0.386864
R11455 SUNSAR_SAR8B_CV_0.D<7>.n12 SUNSAR_SAR8B_CV_0.D<7> 0.34488
R11456 SUNSAR_SAR8B_CV_0.D<7>.n12 SUNSAR_SAR8B_CV_0.D<7> 0.254071
R11457 SUNSAR_SAR8B_CV_0.D<7>.n17 SUNSAR_SAR8B_CV_0.D<7> 0.168144
R11458 SUNSAR_SAR8B_CV_0.D<7>.n15 SUNSAR_SAR8B_CV_0.D<7>.n13 0.10523
R11459 SUNSAR_SAR8B_CV_0.D<7>.n13 SUNSAR_SAR8B_CV_0.D<7>.n12 0.0579324
R11460 SUNSAR_SAR8B_CV_0.D<7>.n15 SUNSAR_SAR8B_CV_0.D<7>.n14 0.0511757
R11461 SUNSAR_SAR8B_CV_0.D<7>.n30 SUNSAR_SAR8B_CV_0.D<7> 0.0481912
R11462 SUNSAR_SAR8B_CV_0.D<7>.n14 SUNSAR_SAR8B_CV_0.D<7> 0.027527
R11463 SUNSAR_SAR8B_CV_0.D<7>.n30 SUNSAR_SAR8B_CV_0.D<7> 0.0233286
R11464 SUNSAR_SAR8B_CV_0.D<7>.n28 SUNSAR_SAR8B_CV_0.D<7> 0.00726261
R11465 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t13 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t12 1060.4
R11466 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t9 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t14 1060.4
R11467 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t15 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t10 1060.4
R11468 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t8 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t11 1060.4
R11469 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t12 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n3 568.956
R11470 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t13 568.956
R11471 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t14 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n5 568.956
R11472 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t9 568.956
R11473 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t15 568.956
R11474 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n8 568.956
R11475 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t8 568.956
R11476 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n2 568.956
R11477 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n1 312.829
R11478 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n0 312.829
R11479 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n21 184.471
R11480 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n23 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n22 92.5005
R11481 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n26 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n25 92.5005
R11482 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n24 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 90.7299
R11483 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n27 90.7299
R11484 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t1 63.8431
R11485 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t2 63.8431
R11486 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t7 63.8431
R11487 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t3 63.8431
R11488 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n27 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n24 53.4593
R11489 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n22 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t4 38.8894
R11490 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n22 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t6 38.8894
R11491 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n25 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t0 38.8894
R11492 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n25 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.t5 38.8894
R11493 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n24 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n23 38.024
R11494 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n27 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n26 38.024
R11495 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n18 32.5933
R11496 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n3 20.3299
R11497 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11498 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11499 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n2 20.3299
R11500 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n4 20.3299
R11501 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11502 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11503 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11504 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n7 20.3299
R11505 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n6 20.3299
R11506 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11507 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11508 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n2 20.3299
R11509 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n23 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11510 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n26 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 20.3299
R11511 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 13.5534
R11512 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n21 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n9 12.8005
R11513 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.325
R11514 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.325
R11515 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.325
R11516 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.325
R11517 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.323
R11518 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.323
R11519 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.323
R11520 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 12.323
R11521 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n21 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n20 9.39466
R11522 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n10 9.39462
R11523 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n11 8.60658
R11524 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n13 8.60658
R11525 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n15 8.60658
R11526 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n17 8.60658
R11527 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n9 6.77697
R11528 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n19 3.93187
R11529 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n14 2.21814
R11530 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n12 2.21814
R11531 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n16 1.10785
R11532 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.168144
R11533 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.024
R11534 SUNSAR_SAR8B_CV_0.D<5>.t11 SUNSAR_SAR8B_CV_0.D<5>.t9 1060.4
R11535 SUNSAR_SAR8B_CV_0.D<5>.t9 SUNSAR_SAR8B_CV_0.D<5> 589.284
R11536 SUNSAR_SAR8B_CV_0.D<5>.n10 SUNSAR_SAR8B_CV_0.D<5>.t11 573.85
R11537 SUNSAR_SAR8B_CV_0.D<5>.n5 SUNSAR_SAR8B_CV_0.D<5>.t8 568.956
R11538 SUNSAR_SAR8B_CV_0.D<5>.n4 SUNSAR_SAR8B_CV_0.D<5>.t10 568.956
R11539 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<5>.n0 312.829
R11540 SUNSAR_SAR8B_CV_0.D<5>.n7 SUNSAR_SAR8B_CV_0.D<5>.n3 297.865
R11541 SUNSAR_SAR8B_CV_0.D<5>.n2 SUNSAR_SAR8B_CV_0.D<5>.n1 92.5005
R11542 SUNSAR_SAR8B_CV_0.D<5>.n27 SUNSAR_SAR8B_CV_0.D<5>.n26 92.5005
R11543 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<5>.n28 90.7299
R11544 SUNSAR_SAR8B_CV_0.D<5>.n8 SUNSAR_SAR8B_CV_0.D<5> 81.6946
R11545 SUNSAR_SAR8B_CV_0.D<5>.n0 SUNSAR_SAR8B_CV_0.D<5>.t6 63.8431
R11546 SUNSAR_SAR8B_CV_0.D<5>.n0 SUNSAR_SAR8B_CV_0.D<5>.t4 63.8431
R11547 SUNSAR_SAR8B_CV_0.D<5>.n3 SUNSAR_SAR8B_CV_0.D<5>.t7 63.8431
R11548 SUNSAR_SAR8B_CV_0.D<5>.n3 SUNSAR_SAR8B_CV_0.D<5>.t5 63.8431
R11549 SUNSAR_SAR8B_CV_0.D<5>.n28 SUNSAR_SAR8B_CV_0.D<5>.n25 48.7856
R11550 SUNSAR_SAR8B_CV_0.D<5>.n1 SUNSAR_SAR8B_CV_0.D<5>.t1 38.8894
R11551 SUNSAR_SAR8B_CV_0.D<5>.n1 SUNSAR_SAR8B_CV_0.D<5>.t0 38.8894
R11552 SUNSAR_SAR8B_CV_0.D<5>.n26 SUNSAR_SAR8B_CV_0.D<5>.t3 38.8894
R11553 SUNSAR_SAR8B_CV_0.D<5>.n26 SUNSAR_SAR8B_CV_0.D<5>.t2 38.8894
R11554 SUNSAR_SAR8B_CV_0.D<5>.n28 SUNSAR_SAR8B_CV_0.D<5>.n27 38.024
R11555 SUNSAR_SAR8B_CV_0.D<5>.n8 SUNSAR_SAR8B_CV_0.D<5>.n2 31.624
R11556 SUNSAR_SAR8B_CV_0.D<5>.n20 SUNSAR_SAR8B_CV_0.D<5>.n19 21.9321
R11557 SUNSAR_SAR8B_CV_0.D<5>.n16 SUNSAR_SAR8B_CV_0.D<5> 20.931
R11558 SUNSAR_SAR8B_CV_0.D<5>.n17 SUNSAR_SAR8B_CV_0.D<5> 20.931
R11559 SUNSAR_SAR8B_CV_0.D<5>.n18 SUNSAR_SAR8B_CV_0.D<5> 20.931
R11560 SUNSAR_SAR8B_CV_0.D<5>.n19 SUNSAR_SAR8B_CV_0.D<5> 20.931
R11561 SUNSAR_SAR8B_CV_0.D<5>.n4 SUNSAR_SAR8B_CV_0.D<5> 20.3299
R11562 SUNSAR_SAR8B_CV_0.D<5>.n5 SUNSAR_SAR8B_CV_0.D<5>.n4 20.3299
R11563 SUNSAR_SAR8B_CV_0.D<5>.n2 SUNSAR_SAR8B_CV_0.D<5> 20.3299
R11564 SUNSAR_SAR8B_CV_0.D<5>.n27 SUNSAR_SAR8B_CV_0.D<5> 20.3299
R11565 SUNSAR_SAR8B_CV_0.D<5>.n23 SUNSAR_SAR8B_CV_0.D<5>.n8 17.9961
R11566 SUNSAR_SAR8B_CV_0.D<5>.n15 SUNSAR_SAR8B_CV_0.D<5>.n14 16.878
R11567 SUNSAR_SAR8B_CV_0.D<5>.n7 SUNSAR_SAR8B_CV_0.D<5>.n6 13.7377
R11568 SUNSAR_SAR8B_CV_0.D<5>.n10 SUNSAR_SAR8B_CV_0.D<5> 12.939
R11569 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<5>.n7 10.6968
R11570 SUNSAR_SAR8B_CV_0.D<5>.n6 SUNSAR_SAR8B_CV_0.D<5> 10.633
R11571 SUNSAR_SAR8B_CV_0.D<5>.n12 SUNSAR_SAR8B_CV_0.D<5>.n10 10.3282
R11572 SUNSAR_SAR8B_CV_0.D<5>.n25 SUNSAR_SAR8B_CV_0.D<5>.n24 9.3005
R11573 SUNSAR_SAR8B_CV_0.D<5>.n25 SUNSAR_SAR8B_CV_0.D<5>.n8 8.11757
R11574 SUNSAR_SAR8B_CV_0.D<5>.n6 SUNSAR_SAR8B_CV_0.D<5>.n5 5.42812
R11575 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<5>.n20 5.42183
R11576 SUNSAR_SAR8B_CV_0.D<5>.n24 SUNSAR_SAR8B_CV_0.D<5>.n9 4.5005
R11577 SUNSAR_SAR8B_CV_0.D<5>.n23 SUNSAR_SAR8B_CV_0.D<5>.n22 4.5005
R11578 SUNSAR_SAR8B_CV_0.D<5>.n15 SUNSAR_SAR8B_CV_0.D<5>.n9 3.4105
R11579 SUNSAR_SAR8B_CV_0.D<5>.n22 SUNSAR_SAR8B_CV_0.D<5>.n21 3.4105
R11580 SUNSAR_SAR8B_CV_0.D<5>.n18 SUNSAR_SAR8B_CV_0.D<5>.n17 2.21814
R11581 SUNSAR_SAR8B_CV_0.D<5>.n17 SUNSAR_SAR8B_CV_0.D<5>.n16 2.21814
R11582 SUNSAR_SAR8B_CV_0.D<5>.n19 SUNSAR_SAR8B_CV_0.D<5>.n18 1.10785
R11583 SUNSAR_SAR8B_CV_0.D<5>.n13 SUNSAR_SAR8B_CV_0.D<5> 0.315348
R11584 SUNSAR_SAR8B_CV_0.D<5>.n13 SUNSAR_SAR8B_CV_0.D<5> 0.247488
R11585 SUNSAR_SAR8B_CV_0.D<5>.n22 SUNSAR_SAR8B_CV_0.D<5>.n9 0.191676
R11586 SUNSAR_SAR8B_CV_0.D<5>.n24 SUNSAR_SAR8B_CV_0.D<5>.n23 0.191676
R11587 SUNSAR_SAR8B_CV_0.D<5>.n16 SUNSAR_SAR8B_CV_0.D<5> 0.168144
R11588 SUNSAR_SAR8B_CV_0.D<5>.n11 SUNSAR_SAR8B_CV_0.D<5> 0.136529
R11589 SUNSAR_SAR8B_CV_0.D<5>.n21 SUNSAR_SAR8B_CV_0.D<5>.n15 0.0723824
R11590 SUNSAR_SAR8B_CV_0.D<5>.n11 SUNSAR_SAR8B_CV_0.D<5> 0.063
R11591 SUNSAR_SAR8B_CV_0.D<5>.n12 SUNSAR_SAR8B_CV_0.D<5>.n11 0.0292162
R11592 SUNSAR_SAR8B_CV_0.D<5>.n21 SUNSAR_SAR8B_CV_0.D<5> 0.0281471
R11593 SUNSAR_SAR8B_CV_0.D<5>.n14 SUNSAR_SAR8B_CV_0.D<5>.n13 0.0270736
R11594 SUNSAR_SAR8B_CV_0.D<5>.n14 SUNSAR_SAR8B_CV_0.D<5>.n12 0.0194256
R11595 SUNSAR_SAR8B_CV_0.D<5>.n20 SUNSAR_SAR8B_CV_0.D<5> 0.00726261
R11596 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.G SUNSAR_SAR8B_CV_0.EN.t57 589.284
R11597 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.G SUNSAR_SAR8B_CV_0.EN.t12 589.284
R11598 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.G SUNSAR_SAR8B_CV_0.EN.t4 589.284
R11599 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.G SUNSAR_SAR8B_CV_0.EN.t35 589.284
R11600 SUNSAR_SAR8B_CV_0.EN.n6 SUNSAR_SAR8B_CV_0.EN.t29 574.383
R11601 SUNSAR_SAR8B_CV_0.EN.n10 SUNSAR_SAR8B_CV_0.EN.t41 568.956
R11602 SUNSAR_SAR8B_CV_0.EN.n3 SUNSAR_SAR8B_CV_0.EN.t19 568.956
R11603 SUNSAR_SAR8B_CV_0.EN.n21 SUNSAR_SAR8B_CV_0.EN.t59 568.956
R11604 SUNSAR_SAR8B_CV_0.EN.n19 SUNSAR_SAR8B_CV_0.EN.t15 568.956
R11605 SUNSAR_SAR8B_CV_0.EN.n20 SUNSAR_SAR8B_CV_0.EN.t7 568.956
R11606 SUNSAR_SAR8B_CV_0.EN.n13 SUNSAR_SAR8B_CV_0.EN.t5 568.956
R11607 SUNSAR_SAR8B_CV_0.EN.n16 SUNSAR_SAR8B_CV_0.EN.t18 568.956
R11608 SUNSAR_SAR8B_CV_0.EN.n14 SUNSAR_SAR8B_CV_0.EN.t9 568.956
R11609 SUNSAR_SAR8B_CV_0.EN.n15 SUNSAR_SAR8B_CV_0.EN.t54 568.956
R11610 SUNSAR_SAR8B_CV_0.EN.n29 SUNSAR_SAR8B_CV_0.EN.t31 568.956
R11611 SUNSAR_SAR8B_CV_0.EN.n27 SUNSAR_SAR8B_CV_0.EN.t43 568.956
R11612 SUNSAR_SAR8B_CV_0.EN.n28 SUNSAR_SAR8B_CV_0.EN.t26 568.956
R11613 SUNSAR_SAR8B_CV_0.EN.n32 SUNSAR_SAR8B_CV_0.EN.t13 568.956
R11614 SUNSAR_SAR8B_CV_0.EN.n30 SUNSAR_SAR8B_CV_0.EN.t33 568.956
R11615 SUNSAR_SAR8B_CV_0.EN.n31 SUNSAR_SAR8B_CV_0.EN.t14 568.956
R11616 SUNSAR_SAR8B_CV_0.EN.n47 SUNSAR_SAR8B_CV_0.EN.t58 568.956
R11617 SUNSAR_SAR8B_CV_0.EN.n45 SUNSAR_SAR8B_CV_0.EN.t21 568.956
R11618 SUNSAR_SAR8B_CV_0.EN.n46 SUNSAR_SAR8B_CV_0.EN.t34 568.956
R11619 SUNSAR_SAR8B_CV_0.EN.n39 SUNSAR_SAR8B_CV_0.EN.t56 568.956
R11620 SUNSAR_SAR8B_CV_0.EN.n42 SUNSAR_SAR8B_CV_0.EN.t32 568.956
R11621 SUNSAR_SAR8B_CV_0.EN.n40 SUNSAR_SAR8B_CV_0.EN.t3 568.956
R11622 SUNSAR_SAR8B_CV_0.EN.n41 SUNSAR_SAR8B_CV_0.EN.t24 568.956
R11623 SUNSAR_SAR8B_CV_0.EN.n55 SUNSAR_SAR8B_CV_0.EN.t22 568.956
R11624 SUNSAR_SAR8B_CV_0.EN.n53 SUNSAR_SAR8B_CV_0.EN.t38 568.956
R11625 SUNSAR_SAR8B_CV_0.EN.n54 SUNSAR_SAR8B_CV_0.EN.t23 568.956
R11626 SUNSAR_SAR8B_CV_0.EN.n58 SUNSAR_SAR8B_CV_0.EN.t44 568.956
R11627 SUNSAR_SAR8B_CV_0.EN.n56 SUNSAR_SAR8B_CV_0.EN.t40 568.956
R11628 SUNSAR_SAR8B_CV_0.EN.n57 SUNSAR_SAR8B_CV_0.EN.t51 568.956
R11629 SUNSAR_SAR8B_CV_0.EN.n73 SUNSAR_SAR8B_CV_0.EN.t10 568.956
R11630 SUNSAR_SAR8B_CV_0.EN.n71 SUNSAR_SAR8B_CV_0.EN.t36 568.956
R11631 SUNSAR_SAR8B_CV_0.EN.n72 SUNSAR_SAR8B_CV_0.EN.t49 568.956
R11632 SUNSAR_SAR8B_CV_0.EN.n65 SUNSAR_SAR8B_CV_0.EN.t17 568.956
R11633 SUNSAR_SAR8B_CV_0.EN.n68 SUNSAR_SAR8B_CV_0.EN.t39 568.956
R11634 SUNSAR_SAR8B_CV_0.EN.n66 SUNSAR_SAR8B_CV_0.EN.t37 568.956
R11635 SUNSAR_SAR8B_CV_0.EN.n67 SUNSAR_SAR8B_CV_0.EN.t50 568.956
R11636 SUNSAR_SAR8B_CV_0.EN.n81 SUNSAR_SAR8B_CV_0.EN.t28 568.956
R11637 SUNSAR_SAR8B_CV_0.EN.n79 SUNSAR_SAR8B_CV_0.EN.t46 568.956
R11638 SUNSAR_SAR8B_CV_0.EN.n80 SUNSAR_SAR8B_CV_0.EN.t60 568.956
R11639 SUNSAR_SAR8B_CV_0.EN.n84 SUNSAR_SAR8B_CV_0.EN.t11 568.956
R11640 SUNSAR_SAR8B_CV_0.EN.n82 SUNSAR_SAR8B_CV_0.EN.t20 568.956
R11641 SUNSAR_SAR8B_CV_0.EN.n83 SUNSAR_SAR8B_CV_0.EN.t55 568.956
R11642 SUNSAR_SAR8B_CV_0.EN.n99 SUNSAR_SAR8B_CV_0.EN.t25 568.956
R11643 SUNSAR_SAR8B_CV_0.EN.n97 SUNSAR_SAR8B_CV_0.EN.t2 568.956
R11644 SUNSAR_SAR8B_CV_0.EN.n98 SUNSAR_SAR8B_CV_0.EN.t53 568.956
R11645 SUNSAR_SAR8B_CV_0.EN.n91 SUNSAR_SAR8B_CV_0.EN.t45 568.956
R11646 SUNSAR_SAR8B_CV_0.EN.n94 SUNSAR_SAR8B_CV_0.EN.t47 568.956
R11647 SUNSAR_SAR8B_CV_0.EN.n92 SUNSAR_SAR8B_CV_0.EN.t27 568.956
R11648 SUNSAR_SAR8B_CV_0.EN.n93 SUNSAR_SAR8B_CV_0.EN.t52 568.956
R11649 SUNSAR_SAR8B_CV_0.EN.n107 SUNSAR_SAR8B_CV_0.EN.t16 568.956
R11650 SUNSAR_SAR8B_CV_0.EN.n105 SUNSAR_SAR8B_CV_0.EN.t48 568.956
R11651 SUNSAR_SAR8B_CV_0.EN.n106 SUNSAR_SAR8B_CV_0.EN.t30 568.956
R11652 SUNSAR_SAR8B_CV_0.EN.n110 SUNSAR_SAR8B_CV_0.EN.t42 568.956
R11653 SUNSAR_SAR8B_CV_0.EN.n108 SUNSAR_SAR8B_CV_0.EN.t8 568.956
R11654 SUNSAR_SAR8B_CV_0.EN.n109 SUNSAR_SAR8B_CV_0.EN.t6 568.956
R11655 SUNSAR_SAR8B_CV_0.EN.n17 SUNSAR_SAR8B_CV_0.EN.n13 422.776
R11656 SUNSAR_SAR8B_CV_0.EN.n43 SUNSAR_SAR8B_CV_0.EN.n39 422.776
R11657 SUNSAR_SAR8B_CV_0.EN.n69 SUNSAR_SAR8B_CV_0.EN.n65 422.776
R11658 SUNSAR_SAR8B_CV_0.EN.n95 SUNSAR_SAR8B_CV_0.EN.n91 422.776
R11659 SUNSAR_SAR8B_CV_0.EN.n33 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.G 402.447
R11660 SUNSAR_SAR8B_CV_0.EN.n59 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.G 402.447
R11661 SUNSAR_SAR8B_CV_0.EN.n85 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.G 402.447
R11662 SUNSAR_SAR8B_CV_0.EN.n111 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.G 402.447
R11663 SUNSAR_CAPT8B_CV_0.XA5a.MP0.D SUNSAR_SAR8B_CV_0.EN.t1 376.673
R11664 SUNSAR_SAR8B_CV_0.EN.n18 SUNSAR_SAR8B_CV_0.EN.n17 150.965
R11665 SUNSAR_SAR8B_CV_0.EN.n44 SUNSAR_SAR8B_CV_0.EN.n43 150.965
R11666 SUNSAR_SAR8B_CV_0.EN.n70 SUNSAR_SAR8B_CV_0.EN.n69 150.965
R11667 SUNSAR_SAR8B_CV_0.EN.n96 SUNSAR_SAR8B_CV_0.EN.n95 150.965
R11668 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.G SUNSAR_SAR8B_CV_0.EN.n33 137.412
R11669 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.G SUNSAR_SAR8B_CV_0.EN.n59 137.412
R11670 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.G SUNSAR_SAR8B_CV_0.EN.n85 137.412
R11671 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.G SUNSAR_SAR8B_CV_0.EN.n111 137.412
R11672 SUNSAR_SAR8B_CV_0.EN.n0 SUNSAR_SAR8B_CV_0.EN.t0 131.389
R11673 SUNSAR_SAR8B_CV_0.EN.n1 SUNSAR_CAPT8B_CV_0.XA5a.MP0.D 121.977
R11674 SUNSAR_SAR8B_CV_0.EN.n17 SUNSAR_SAR8B_CV_0.EN.n16 38.024
R11675 SUNSAR_SAR8B_CV_0.EN.n43 SUNSAR_SAR8B_CV_0.EN.n42 38.024
R11676 SUNSAR_SAR8B_CV_0.EN.n69 SUNSAR_SAR8B_CV_0.EN.n68 38.024
R11677 SUNSAR_SAR8B_CV_0.EN.n95 SUNSAR_SAR8B_CV_0.EN.n94 38.024
R11678 SUNSAR_CAPT8B_CV_0.EN SUNSAR_SAR8B_CV_0.EN.n115 35.7616
R11679 SUNSAR_SAR8B_CV_0.EN.n19 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP0.G 20.3299
R11680 SUNSAR_SAR8B_CV_0.EN.n20 SUNSAR_SAR8B_CV_0.EN.n19 20.3299
R11681 SUNSAR_SAR8B_CV_0.EN.n20 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.G 20.3299
R11682 SUNSAR_SAR8B_CV_0.EN.n21 SUNSAR_SAR8B_CV_0.EN.n20 20.3299
R11683 SUNSAR_SAR8B_CV_0.EN.n13 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP0.G 20.3299
R11684 SUNSAR_SAR8B_CV_0.EN.n14 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP0.G 20.3299
R11685 SUNSAR_SAR8B_CV_0.EN.n15 SUNSAR_SAR8B_CV_0.EN.n14 20.3299
R11686 SUNSAR_SAR8B_CV_0.EN.n15 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.G 20.3299
R11687 SUNSAR_SAR8B_CV_0.EN.n16 SUNSAR_SAR8B_CV_0.EN.n15 20.3299
R11688 SUNSAR_SAR8B_CV_0.EN.n16 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.G 20.3299
R11689 SUNSAR_SAR8B_CV_0.EN.n27 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP0.G 20.3299
R11690 SUNSAR_SAR8B_CV_0.EN.n28 SUNSAR_SAR8B_CV_0.EN.n27 20.3299
R11691 SUNSAR_SAR8B_CV_0.EN.n28 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.G 20.3299
R11692 SUNSAR_SAR8B_CV_0.EN.n29 SUNSAR_SAR8B_CV_0.EN.n28 20.3299
R11693 SUNSAR_SAR8B_CV_0.EN.n30 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP0.G 20.3299
R11694 SUNSAR_SAR8B_CV_0.EN.n31 SUNSAR_SAR8B_CV_0.EN.n30 20.3299
R11695 SUNSAR_SAR8B_CV_0.EN.n31 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.G 20.3299
R11696 SUNSAR_SAR8B_CV_0.EN.n32 SUNSAR_SAR8B_CV_0.EN.n31 20.3299
R11697 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.G SUNSAR_SAR8B_CV_0.EN.n32 20.3299
R11698 SUNSAR_SAR8B_CV_0.EN.n45 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP0.G 20.3299
R11699 SUNSAR_SAR8B_CV_0.EN.n46 SUNSAR_SAR8B_CV_0.EN.n45 20.3299
R11700 SUNSAR_SAR8B_CV_0.EN.n46 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.G 20.3299
R11701 SUNSAR_SAR8B_CV_0.EN.n47 SUNSAR_SAR8B_CV_0.EN.n46 20.3299
R11702 SUNSAR_SAR8B_CV_0.EN.n39 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP0.G 20.3299
R11703 SUNSAR_SAR8B_CV_0.EN.n40 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP0.G 20.3299
R11704 SUNSAR_SAR8B_CV_0.EN.n41 SUNSAR_SAR8B_CV_0.EN.n40 20.3299
R11705 SUNSAR_SAR8B_CV_0.EN.n41 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.G 20.3299
R11706 SUNSAR_SAR8B_CV_0.EN.n42 SUNSAR_SAR8B_CV_0.EN.n41 20.3299
R11707 SUNSAR_SAR8B_CV_0.EN.n42 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.G 20.3299
R11708 SUNSAR_SAR8B_CV_0.EN.n53 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP0.G 20.3299
R11709 SUNSAR_SAR8B_CV_0.EN.n54 SUNSAR_SAR8B_CV_0.EN.n53 20.3299
R11710 SUNSAR_SAR8B_CV_0.EN.n54 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.G 20.3299
R11711 SUNSAR_SAR8B_CV_0.EN.n55 SUNSAR_SAR8B_CV_0.EN.n54 20.3299
R11712 SUNSAR_SAR8B_CV_0.EN.n56 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP0.G 20.3299
R11713 SUNSAR_SAR8B_CV_0.EN.n57 SUNSAR_SAR8B_CV_0.EN.n56 20.3299
R11714 SUNSAR_SAR8B_CV_0.EN.n57 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.G 20.3299
R11715 SUNSAR_SAR8B_CV_0.EN.n58 SUNSAR_SAR8B_CV_0.EN.n57 20.3299
R11716 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.G SUNSAR_SAR8B_CV_0.EN.n58 20.3299
R11717 SUNSAR_SAR8B_CV_0.EN.n71 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP0.G 20.3299
R11718 SUNSAR_SAR8B_CV_0.EN.n72 SUNSAR_SAR8B_CV_0.EN.n71 20.3299
R11719 SUNSAR_SAR8B_CV_0.EN.n72 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.G 20.3299
R11720 SUNSAR_SAR8B_CV_0.EN.n73 SUNSAR_SAR8B_CV_0.EN.n72 20.3299
R11721 SUNSAR_SAR8B_CV_0.EN.n65 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP0.G 20.3299
R11722 SUNSAR_SAR8B_CV_0.EN.n66 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP0.G 20.3299
R11723 SUNSAR_SAR8B_CV_0.EN.n67 SUNSAR_SAR8B_CV_0.EN.n66 20.3299
R11724 SUNSAR_SAR8B_CV_0.EN.n67 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.G 20.3299
R11725 SUNSAR_SAR8B_CV_0.EN.n68 SUNSAR_SAR8B_CV_0.EN.n67 20.3299
R11726 SUNSAR_SAR8B_CV_0.EN.n68 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.G 20.3299
R11727 SUNSAR_SAR8B_CV_0.EN.n79 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP0.G 20.3299
R11728 SUNSAR_SAR8B_CV_0.EN.n80 SUNSAR_SAR8B_CV_0.EN.n79 20.3299
R11729 SUNSAR_SAR8B_CV_0.EN.n80 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.G 20.3299
R11730 SUNSAR_SAR8B_CV_0.EN.n81 SUNSAR_SAR8B_CV_0.EN.n80 20.3299
R11731 SUNSAR_SAR8B_CV_0.EN.n82 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP0.G 20.3299
R11732 SUNSAR_SAR8B_CV_0.EN.n83 SUNSAR_SAR8B_CV_0.EN.n82 20.3299
R11733 SUNSAR_SAR8B_CV_0.EN.n83 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.G 20.3299
R11734 SUNSAR_SAR8B_CV_0.EN.n84 SUNSAR_SAR8B_CV_0.EN.n83 20.3299
R11735 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.G SUNSAR_SAR8B_CV_0.EN.n84 20.3299
R11736 SUNSAR_SAR8B_CV_0.EN.n97 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP0.G 20.3299
R11737 SUNSAR_SAR8B_CV_0.EN.n98 SUNSAR_SAR8B_CV_0.EN.n97 20.3299
R11738 SUNSAR_SAR8B_CV_0.EN.n98 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.G 20.3299
R11739 SUNSAR_SAR8B_CV_0.EN.n99 SUNSAR_SAR8B_CV_0.EN.n98 20.3299
R11740 SUNSAR_SAR8B_CV_0.EN.n91 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP0.G 20.3299
R11741 SUNSAR_SAR8B_CV_0.EN.n92 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP0.G 20.3299
R11742 SUNSAR_SAR8B_CV_0.EN.n93 SUNSAR_SAR8B_CV_0.EN.n92 20.3299
R11743 SUNSAR_SAR8B_CV_0.EN.n93 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.G 20.3299
R11744 SUNSAR_SAR8B_CV_0.EN.n94 SUNSAR_SAR8B_CV_0.EN.n93 20.3299
R11745 SUNSAR_SAR8B_CV_0.EN.n94 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.G 20.3299
R11746 SUNSAR_SAR8B_CV_0.EN.n105 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP0.G 20.3299
R11747 SUNSAR_SAR8B_CV_0.EN.n106 SUNSAR_SAR8B_CV_0.EN.n105 20.3299
R11748 SUNSAR_SAR8B_CV_0.EN.n106 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.G 20.3299
R11749 SUNSAR_SAR8B_CV_0.EN.n107 SUNSAR_SAR8B_CV_0.EN.n106 20.3299
R11750 SUNSAR_SAR8B_CV_0.EN.n108 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP0.G 20.3299
R11751 SUNSAR_SAR8B_CV_0.EN.n109 SUNSAR_SAR8B_CV_0.EN.n108 20.3299
R11752 SUNSAR_SAR8B_CV_0.EN.n109 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.G 20.3299
R11753 SUNSAR_SAR8B_CV_0.EN.n110 SUNSAR_SAR8B_CV_0.EN.n109 20.3299
R11754 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.G SUNSAR_SAR8B_CV_0.EN.n110 20.3299
R11755 SUNSAR_SAR8B_CV_0.EN.n33 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.G 17.6946
R11756 SUNSAR_SAR8B_CV_0.EN.n59 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.G 17.6946
R11757 SUNSAR_SAR8B_CV_0.EN.n85 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.G 17.6946
R11758 SUNSAR_SAR8B_CV_0.EN.n111 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.G 17.6946
R11759 SUNSAR_SAR8B_CV_0.EN.n11 SUNSAR_SAR8B_CV_0.EN.n10 16.1692
R11760 SUNSAR_SAR8B_CV_0.EN.n3 SUNSAR_SAR8B_CV_0.EN.n2 16.1445
R11761 SUNSAR_SAR8B_CV_0.EN.n36 SUNSAR_SAR8B_CV_0.EN.n29 16.077
R11762 SUNSAR_SAR8B_CV_0.EN.n62 SUNSAR_SAR8B_CV_0.EN.n55 16.077
R11763 SUNSAR_SAR8B_CV_0.EN.n88 SUNSAR_SAR8B_CV_0.EN.n81 16.077
R11764 SUNSAR_SAR8B_CV_0.EN.n114 SUNSAR_SAR8B_CV_0.EN.n107 16.077
R11765 SUNSAR_SAR8B_CV_0.EN.n10 SUNSAR_SAR8B_CV_0.EN.n9 12.8005
R11766 SUNSAR_SAR8B_CV_0.EN.n4 SUNSAR_SAR8B_CV_0.EN.n3 12.8005
R11767 SUNSAR_SAR8B_CV_0.EN.n22 SUNSAR_SAR8B_CV_0.EN.n21 12.8005
R11768 SUNSAR_SAR8B_CV_0.EN.n34 SUNSAR_SAR8B_CV_0.EN.n29 12.8005
R11769 SUNSAR_SAR8B_CV_0.EN.n48 SUNSAR_SAR8B_CV_0.EN.n47 12.8005
R11770 SUNSAR_SAR8B_CV_0.EN.n60 SUNSAR_SAR8B_CV_0.EN.n55 12.8005
R11771 SUNSAR_SAR8B_CV_0.EN.n74 SUNSAR_SAR8B_CV_0.EN.n73 12.8005
R11772 SUNSAR_SAR8B_CV_0.EN.n86 SUNSAR_SAR8B_CV_0.EN.n81 12.8005
R11773 SUNSAR_SAR8B_CV_0.EN.n100 SUNSAR_SAR8B_CV_0.EN.n99 12.8005
R11774 SUNSAR_SAR8B_CV_0.EN.n112 SUNSAR_SAR8B_CV_0.EN.n107 12.8005
R11775 SUNSAR_SAR8B_CV_0.EN.n117 SUNSAR_SAR8B_CV_0.EN.n0 12.8005
R11776 SUNSAR_SAR8B_CV_0.EN.n6 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.G 10.633
R11777 SUNSAR_SAR8B_CV_0.EN.n117 SUNSAR_SAR8B_CV_0.EN.n116 9.39659
R11778 SUNSAR_SAR8B_CV_0.EN.n116 SUNSAR_SAR8B_CV_0.EN.n1 9.39269
R11779 SUNSAR_SAR8B_CV_0.EN.n5 SUNSAR_SAR8B_CV_0.EN.n4 9.3005
R11780 SUNSAR_SAR8B_CV_0.EN.n9 SUNSAR_SAR8B_CV_0.EN.n8 9.3005
R11781 SUNSAR_SAR8B_CV_0.EN.n24 SUNSAR_SAR8B_CV_0.EN.n18 9.3005
R11782 SUNSAR_SAR8B_CV_0.EN.n23 SUNSAR_SAR8B_CV_0.EN.n22 9.3005
R11783 SUNSAR_SAR8B_CV_0.EN.n35 SUNSAR_SAR8B_CV_0.EN.n34 9.3005
R11784 SUNSAR_SAR8B_CV_0.EN.n50 SUNSAR_SAR8B_CV_0.EN.n44 9.3005
R11785 SUNSAR_SAR8B_CV_0.EN.n49 SUNSAR_SAR8B_CV_0.EN.n48 9.3005
R11786 SUNSAR_SAR8B_CV_0.EN.n61 SUNSAR_SAR8B_CV_0.EN.n60 9.3005
R11787 SUNSAR_SAR8B_CV_0.EN.n76 SUNSAR_SAR8B_CV_0.EN.n70 9.3005
R11788 SUNSAR_SAR8B_CV_0.EN.n75 SUNSAR_SAR8B_CV_0.EN.n74 9.3005
R11789 SUNSAR_SAR8B_CV_0.EN.n87 SUNSAR_SAR8B_CV_0.EN.n86 9.3005
R11790 SUNSAR_SAR8B_CV_0.EN.n102 SUNSAR_SAR8B_CV_0.EN.n96 9.3005
R11791 SUNSAR_SAR8B_CV_0.EN.n101 SUNSAR_SAR8B_CV_0.EN.n100 9.3005
R11792 SUNSAR_SAR8B_CV_0.EN.n113 SUNSAR_SAR8B_CV_0.EN.n112 9.3005
R11793 SUNSAR_SAR8B_CV_0.EN.n9 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.G 7.52991
R11794 SUNSAR_SAR8B_CV_0.EN.n4 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN0.G 7.52991
R11795 SUNSAR_SAR8B_CV_0.EN.n22 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.G 7.52991
R11796 SUNSAR_SAR8B_CV_0.EN.n34 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.G 7.52991
R11797 SUNSAR_SAR8B_CV_0.EN.n48 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.G 7.52991
R11798 SUNSAR_SAR8B_CV_0.EN.n60 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.G 7.52991
R11799 SUNSAR_SAR8B_CV_0.EN.n74 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.G 7.52991
R11800 SUNSAR_SAR8B_CV_0.EN.n86 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.G 7.52991
R11801 SUNSAR_SAR8B_CV_0.EN.n100 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.G 7.52991
R11802 SUNSAR_SAR8B_CV_0.EN.n112 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.G 7.52991
R11803 SUNSAR_CAPT8B_CV_0.XA5a.MN0.D SUNSAR_SAR8B_CV_0.EN.n117 7.52991
R11804 SUNSAR_SAR8B_CV_0.EN.n90 SUNSAR_SAR8B_CV_0.EN.n89 7.48579
R11805 SUNSAR_SAR8B_CV_0.EN.n64 SUNSAR_SAR8B_CV_0.EN.n63 7.48579
R11806 SUNSAR_SAR8B_CV_0.EN.n38 SUNSAR_SAR8B_CV_0.EN.n37 7.48579
R11807 SUNSAR_SAR8B_CV_0.EN.n21 SUNSAR_SAR8B_CV_0.EN.n18 6.77697
R11808 SUNSAR_SAR8B_CV_0.EN.n47 SUNSAR_SAR8B_CV_0.EN.n44 6.77697
R11809 SUNSAR_SAR8B_CV_0.EN.n73 SUNSAR_SAR8B_CV_0.EN.n70 6.77697
R11810 SUNSAR_SAR8B_CV_0.EN.n99 SUNSAR_SAR8B_CV_0.EN.n96 6.77697
R11811 SUNSAR_SAR8B_CV_0.EN.n1 SUNSAR_SAR8B_CV_0.EN.n0 6.77697
R11812 SUNSAR_SAR8B_CV_0.EN.n12 SUNSAR_SAR8B_CV_0.EN.n11 5.10394
R11813 SUNSAR_SAR8B_CV_0.EN.n116 SUNSAR_CAPT8B_CV_0.EN 4.83188
R11814 SUNSAR_SAR8B_CV_0.EN.n115 SUNSAR_SAR8B_CV_0.EN.n114 4.5005
R11815 SUNSAR_SAR8B_CV_0.EN.n113 SUNSAR_SAR8B_CV_0.EN.n104 4.5005
R11816 SUNSAR_SAR8B_CV_0.EN.n103 SUNSAR_SAR8B_CV_0.EN.n102 4.5005
R11817 SUNSAR_SAR8B_CV_0.EN.n101 SUNSAR_SAR8B_CV_0.EN.n90 4.5005
R11818 SUNSAR_SAR8B_CV_0.EN.n89 SUNSAR_SAR8B_CV_0.EN.n88 4.5005
R11819 SUNSAR_SAR8B_CV_0.EN.n87 SUNSAR_SAR8B_CV_0.EN.n78 4.5005
R11820 SUNSAR_SAR8B_CV_0.EN.n77 SUNSAR_SAR8B_CV_0.EN.n76 4.5005
R11821 SUNSAR_SAR8B_CV_0.EN.n75 SUNSAR_SAR8B_CV_0.EN.n64 4.5005
R11822 SUNSAR_SAR8B_CV_0.EN.n63 SUNSAR_SAR8B_CV_0.EN.n62 4.5005
R11823 SUNSAR_SAR8B_CV_0.EN.n61 SUNSAR_SAR8B_CV_0.EN.n52 4.5005
R11824 SUNSAR_SAR8B_CV_0.EN.n51 SUNSAR_SAR8B_CV_0.EN.n50 4.5005
R11825 SUNSAR_SAR8B_CV_0.EN.n49 SUNSAR_SAR8B_CV_0.EN.n38 4.5005
R11826 SUNSAR_SAR8B_CV_0.EN.n37 SUNSAR_SAR8B_CV_0.EN.n36 4.5005
R11827 SUNSAR_SAR8B_CV_0.EN.n35 SUNSAR_SAR8B_CV_0.EN.n26 4.5005
R11828 SUNSAR_SAR8B_CV_0.EN.n25 SUNSAR_SAR8B_CV_0.EN.n24 4.5005
R11829 SUNSAR_SAR8B_CV_0.EN.n23 SUNSAR_SAR8B_CV_0.EN.n12 4.5005
R11830 SUNSAR_SAR8B_CV_0.EN.n7 SUNSAR_SAR8B_CV_0.EN.n6 4.19047
R11831 SUNSAR_SAR8B_CV_0.EN.n7 SUNSAR_SAR8B_CV_0.EN.n5 4.00418
R11832 SUNSAR_SAR8B_CV_0.EN.n2 SUNSAR_SAR8B_CV_0.XA0.EN 2.35274
R11833 SUNSAR_SAR8B_CV_0.EN.n8 SUNSAR_SAR8B_CV_0.EN.n7 1.41594
R11834 SUNSAR_SAR8B_CV_0.EN.n104 SUNSAR_SAR8B_CV_0.EN.n103 1.39756
R11835 SUNSAR_SAR8B_CV_0.EN.n78 SUNSAR_SAR8B_CV_0.EN.n77 1.39756
R11836 SUNSAR_SAR8B_CV_0.EN.n52 SUNSAR_SAR8B_CV_0.EN.n51 1.39756
R11837 SUNSAR_SAR8B_CV_0.EN.n26 SUNSAR_SAR8B_CV_0.EN.n25 1.39756
R11838 SUNSAR_SAR8B_CV_0.EN.n24 SUNSAR_SAR8B_CV_0.EN.n23 0.191676
R11839 SUNSAR_SAR8B_CV_0.EN.n36 SUNSAR_SAR8B_CV_0.EN.n35 0.191676
R11840 SUNSAR_SAR8B_CV_0.EN.n50 SUNSAR_SAR8B_CV_0.EN.n49 0.191676
R11841 SUNSAR_SAR8B_CV_0.EN.n62 SUNSAR_SAR8B_CV_0.EN.n61 0.191676
R11842 SUNSAR_SAR8B_CV_0.EN.n76 SUNSAR_SAR8B_CV_0.EN.n75 0.191676
R11843 SUNSAR_SAR8B_CV_0.EN.n88 SUNSAR_SAR8B_CV_0.EN.n87 0.191676
R11844 SUNSAR_SAR8B_CV_0.EN.n102 SUNSAR_SAR8B_CV_0.EN.n101 0.191676
R11845 SUNSAR_SAR8B_CV_0.EN.n114 SUNSAR_SAR8B_CV_0.EN.n113 0.191676
R11846 SUNSAR_SAR8B_CV_0.EN.n115 SUNSAR_SAR8B_CV_0.EN.n104 0.191676
R11847 SUNSAR_SAR8B_CV_0.EN.n103 SUNSAR_SAR8B_CV_0.EN.n90 0.191676
R11848 SUNSAR_SAR8B_CV_0.EN.n89 SUNSAR_SAR8B_CV_0.EN.n78 0.191676
R11849 SUNSAR_SAR8B_CV_0.EN.n77 SUNSAR_SAR8B_CV_0.EN.n64 0.191676
R11850 SUNSAR_SAR8B_CV_0.EN.n63 SUNSAR_SAR8B_CV_0.EN.n52 0.191676
R11851 SUNSAR_SAR8B_CV_0.EN.n51 SUNSAR_SAR8B_CV_0.EN.n38 0.191676
R11852 SUNSAR_SAR8B_CV_0.EN.n37 SUNSAR_SAR8B_CV_0.EN.n26 0.191676
R11853 SUNSAR_SAR8B_CV_0.EN.n25 SUNSAR_SAR8B_CV_0.EN.n12 0.191676
R11854 SUNSAR_SAR8B_CV_0.EN.n5 SUNSAR_SAR8B_CV_0.EN.n2 0.123303
R11855 SUNSAR_SAR8B_CV_0.EN.n11 SUNSAR_SAR8B_CV_0.EN.n8 0.0965882
R11856 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t4 1060.4
R11857 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t5 1060.4
R11858 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t9 1060.4
R11859 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t6 1060.4
R11860 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n1 568.956
R11861 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t8 568.956
R11862 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n3 568.956
R11863 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t2 568.956
R11864 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t7 568.956
R11865 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n6 568.956
R11866 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t3 568.956
R11867 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n0 568.956
R11868 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t0 356.344
R11869 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.t1 131.389
R11870 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n9 128.754
R11871 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA0.XA2.MP0.G 97.8829
R11872 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n1 20.3299
R11873 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA0.XA2.MN3.G 20.3299
R11874 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA0.XA2.MP3.G 20.3299
R11875 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n0 20.3299
R11876 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n2 20.3299
R11877 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA0.XA2.MP2.G 20.3299
R11878 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA0.XA2.MN2.G 20.3299
R11879 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA0.XA2.MN0.G 20.3299
R11880 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n5 20.3299
R11881 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n4 20.3299
R11882 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA0.XA2.MN1.G 20.3299
R11883 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA0.XA2.MP1.G 20.3299
R11884 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n0 20.3299
R11885 SUNSAR_SAR8B_CV_0.XA0.XA2.MP0.G SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n7 20.3299
R11886 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n8 20.3299
R11887 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.D 20.3299
R11888 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t9 1060.4
R11889 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t4 1060.4
R11890 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t5 1060.4
R11891 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t8 1060.4
R11892 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n2 568.956
R11893 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t3 568.956
R11894 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n4 568.956
R11895 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t2 568.956
R11896 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t6 568.956
R11897 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n7 568.956
R11898 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t7 568.956
R11899 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n1 568.956
R11900 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t0 356.344
R11901 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.D SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.t1 151.719
R11902 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.D 128.754
R11903 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n8 97.8829
R11904 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n2 20.3299
R11905 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA7.XA2.MN3.G 20.3299
R11906 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA7.XA2.MP3.G 20.3299
R11907 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n1 20.3299
R11908 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n3 20.3299
R11909 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA7.XA2.MP2.G 20.3299
R11910 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA7.XA2.MN2.G 20.3299
R11911 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA7.XA2.MN0.G 20.3299
R11912 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n6 20.3299
R11913 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n5 20.3299
R11914 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA7.XA2.MN1.G 20.3299
R11915 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA7.XA2.MP1.G 20.3299
R11916 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n1 20.3299
R11917 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA7.XA2.MP0.G 20.3299
R11918 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n0 20.3299
R11919 SUNSAR_SAR8B_CV_0.XA7.CN1.t15 SUNSAR_SAR8B_CV_0.XA7.CN1.t13 1060.4
R11920 SUNSAR_SAR8B_CV_0.XA7.CN1.t10 SUNSAR_SAR8B_CV_0.XA7.CN1.t11 1060.4
R11921 SUNSAR_SAR8B_CV_0.XA7.CN1.t9 SUNSAR_SAR8B_CV_0.XA7.CN1.t12 1060.4
R11922 SUNSAR_SAR8B_CV_0.XA7.CN1.t8 SUNSAR_SAR8B_CV_0.XA7.CN1.t14 1060.4
R11923 SUNSAR_SAR8B_CV_0.XA7.CN1.t13 SUNSAR_SAR8B_CV_0.XA7.CN1.n1 568.956
R11924 SUNSAR_SAR8B_CV_0.XA7.CN1.n2 SUNSAR_SAR8B_CV_0.XA7.CN1.t15 568.956
R11925 SUNSAR_SAR8B_CV_0.XA7.CN1.t11 SUNSAR_SAR8B_CV_0.XA7.CN1.n3 568.956
R11926 SUNSAR_SAR8B_CV_0.XA7.CN1.n4 SUNSAR_SAR8B_CV_0.XA7.CN1.t10 568.956
R11927 SUNSAR_SAR8B_CV_0.XA7.CN1.n7 SUNSAR_SAR8B_CV_0.XA7.CN1.t9 568.956
R11928 SUNSAR_SAR8B_CV_0.XA7.CN1.t12 SUNSAR_SAR8B_CV_0.XA7.CN1.n6 568.956
R11929 SUNSAR_SAR8B_CV_0.XA7.CN1.n5 SUNSAR_SAR8B_CV_0.XA7.CN1.t8 568.956
R11930 SUNSAR_SAR8B_CV_0.XA7.CN1.t14 SUNSAR_SAR8B_CV_0.XA7.CN1.n0 568.956
R11931 SUNSAR_SAR8B_CV_0.XA7.CN1.n12 SUNSAR_SAR8B_CV_0.XA7.CN1.n11 292.5
R11932 SUNSAR_SAR8B_CV_0.XA7.CN1.n17 SUNSAR_SAR8B_CV_0.XA7.CN1.n16 292.5
R11933 SUNSAR_SAR8B_CV_0.XA7.CN1.n10 SUNSAR_SAR8B_CV_0.XA7.CN1 197.272
R11934 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.CN1.n14 112.829
R11935 SUNSAR_SAR8B_CV_0.XA7.CN1.n13 SUNSAR_SAR8B_CV_0.XA7.CN1.n12 111.059
R11936 SUNSAR_SAR8B_CV_0.XA7.CN1.n17 SUNSAR_SAR8B_CV_0.XA7.CN1.n15 111.059
R11937 SUNSAR_SAR8B_CV_0.XA7.CN1.n10 SUNSAR_SAR8B_CV_0.XA7.CN1.n9 92.5005
R11938 SUNSAR_SAR8B_CV_0.XA7.CN1.n16 SUNSAR_SAR8B_CV_0.XA7.CN1.t5 63.8431
R11939 SUNSAR_SAR8B_CV_0.XA7.CN1.n16 SUNSAR_SAR8B_CV_0.XA7.CN1.t4 63.8431
R11940 SUNSAR_SAR8B_CV_0.XA7.CN1.n11 SUNSAR_SAR8B_CV_0.XA7.CN1.t7 63.8431
R11941 SUNSAR_SAR8B_CV_0.XA7.CN1.n11 SUNSAR_SAR8B_CV_0.XA7.CN1.t6 63.8431
R11942 SUNSAR_SAR8B_CV_0.XA7.CN1.n15 SUNSAR_SAR8B_CV_0.XA7.CN1.n13 53.4593
R11943 SUNSAR_SAR8B_CV_0.XA7.CN1.n9 SUNSAR_SAR8B_CV_0.XA7.CN1.t0 38.8894
R11944 SUNSAR_SAR8B_CV_0.XA7.CN1.n9 SUNSAR_SAR8B_CV_0.XA7.CN1.t2 38.8894
R11945 SUNSAR_SAR8B_CV_0.XA7.CN1.n14 SUNSAR_SAR8B_CV_0.XA7.CN1.t3 38.8894
R11946 SUNSAR_SAR8B_CV_0.XA7.CN1.n14 SUNSAR_SAR8B_CV_0.XA7.CN1.t1 38.8894
R11947 SUNSAR_SAR8B_CV_0.XA7.CN1.n4 SUNSAR_SAR8B_CV_0.XA7.CN1.n1 20.3299
R11948 SUNSAR_SAR8B_CV_0.XA7.CN1.n1 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11949 SUNSAR_SAR8B_CV_0.XA7.CN1.n2 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11950 SUNSAR_SAR8B_CV_0.XA7.CN1.n3 SUNSAR_SAR8B_CV_0.XA7.CN1.n0 20.3299
R11951 SUNSAR_SAR8B_CV_0.XA7.CN1.n3 SUNSAR_SAR8B_CV_0.XA7.CN1.n2 20.3299
R11952 SUNSAR_SAR8B_CV_0.XA7.CN1.n3 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11953 SUNSAR_SAR8B_CV_0.XA7.CN1.n4 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11954 SUNSAR_SAR8B_CV_0.XA7.CN1.n6 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11955 SUNSAR_SAR8B_CV_0.XA7.CN1.n6 SUNSAR_SAR8B_CV_0.XA7.CN1.n5 20.3299
R11956 SUNSAR_SAR8B_CV_0.XA7.CN1.n5 SUNSAR_SAR8B_CV_0.XA7.CN1.n4 20.3299
R11957 SUNSAR_SAR8B_CV_0.XA7.CN1.n5 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11958 SUNSAR_SAR8B_CV_0.XA7.CN1.n0 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11959 SUNSAR_SAR8B_CV_0.XA7.CN1.n7 SUNSAR_SAR8B_CV_0.XA7.CN1.n0 20.3299
R11960 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.CN1.n10 20.3299
R11961 SUNSAR_SAR8B_CV_0.XA7.CN1.n12 SUNSAR_SAR8B_CV_0.XA7.CN1 20.3299
R11962 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.CN1.n17 20.3299
R11963 SUNSAR_SAR8B_CV_0.XA7.CN1.n13 SUNSAR_SAR8B_CV_0.XA7.CN1 17.6946
R11964 SUNSAR_SAR8B_CV_0.XA7.CN1.n15 SUNSAR_SAR8B_CV_0.XA7.CN1 17.6946
R11965 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.CN1.n8 10.6647
R11966 SUNSAR_SAR8B_CV_0.XA7.CN1.n8 SUNSAR_SAR8B_CV_0.XA7.CN1 7.91546
R11967 SUNSAR_SAR8B_CV_0.XA7.CN1.n8 SUNSAR_SAR8B_CV_0.XA7.CN1.n7 5.39616
R11968 SUNSAR_SAR8B_CV_0.XA6.CN1.t13 SUNSAR_SAR8B_CV_0.XA6.CN1.t8 1060.4
R11969 SUNSAR_SAR8B_CV_0.XA6.CN1.t14 SUNSAR_SAR8B_CV_0.XA6.CN1.t9 1060.4
R11970 SUNSAR_SAR8B_CV_0.XA6.CN1.t11 SUNSAR_SAR8B_CV_0.XA6.CN1.t15 1060.4
R11971 SUNSAR_SAR8B_CV_0.XA6.CN1.t12 SUNSAR_SAR8B_CV_0.XA6.CN1.t10 1060.4
R11972 SUNSAR_SAR8B_CV_0.XA6.CN1.t8 SUNSAR_SAR8B_CV_0.XA6.CN1.n3 568.956
R11973 SUNSAR_SAR8B_CV_0.XA6.CN1.n4 SUNSAR_SAR8B_CV_0.XA6.CN1.t13 568.956
R11974 SUNSAR_SAR8B_CV_0.XA6.CN1.t9 SUNSAR_SAR8B_CV_0.XA6.CN1.n5 568.956
R11975 SUNSAR_SAR8B_CV_0.XA6.CN1.n6 SUNSAR_SAR8B_CV_0.XA6.CN1.t14 568.956
R11976 SUNSAR_SAR8B_CV_0.XA6.CN1.n9 SUNSAR_SAR8B_CV_0.XA6.CN1.t11 568.956
R11977 SUNSAR_SAR8B_CV_0.XA6.CN1.t15 SUNSAR_SAR8B_CV_0.XA6.CN1.n8 568.956
R11978 SUNSAR_SAR8B_CV_0.XA6.CN1.n7 SUNSAR_SAR8B_CV_0.XA6.CN1.t12 568.956
R11979 SUNSAR_SAR8B_CV_0.XA6.CN1.t10 SUNSAR_SAR8B_CV_0.XA6.CN1.n2 568.956
R11980 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.CN1.n1 312.829
R11981 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.CN1.n0 312.829
R11982 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.CN1.n12 184.471
R11983 SUNSAR_SAR8B_CV_0.XA6.CN1.n14 SUNSAR_SAR8B_CV_0.XA6.CN1.n13 92.5005
R11984 SUNSAR_SAR8B_CV_0.XA6.CN1.n17 SUNSAR_SAR8B_CV_0.XA6.CN1.n16 92.5005
R11985 SUNSAR_SAR8B_CV_0.XA6.CN1.n15 SUNSAR_SAR8B_CV_0.XA6.CN1 90.7299
R11986 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.CN1.n18 90.7299
R11987 SUNSAR_SAR8B_CV_0.XA6.CN1.n1 SUNSAR_SAR8B_CV_0.XA6.CN1.t5 63.8431
R11988 SUNSAR_SAR8B_CV_0.XA6.CN1.n1 SUNSAR_SAR8B_CV_0.XA6.CN1.t6 63.8431
R11989 SUNSAR_SAR8B_CV_0.XA6.CN1.n0 SUNSAR_SAR8B_CV_0.XA6.CN1.t2 63.8431
R11990 SUNSAR_SAR8B_CV_0.XA6.CN1.n0 SUNSAR_SAR8B_CV_0.XA6.CN1.t0 63.8431
R11991 SUNSAR_SAR8B_CV_0.XA6.CN1.n18 SUNSAR_SAR8B_CV_0.XA6.CN1.n15 53.4593
R11992 SUNSAR_SAR8B_CV_0.XA6.CN1.n16 SUNSAR_SAR8B_CV_0.XA6.CN1.t4 38.8894
R11993 SUNSAR_SAR8B_CV_0.XA6.CN1.n16 SUNSAR_SAR8B_CV_0.XA6.CN1.t7 38.8894
R11994 SUNSAR_SAR8B_CV_0.XA6.CN1.n13 SUNSAR_SAR8B_CV_0.XA6.CN1.t1 38.8894
R11995 SUNSAR_SAR8B_CV_0.XA6.CN1.n13 SUNSAR_SAR8B_CV_0.XA6.CN1.t3 38.8894
R11996 SUNSAR_SAR8B_CV_0.XA6.CN1.n15 SUNSAR_SAR8B_CV_0.XA6.CN1.n14 38.024
R11997 SUNSAR_SAR8B_CV_0.XA6.CN1.n18 SUNSAR_SAR8B_CV_0.XA6.CN1.n17 38.024
R11998 SUNSAR_SAR8B_CV_0.XA6.CN1.n6 SUNSAR_SAR8B_CV_0.XA6.CN1.n3 20.3299
R11999 SUNSAR_SAR8B_CV_0.XA6.CN1.n3 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12000 SUNSAR_SAR8B_CV_0.XA6.CN1.n4 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12001 SUNSAR_SAR8B_CV_0.XA6.CN1.n5 SUNSAR_SAR8B_CV_0.XA6.CN1.n2 20.3299
R12002 SUNSAR_SAR8B_CV_0.XA6.CN1.n5 SUNSAR_SAR8B_CV_0.XA6.CN1.n4 20.3299
R12003 SUNSAR_SAR8B_CV_0.XA6.CN1.n5 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12004 SUNSAR_SAR8B_CV_0.XA6.CN1.n6 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12005 SUNSAR_SAR8B_CV_0.XA6.CN1.n8 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12006 SUNSAR_SAR8B_CV_0.XA6.CN1.n8 SUNSAR_SAR8B_CV_0.XA6.CN1.n7 20.3299
R12007 SUNSAR_SAR8B_CV_0.XA6.CN1.n7 SUNSAR_SAR8B_CV_0.XA6.CN1.n6 20.3299
R12008 SUNSAR_SAR8B_CV_0.XA6.CN1.n7 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12009 SUNSAR_SAR8B_CV_0.XA6.CN1.n2 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12010 SUNSAR_SAR8B_CV_0.XA6.CN1.n9 SUNSAR_SAR8B_CV_0.XA6.CN1.n2 20.3299
R12011 SUNSAR_SAR8B_CV_0.XA6.CN1.n14 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12012 SUNSAR_SAR8B_CV_0.XA6.CN1.n17 SUNSAR_SAR8B_CV_0.XA6.CN1 20.3299
R12013 SUNSAR_SAR8B_CV_0.XA6.CN1.n10 SUNSAR_SAR8B_CV_0.XA6.CN1 13.5534
R12014 SUNSAR_SAR8B_CV_0.XA6.CN1.n12 SUNSAR_SAR8B_CV_0.XA6.CN1.n9 12.8005
R12015 SUNSAR_SAR8B_CV_0.XA6.CN1.n12 SUNSAR_SAR8B_CV_0.XA6.CN1.n11 9.39466
R12016 SUNSAR_SAR8B_CV_0.XA6.CN1.n11 SUNSAR_SAR8B_CV_0.XA6.CN1.n10 9.39462
R12017 SUNSAR_SAR8B_CV_0.XA6.CN1.n10 SUNSAR_SAR8B_CV_0.XA6.CN1.n9 6.77697
R12018 SUNSAR_SAR8B_CV_0.XA6.CN1.n11 SUNSAR_SAR8B_CV_0.XA6.CN1 3.95537
R12019 SUNSAR_SAR8B_CV_0.D<1>.t8 SUNSAR_SAR8B_CV_0.D<1>.t11 1060.4
R12020 SUNSAR_SAR8B_CV_0.D<1>.t11 SUNSAR_SAR8B_CV_0.D<1> 589.284
R12021 SUNSAR_SAR8B_CV_0.D<1>.n10 SUNSAR_SAR8B_CV_0.D<1>.t8 573.85
R12022 SUNSAR_SAR8B_CV_0.D<1>.n5 SUNSAR_SAR8B_CV_0.D<1>.t10 568.956
R12023 SUNSAR_SAR8B_CV_0.D<1>.n4 SUNSAR_SAR8B_CV_0.D<1>.t9 568.956
R12024 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.D<1>.n0 312.829
R12025 SUNSAR_SAR8B_CV_0.D<1>.n7 SUNSAR_SAR8B_CV_0.D<1>.n3 297.865
R12026 SUNSAR_SAR8B_CV_0.D<1>.n2 SUNSAR_SAR8B_CV_0.D<1>.n1 92.5005
R12027 SUNSAR_SAR8B_CV_0.D<1>.n23 SUNSAR_SAR8B_CV_0.D<1>.n22 92.5005
R12028 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.D<1>.n24 90.7299
R12029 SUNSAR_SAR8B_CV_0.D<1>.n8 SUNSAR_SAR8B_CV_0.D<1> 81.6946
R12030 SUNSAR_SAR8B_CV_0.D<1>.n0 SUNSAR_SAR8B_CV_0.D<1>.t6 63.8431
R12031 SUNSAR_SAR8B_CV_0.D<1>.n0 SUNSAR_SAR8B_CV_0.D<1>.t5 63.8431
R12032 SUNSAR_SAR8B_CV_0.D<1>.n3 SUNSAR_SAR8B_CV_0.D<1>.t7 63.8431
R12033 SUNSAR_SAR8B_CV_0.D<1>.n3 SUNSAR_SAR8B_CV_0.D<1>.t4 63.8431
R12034 SUNSAR_SAR8B_CV_0.D<1>.n24 SUNSAR_SAR8B_CV_0.D<1>.n21 48.7856
R12035 SUNSAR_SAR8B_CV_0.D<1>.n1 SUNSAR_SAR8B_CV_0.D<1>.t1 38.8894
R12036 SUNSAR_SAR8B_CV_0.D<1>.n1 SUNSAR_SAR8B_CV_0.D<1>.t2 38.8894
R12037 SUNSAR_SAR8B_CV_0.D<1>.n22 SUNSAR_SAR8B_CV_0.D<1>.t3 38.8894
R12038 SUNSAR_SAR8B_CV_0.D<1>.n22 SUNSAR_SAR8B_CV_0.D<1>.t0 38.8894
R12039 SUNSAR_SAR8B_CV_0.D<1>.n24 SUNSAR_SAR8B_CV_0.D<1>.n23 38.024
R12040 SUNSAR_SAR8B_CV_0.D<1>.n16 SUNSAR_SAR8B_CV_0.D<1>.n15 31.7924
R12041 SUNSAR_SAR8B_CV_0.D<1>.n8 SUNSAR_SAR8B_CV_0.D<1>.n2 31.624
R12042 SUNSAR_SAR8B_CV_0.D<1>.n15 SUNSAR_SAR8B_CV_0.D<1> 22.6589
R12043 SUNSAR_SAR8B_CV_0.D<1>.n4 SUNSAR_SAR8B_CV_0.D<1> 20.3299
R12044 SUNSAR_SAR8B_CV_0.D<1>.n5 SUNSAR_SAR8B_CV_0.D<1>.n4 20.3299
R12045 SUNSAR_SAR8B_CV_0.D<1>.n2 SUNSAR_SAR8B_CV_0.D<1> 20.3299
R12046 SUNSAR_SAR8B_CV_0.D<1>.n23 SUNSAR_SAR8B_CV_0.D<1> 20.3299
R12047 SUNSAR_SAR8B_CV_0.D<1>.n19 SUNSAR_SAR8B_CV_0.D<1>.n8 17.9961
R12048 SUNSAR_SAR8B_CV_0.D<1>.n14 SUNSAR_SAR8B_CV_0.D<1>.n13 16.9417
R12049 SUNSAR_SAR8B_CV_0.D<1>.n7 SUNSAR_SAR8B_CV_0.D<1>.n6 13.7377
R12050 SUNSAR_SAR8B_CV_0.D<1>.n10 SUNSAR_SAR8B_CV_0.D<1> 12.939
R12051 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.D<1>.n7 10.6968
R12052 SUNSAR_SAR8B_CV_0.D<1>.n6 SUNSAR_SAR8B_CV_0.D<1> 10.633
R12053 SUNSAR_SAR8B_CV_0.D<1>.n12 SUNSAR_SAR8B_CV_0.D<1>.n10 10.4477
R12054 SUNSAR_SAR8B_CV_0.D<1>.n21 SUNSAR_SAR8B_CV_0.D<1>.n20 9.3005
R12055 SUNSAR_SAR8B_CV_0.D<1>.n21 SUNSAR_SAR8B_CV_0.D<1>.n8 8.11757
R12056 SUNSAR_SAR8B_CV_0.D<1>.n6 SUNSAR_SAR8B_CV_0.D<1>.n5 5.42812
R12057 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.D<1>.n16 4.9076
R12058 SUNSAR_SAR8B_CV_0.D<1>.n20 SUNSAR_SAR8B_CV_0.D<1>.n9 4.5005
R12059 SUNSAR_SAR8B_CV_0.D<1>.n19 SUNSAR_SAR8B_CV_0.D<1>.n18 4.5005
R12060 SUNSAR_SAR8B_CV_0.D<1>.n14 SUNSAR_SAR8B_CV_0.D<1>.n9 3.4105
R12061 SUNSAR_SAR8B_CV_0.D<1>.n18 SUNSAR_SAR8B_CV_0.D<1>.n17 3.4105
R12062 SUNSAR_SAR8B_CV_0.D<1>.n13 SUNSAR_SAR8B_CV_0.D<1> 0.329788
R12063 SUNSAR_SAR8B_CV_0.D<1>.n18 SUNSAR_SAR8B_CV_0.D<1>.n9 0.191676
R12064 SUNSAR_SAR8B_CV_0.D<1>.n20 SUNSAR_SAR8B_CV_0.D<1>.n19 0.191676
R12065 SUNSAR_SAR8B_CV_0.D<1>.n15 SUNSAR_SAR8B_CV_0.D<1> 0.168144
R12066 SUNSAR_SAR8B_CV_0.D<1>.n11 SUNSAR_SAR8B_CV_0.D<1> 0.132853
R12067 SUNSAR_SAR8B_CV_0.D<1>.n11 SUNSAR_SAR8B_CV_0.D<1> 0.108934
R12068 SUNSAR_SAR8B_CV_0.D<1>.n17 SUNSAR_SAR8B_CV_0.D<1>.n14 0.0723824
R12069 SUNSAR_SAR8B_CV_0.D<1>.n12 SUNSAR_SAR8B_CV_0.D<1>.n11 0.0547169
R12070 SUNSAR_SAR8B_CV_0.D<1>.n17 SUNSAR_SAR8B_CV_0.D<1> 0.0281471
R12071 SUNSAR_SAR8B_CV_0.D<1>.n16 SUNSAR_SAR8B_CV_0.D<1> 0.00726261
R12072 SUNSAR_SAR8B_CV_0.D<1>.n13 SUNSAR_SAR8B_CV_0.D<1>.n12 0.00351205
R12073 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t8 568.956
R12074 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t9 568.956
R12075 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n0 312.829
R12076 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n15 292.5
R12077 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n16 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 197.272
R12078 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n18 92.5005
R12079 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n22 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n21 92.5005
R12080 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n23 90.7299
R12081 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t4 63.8431
R12082 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t5 63.8431
R12083 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t6 63.8431
R12084 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n15 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t7 63.8431
R12085 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n17 59.1064
R12086 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n12 57.1591
R12087 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n23 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n20 53.4593
R12088 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t2 38.8894
R12089 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n18 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t0 38.8894
R12090 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n21 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t1 38.8894
R12091 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n21 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.t3 38.8894
R12092 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n20 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n19 38.024
R12093 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n23 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n22 38.024
R12094 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 31.624
R12095 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 20.3299
R12096 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n14 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n13 20.3299
R12097 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n14 20.3299
R12098 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n16 20.3299
R12099 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n19 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 20.3299
R12100 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n22 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 20.3299
R12101 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12102 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12103 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12104 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12105 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12106 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.325
R12107 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12108 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12109 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12110 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12111 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12112 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 12.323
R12113 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n17 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 10.3476
R12114 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n1 7.56982
R12115 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n3 7.56982
R12116 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n5 7.56982
R12117 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n7 7.56982
R12118 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n9 7.56982
R12119 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n11 7.56982
R12120 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n10 1.10785
R12121 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n8 1.10785
R12122 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n6 1.10785
R12123 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n4 1.10785
R12124 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n2 1.10785
R12125 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.168144
R12126 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t15 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t13 1060.4
R12127 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t9 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t8 1060.4
R12128 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t11 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t10 1060.4
R12129 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t12 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t14 1060.4
R12130 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t13 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n11 568.956
R12131 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t15 568.956
R12132 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t8 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n13 568.956
R12133 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t9 568.956
R12134 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t11 568.956
R12135 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t10 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n16 568.956
R12136 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t12 568.956
R12137 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t14 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n10 568.956
R12138 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n0 312.829
R12139 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n5 312.829
R12140 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n17 197.272
R12141 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n1 92.5005
R12142 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n8 92.5005
R12143 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 90.7299
R12144 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t7 63.8431
R12145 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n0 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t2 63.8431
R12146 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t0 63.8431
R12147 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n5 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t5 63.8431
R12148 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 61.177
R12149 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n3 53.4593
R12150 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t6 38.8894
R12151 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n8 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t4 38.8894
R12152 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t1 38.8894
R12153 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n1 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t3 38.8894
R12154 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n3 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n2 38.024
R12155 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n9 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n7 38.024
R12156 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n4 31.7584
R12157 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n7 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n6 29.5534
R12158 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 21.2766
R12159 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n2 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12160 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n11 20.3299
R12161 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n11 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12162 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n12 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12163 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n10 20.3299
R12164 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n12 20.3299
R12165 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n13 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12166 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n14 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12167 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12168 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n16 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n15 20.3299
R12169 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n14 20.3299
R12170 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n15 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12171 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n10 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12172 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n10 20.3299
R12173 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n17 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 20.3299
R12174 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n9 20.3299
R12175 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n6 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 10.3476
R12176 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n4 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.168144
R12177 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t9 568.956
R12178 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t8 568.956
R12179 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n0 312.829
R12180 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n5 292.5
R12181 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 197.272
R12182 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n8 92.5005
R12183 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n11 92.5005
R12184 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n13 90.7299
R12185 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t4 63.8431
R12186 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t7 63.8431
R12187 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t5 63.8431
R12188 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t6 63.8431
R12189 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n7 59.1064
R12190 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n10 53.4593
R12191 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t0 38.8894
R12192 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t1 38.8894
R12193 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t2 38.8894
R12194 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.t3 38.8894
R12195 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n9 38.024
R12196 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n12 38.024
R12197 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n2 36.6593
R12198 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 31.624
R12199 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 20.3299
R12200 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n3 20.3299
R12201 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n4 20.3299
R12202 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n6 20.3299
R12203 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 20.3299
R12204 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 20.3299
R12205 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 12.325
R12206 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 12.323
R12207 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 10.3476
R12208 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n1 8.95217
R12209 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.168144
R12210 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t7 1060.4
R12211 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t5 1060.4
R12212 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t8 1060.4
R12213 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t4 1060.4
R12214 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n1 568.956
R12215 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t3 568.956
R12216 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n3 568.956
R12217 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t6 568.956
R12218 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t2 568.956
R12219 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n6 568.956
R12220 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t9 568.956
R12221 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n0 568.956
R12222 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t0 356.344
R12223 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.t1 135.293
R12224 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n10 128.754
R12225 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n1 20.3299
R12226 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA1.XA4.MP3.G 20.3299
R12227 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA1.XA4.MN3.G 20.3299
R12228 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n0 20.3299
R12229 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n2 20.3299
R12230 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA1.XA4.MN2.G 20.3299
R12231 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA1.XA4.MP2.G 20.3299
R12232 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA1.XA4.MP0.G 20.3299
R12233 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n5 20.3299
R12234 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n4 20.3299
R12235 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA1.XA4.MP1.G 20.3299
R12236 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA1.XA4.MN1.G 20.3299
R12237 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n0 20.3299
R12238 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.D 20.3299
R12239 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n8 16.3643
R12240 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n9 15.2303
R12241 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA1.XA4.MN0.G 15.1965
R12242 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n7 3.93805
R12243 SUNSAR_SAR8B_CV_0.XA6.CP0.t14 SUNSAR_SAR8B_CV_0.XA6.CP0.t8 1060.4
R12244 SUNSAR_SAR8B_CV_0.XA6.CP0.t15 SUNSAR_SAR8B_CV_0.XA6.CP0.t12 1060.4
R12245 SUNSAR_SAR8B_CV_0.XA6.CP0.t13 SUNSAR_SAR8B_CV_0.XA6.CP0.t11 1060.4
R12246 SUNSAR_SAR8B_CV_0.XA6.CP0.t9 SUNSAR_SAR8B_CV_0.XA6.CP0.t10 1060.4
R12247 SUNSAR_SAR8B_CV_0.XA6.CP0.t8 SUNSAR_SAR8B_CV_0.XA6.CP0.n4 568.956
R12248 SUNSAR_SAR8B_CV_0.XA6.CP0.n5 SUNSAR_SAR8B_CV_0.XA6.CP0.t14 568.956
R12249 SUNSAR_SAR8B_CV_0.XA6.CP0.t12 SUNSAR_SAR8B_CV_0.XA6.CP0.n6 568.956
R12250 SUNSAR_SAR8B_CV_0.XA6.CP0.n7 SUNSAR_SAR8B_CV_0.XA6.CP0.t15 568.956
R12251 SUNSAR_SAR8B_CV_0.XA6.CP0.n10 SUNSAR_SAR8B_CV_0.XA6.CP0.t13 568.956
R12252 SUNSAR_SAR8B_CV_0.XA6.CP0.t11 SUNSAR_SAR8B_CV_0.XA6.CP0.n9 568.956
R12253 SUNSAR_SAR8B_CV_0.XA6.CP0.n8 SUNSAR_SAR8B_CV_0.XA6.CP0.t9 568.956
R12254 SUNSAR_SAR8B_CV_0.XA6.CP0.t10 SUNSAR_SAR8B_CV_0.XA6.CP0.n3 568.956
R12255 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.CP0.n1 312.829
R12256 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.CP0.n0 312.829
R12257 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.CP0.n10 197.272
R12258 SUNSAR_SAR8B_CV_0.XA6.CP0.n12 SUNSAR_SAR8B_CV_0.XA6.CP0.n11 92.5005
R12259 SUNSAR_SAR8B_CV_0.XA6.CP0.n15 SUNSAR_SAR8B_CV_0.XA6.CP0.n14 92.5005
R12260 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.CP0.n16 90.7299
R12261 SUNSAR_SAR8B_CV_0.XA6.CP0.n0 SUNSAR_SAR8B_CV_0.XA6.CP0.t1 63.8431
R12262 SUNSAR_SAR8B_CV_0.XA6.CP0.n0 SUNSAR_SAR8B_CV_0.XA6.CP0.t3 63.8431
R12263 SUNSAR_SAR8B_CV_0.XA6.CP0.n1 SUNSAR_SAR8B_CV_0.XA6.CP0.t2 63.8431
R12264 SUNSAR_SAR8B_CV_0.XA6.CP0.n1 SUNSAR_SAR8B_CV_0.XA6.CP0.t4 63.8431
R12265 SUNSAR_SAR8B_CV_0.XA6.CP0.n2 SUNSAR_SAR8B_CV_0.XA6.CP0 61.177
R12266 SUNSAR_SAR8B_CV_0.XA6.CP0.n16 SUNSAR_SAR8B_CV_0.XA6.CP0.n13 53.4593
R12267 SUNSAR_SAR8B_CV_0.XA6.CP0.n11 SUNSAR_SAR8B_CV_0.XA6.CP0.t5 38.8894
R12268 SUNSAR_SAR8B_CV_0.XA6.CP0.n11 SUNSAR_SAR8B_CV_0.XA6.CP0.t6 38.8894
R12269 SUNSAR_SAR8B_CV_0.XA6.CP0.n14 SUNSAR_SAR8B_CV_0.XA6.CP0.t0 38.8894
R12270 SUNSAR_SAR8B_CV_0.XA6.CP0.n14 SUNSAR_SAR8B_CV_0.XA6.CP0.t7 38.8894
R12271 SUNSAR_SAR8B_CV_0.XA6.CP0.n13 SUNSAR_SAR8B_CV_0.XA6.CP0.n12 38.024
R12272 SUNSAR_SAR8B_CV_0.XA6.CP0.n16 SUNSAR_SAR8B_CV_0.XA6.CP0.n15 38.024
R12273 SUNSAR_SAR8B_CV_0.XA6.CP0.n13 SUNSAR_SAR8B_CV_0.XA6.CP0.n2 29.5534
R12274 SUNSAR_SAR8B_CV_0.XA6.CP0.n7 SUNSAR_SAR8B_CV_0.XA6.CP0.n4 20.3299
R12275 SUNSAR_SAR8B_CV_0.XA6.CP0.n4 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12276 SUNSAR_SAR8B_CV_0.XA6.CP0.n5 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12277 SUNSAR_SAR8B_CV_0.XA6.CP0.n6 SUNSAR_SAR8B_CV_0.XA6.CP0.n3 20.3299
R12278 SUNSAR_SAR8B_CV_0.XA6.CP0.n6 SUNSAR_SAR8B_CV_0.XA6.CP0.n5 20.3299
R12279 SUNSAR_SAR8B_CV_0.XA6.CP0.n6 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12280 SUNSAR_SAR8B_CV_0.XA6.CP0.n7 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12281 SUNSAR_SAR8B_CV_0.XA6.CP0.n9 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12282 SUNSAR_SAR8B_CV_0.XA6.CP0.n9 SUNSAR_SAR8B_CV_0.XA6.CP0.n8 20.3299
R12283 SUNSAR_SAR8B_CV_0.XA6.CP0.n8 SUNSAR_SAR8B_CV_0.XA6.CP0.n7 20.3299
R12284 SUNSAR_SAR8B_CV_0.XA6.CP0.n8 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12285 SUNSAR_SAR8B_CV_0.XA6.CP0.n3 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12286 SUNSAR_SAR8B_CV_0.XA6.CP0.n10 SUNSAR_SAR8B_CV_0.XA6.CP0.n3 20.3299
R12287 SUNSAR_SAR8B_CV_0.XA6.CP0.n10 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12288 SUNSAR_SAR8B_CV_0.XA6.CP0.n12 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12289 SUNSAR_SAR8B_CV_0.XA6.CP0.n15 SUNSAR_SAR8B_CV_0.XA6.CP0 20.3299
R12290 SUNSAR_SAR8B_CV_0.XA6.CP0.n2 SUNSAR_SAR8B_CV_0.XA6.CP0 10.3476
R12291 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t9 568.956
R12292 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t8 568.956
R12293 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n0 312.829
R12294 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n5 292.5
R12295 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 197.272
R12296 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n8 92.5005
R12297 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n11 92.5005
R12298 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n13 90.7299
R12299 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t5 63.8431
R12300 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t7 63.8431
R12301 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t6 63.8431
R12302 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t4 63.8431
R12303 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n7 59.1064
R12304 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n10 53.4593
R12305 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n2 39.4245
R12306 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t2 38.8894
R12307 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t1 38.8894
R12308 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t3 38.8894
R12309 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.t0 38.8894
R12310 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n9 38.024
R12311 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n12 38.024
R12312 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 31.624
R12313 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 20.3299
R12314 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n3 20.3299
R12315 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n4 20.3299
R12316 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n6 20.3299
R12317 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 20.3299
R12318 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 20.3299
R12319 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 12.325
R12320 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 12.323
R12321 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 10.3476
R12322 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n1 10.3345
R12323 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.168144
R12324 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t5 1060.4
R12325 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t8 1060.4
R12326 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t7 1060.4
R12327 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t4 1060.4
R12328 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n2 568.956
R12329 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t6 568.956
R12330 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n4 568.956
R12331 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t9 568.956
R12332 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t3 568.956
R12333 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n7 568.956
R12334 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t2 568.956
R12335 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n1 568.956
R12336 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t0 356.344
R12337 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.D SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.t1 151.719
R12338 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.D 128.754
R12339 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n8 97.8829
R12340 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n2 20.3299
R12341 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA5.XA2.MN3.G 20.3299
R12342 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA5.XA2.MP3.G 20.3299
R12343 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n1 20.3299
R12344 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n3 20.3299
R12345 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA5.XA2.MP2.G 20.3299
R12346 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA5.XA2.MN2.G 20.3299
R12347 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA5.XA2.MN0.G 20.3299
R12348 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n6 20.3299
R12349 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n5 20.3299
R12350 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA5.XA2.MN1.G 20.3299
R12351 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA5.XA2.MP1.G 20.3299
R12352 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n1 20.3299
R12353 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA5.XA2.MP0.G 20.3299
R12354 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n0 20.3299
R12355 SUNSAR_SAR8B_CV_0.XA5.CN1.t11 SUNSAR_SAR8B_CV_0.XA5.CN1.t12 1060.4
R12356 SUNSAR_SAR8B_CV_0.XA5.CN1.t8 SUNSAR_SAR8B_CV_0.XA5.CN1.t15 1060.4
R12357 SUNSAR_SAR8B_CV_0.XA5.CN1.t13 SUNSAR_SAR8B_CV_0.XA5.CN1.t10 1060.4
R12358 SUNSAR_SAR8B_CV_0.XA5.CN1.t14 SUNSAR_SAR8B_CV_0.XA5.CN1.t9 1060.4
R12359 SUNSAR_SAR8B_CV_0.XA5.CN1.t12 SUNSAR_SAR8B_CV_0.XA5.CN1.n1 568.956
R12360 SUNSAR_SAR8B_CV_0.XA5.CN1.n2 SUNSAR_SAR8B_CV_0.XA5.CN1.t11 568.956
R12361 SUNSAR_SAR8B_CV_0.XA5.CN1.t15 SUNSAR_SAR8B_CV_0.XA5.CN1.n3 568.956
R12362 SUNSAR_SAR8B_CV_0.XA5.CN1.n4 SUNSAR_SAR8B_CV_0.XA5.CN1.t8 568.956
R12363 SUNSAR_SAR8B_CV_0.XA5.CN1.n7 SUNSAR_SAR8B_CV_0.XA5.CN1.t13 568.956
R12364 SUNSAR_SAR8B_CV_0.XA5.CN1.t10 SUNSAR_SAR8B_CV_0.XA5.CN1.n6 568.956
R12365 SUNSAR_SAR8B_CV_0.XA5.CN1.n5 SUNSAR_SAR8B_CV_0.XA5.CN1.t14 568.956
R12366 SUNSAR_SAR8B_CV_0.XA5.CN1.t9 SUNSAR_SAR8B_CV_0.XA5.CN1.n0 568.956
R12367 SUNSAR_SAR8B_CV_0.XA5.CN1.n12 SUNSAR_SAR8B_CV_0.XA5.CN1.n11 292.5
R12368 SUNSAR_SAR8B_CV_0.XA5.CN1.n17 SUNSAR_SAR8B_CV_0.XA5.CN1.n16 292.5
R12369 SUNSAR_SAR8B_CV_0.XA5.CN1.n10 SUNSAR_SAR8B_CV_0.XA5.CN1 197.272
R12370 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.CN1.n14 112.829
R12371 SUNSAR_SAR8B_CV_0.XA5.CN1.n13 SUNSAR_SAR8B_CV_0.XA5.CN1.n12 111.059
R12372 SUNSAR_SAR8B_CV_0.XA5.CN1.n17 SUNSAR_SAR8B_CV_0.XA5.CN1.n15 111.059
R12373 SUNSAR_SAR8B_CV_0.XA5.CN1.n10 SUNSAR_SAR8B_CV_0.XA5.CN1.n9 92.5005
R12374 SUNSAR_SAR8B_CV_0.XA5.CN1.n16 SUNSAR_SAR8B_CV_0.XA5.CN1.t7 63.8431
R12375 SUNSAR_SAR8B_CV_0.XA5.CN1.n16 SUNSAR_SAR8B_CV_0.XA5.CN1.t5 63.8431
R12376 SUNSAR_SAR8B_CV_0.XA5.CN1.n11 SUNSAR_SAR8B_CV_0.XA5.CN1.t6 63.8431
R12377 SUNSAR_SAR8B_CV_0.XA5.CN1.n11 SUNSAR_SAR8B_CV_0.XA5.CN1.t4 63.8431
R12378 SUNSAR_SAR8B_CV_0.XA5.CN1.n15 SUNSAR_SAR8B_CV_0.XA5.CN1.n13 53.4593
R12379 SUNSAR_SAR8B_CV_0.XA5.CN1.n9 SUNSAR_SAR8B_CV_0.XA5.CN1.t1 38.8894
R12380 SUNSAR_SAR8B_CV_0.XA5.CN1.n9 SUNSAR_SAR8B_CV_0.XA5.CN1.t2 38.8894
R12381 SUNSAR_SAR8B_CV_0.XA5.CN1.n14 SUNSAR_SAR8B_CV_0.XA5.CN1.t0 38.8894
R12382 SUNSAR_SAR8B_CV_0.XA5.CN1.n14 SUNSAR_SAR8B_CV_0.XA5.CN1.t3 38.8894
R12383 SUNSAR_SAR8B_CV_0.XA5.CN1.n4 SUNSAR_SAR8B_CV_0.XA5.CN1.n1 20.3299
R12384 SUNSAR_SAR8B_CV_0.XA5.CN1.n1 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12385 SUNSAR_SAR8B_CV_0.XA5.CN1.n2 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12386 SUNSAR_SAR8B_CV_0.XA5.CN1.n3 SUNSAR_SAR8B_CV_0.XA5.CN1.n0 20.3299
R12387 SUNSAR_SAR8B_CV_0.XA5.CN1.n3 SUNSAR_SAR8B_CV_0.XA5.CN1.n2 20.3299
R12388 SUNSAR_SAR8B_CV_0.XA5.CN1.n3 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12389 SUNSAR_SAR8B_CV_0.XA5.CN1.n4 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12390 SUNSAR_SAR8B_CV_0.XA5.CN1.n6 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12391 SUNSAR_SAR8B_CV_0.XA5.CN1.n6 SUNSAR_SAR8B_CV_0.XA5.CN1.n5 20.3299
R12392 SUNSAR_SAR8B_CV_0.XA5.CN1.n5 SUNSAR_SAR8B_CV_0.XA5.CN1.n4 20.3299
R12393 SUNSAR_SAR8B_CV_0.XA5.CN1.n5 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12394 SUNSAR_SAR8B_CV_0.XA5.CN1.n0 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12395 SUNSAR_SAR8B_CV_0.XA5.CN1.n7 SUNSAR_SAR8B_CV_0.XA5.CN1.n0 20.3299
R12396 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.CN1.n10 20.3299
R12397 SUNSAR_SAR8B_CV_0.XA5.CN1.n12 SUNSAR_SAR8B_CV_0.XA5.CN1 20.3299
R12398 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.CN1.n17 20.3299
R12399 SUNSAR_SAR8B_CV_0.XA5.CN1.n13 SUNSAR_SAR8B_CV_0.XA5.CN1 17.6946
R12400 SUNSAR_SAR8B_CV_0.XA5.CN1.n15 SUNSAR_SAR8B_CV_0.XA5.CN1 17.6946
R12401 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.CN1.n8 10.6647
R12402 SUNSAR_SAR8B_CV_0.XA5.CN1.n8 SUNSAR_SAR8B_CV_0.XA5.CN1 7.91546
R12403 SUNSAR_SAR8B_CV_0.XA5.CN1.n8 SUNSAR_SAR8B_CV_0.XA5.CN1.n7 5.39616
R12404 SUNSAR_SAR8B_CV_0.DONE.t14 SUNSAR_SAR8B_CV_0.DONE.t7 1060.4
R12405 SUNSAR_SAR8B_CV_0.DONE.t6 SUNSAR_SAR8B_CV_0.DONE.t11 1060.4
R12406 SUNSAR_SAR8B_CV_0.DONE.t9 SUNSAR_SAR8B_CV_0.DONE.t5 1060.4
R12407 SUNSAR_SAR8B_CV_0.DONE.t21 SUNSAR_SAR8B_CV_0.DONE.t12 1060.4
R12408 SUNSAR_SAR8B_CV_0.DONE.t3 SUNSAR_SAR8B_CV_0.DONE.t4 1060.4
R12409 SUNSAR_SAR8B_CV_0.DONE.t15 SUNSAR_SAR8B_CV_0.DONE.t16 1060.4
R12410 SUNSAR_SAR8B_CV_0.DONE.t13 SUNSAR_SAR8B_CV_0.DONE.t17 1060.4
R12411 SUNSAR_SAR8B_CV_0.DONE.t19 SUNSAR_SAR8B_CV_0.DONE.t8 1060.4
R12412 SUNSAR_SAR8B_CV_0.DONE.t2 SUNSAR_SAR8B_CV_0.DONE.t20 1060.4
R12413 SUNSAR_SAR8B_CV_0.DONE.t18 SUNSAR_SAR8B_CV_0.DONE.t10 1060.4
R12414 SUNSAR_SAR8B_CV_0.DONE.n19 SUNSAR_SAR8B_CV_0.DONE.n17 776.083
R12415 SUNSAR_SAR8B_CV_0.DONE.n15 SUNSAR_SAR8B_CV_0.DONE.n13 776.083
R12416 SUNSAR_SAR8B_CV_0.DONE.n11 SUNSAR_SAR8B_CV_0.DONE.n9 776.083
R12417 SUNSAR_SAR8B_CV_0.DONE.n7 SUNSAR_SAR8B_CV_0.DONE.n5 776.083
R12418 SUNSAR_SAR8B_CV_0.DONE.n20 tt_um_TT06_SAR_done_0.DONE 774.226
R12419 SUNSAR_SAR8B_CV_0.DONE.t11 tt_um_TT06_SAR_done_0.x3.MP0.G 591.995
R12420 SUNSAR_SAR8B_CV_0.DONE.t7 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.G 589.284
R12421 SUNSAR_SAR8B_CV_0.DONE.t5 SUNSAR_CAPT8B_CV_0.XI14.XA1.MP0.G 589.284
R12422 SUNSAR_SAR8B_CV_0.DONE.t12 SUNSAR_CAPT8B_CV_0.XH13.XA1.MP0.G 589.284
R12423 SUNSAR_SAR8B_CV_0.DONE.t4 SUNSAR_CAPT8B_CV_0.XG12.XA1.MP0.G 589.284
R12424 SUNSAR_SAR8B_CV_0.DONE.t16 SUNSAR_CAPT8B_CV_0.XF11.XA1.MP0.G 589.284
R12425 SUNSAR_SAR8B_CV_0.DONE.t17 SUNSAR_CAPT8B_CV_0.XE10.XA1.MP0.G 589.284
R12426 SUNSAR_SAR8B_CV_0.DONE.t8 SUNSAR_CAPT8B_CV_0.XD09.XA1.MP0.G 589.284
R12427 SUNSAR_SAR8B_CV_0.DONE.t20 SUNSAR_CAPT8B_CV_0.XC08.XA1.MP0.G 589.284
R12428 SUNSAR_SAR8B_CV_0.DONE.t10 SUNSAR_CAPT8B_CV_0.XB07.XA1.MP0.G 589.284
R12429 SUNSAR_SAR8B_CV_0.DONE.n0 SUNSAR_SAR8B_CV_0.DONE.t14 574.351
R12430 SUNSAR_SAR8B_CV_0.DONE.n18 SUNSAR_SAR8B_CV_0.DONE.t9 573.85
R12431 SUNSAR_SAR8B_CV_0.DONE.n16 SUNSAR_SAR8B_CV_0.DONE.t21 573.85
R12432 SUNSAR_SAR8B_CV_0.DONE.n14 SUNSAR_SAR8B_CV_0.DONE.t3 573.85
R12433 SUNSAR_SAR8B_CV_0.DONE.n12 SUNSAR_SAR8B_CV_0.DONE.t15 573.85
R12434 SUNSAR_SAR8B_CV_0.DONE.n10 SUNSAR_SAR8B_CV_0.DONE.t13 573.85
R12435 SUNSAR_SAR8B_CV_0.DONE.n8 SUNSAR_SAR8B_CV_0.DONE.t19 573.85
R12436 SUNSAR_SAR8B_CV_0.DONE.n6 SUNSAR_SAR8B_CV_0.DONE.t2 573.85
R12437 SUNSAR_SAR8B_CV_0.DONE.n4 SUNSAR_SAR8B_CV_0.DONE.t18 573.85
R12438 SUNSAR_SAR8B_CV_0.DONE.n2 SUNSAR_SAR8B_CV_0.DONE.t6 568.956
R12439 SUNSAR_SAR8B_CV_0.DONE.n23 SUNSAR_SAR8B_CV_0.DONE.t1 356.344
R12440 SUNSAR_SAR8B_CV_0.DONE.n17 SUNSAR_SAR8B_CV_0.DONE.n15 152.649
R12441 SUNSAR_SAR8B_CV_0.DONE.n13 SUNSAR_SAR8B_CV_0.DONE.n11 152.649
R12442 SUNSAR_SAR8B_CV_0.DONE.n9 SUNSAR_SAR8B_CV_0.DONE.n7 152.649
R12443 SUNSAR_SAR8B_CV_0.DONE.n22 SUNSAR_SAR8B_CV_0.DONE.t0 136.785
R12444 SUNSAR_SAR8B_CV_0.XA7.XA8.MN0.D SUNSAR_SAR8B_CV_0.DONE.n23 128.754
R12445 SUNSAR_SAR8B_CV_0.DONE.n5 SUNSAR_CAPT8B_CV_0.DONE 76.3244
R12446 SUNSAR_SAR8B_CV_0.DONE.n20 SUNSAR_SAR8B_CV_0.DONE.n19 63.9008
R12447 SUNSAR_SAR8B_CV_0.DONE.n21 SUNSAR_SAR8B_CV_0.DONE.n20 24.0308
R12448 SUNSAR_SAR8B_CV_0.DONE.n23 SUNSAR_SAR8B_CV_0.XA7.XA8.MP0.D 20.3299
R12449 SUNSAR_SAR8B_CV_0.DONE.n2 SUNSAR_SAR8B_CV_0.DONE.n1 14.3064
R12450 SUNSAR_SAR8B_CV_0.DONE.n18 SUNSAR_CAPT8B_CV_0.XI14.XA1.MN0.G 12.9392
R12451 SUNSAR_SAR8B_CV_0.DONE.n16 SUNSAR_CAPT8B_CV_0.XH13.XA1.MN0.G 12.9392
R12452 SUNSAR_SAR8B_CV_0.DONE.n14 SUNSAR_CAPT8B_CV_0.XG12.XA1.MN0.G 12.9392
R12453 SUNSAR_SAR8B_CV_0.DONE.n12 SUNSAR_CAPT8B_CV_0.XF11.XA1.MN0.G 12.9392
R12454 SUNSAR_SAR8B_CV_0.DONE.n10 SUNSAR_CAPT8B_CV_0.XE10.XA1.MN0.G 12.9392
R12455 SUNSAR_SAR8B_CV_0.DONE.n8 SUNSAR_CAPT8B_CV_0.XD09.XA1.MN0.G 12.9392
R12456 SUNSAR_SAR8B_CV_0.DONE.n6 SUNSAR_CAPT8B_CV_0.XC08.XA1.MN0.G 12.9392
R12457 SUNSAR_SAR8B_CV_0.DONE.n4 SUNSAR_CAPT8B_CV_0.XB07.XA1.MN0.G 12.9392
R12458 SUNSAR_SAR8B_CV_0.XA7.XA8.MN0.D SUNSAR_SAR8B_CV_0.DONE.n22 10.6653
R12459 SUNSAR_SAR8B_CV_0.DONE.n0 SUNSAR_SAR8B_CV_0.XA20.XA11.MN1.G 10.664
R12460 SUNSAR_SAR8B_CV_0.DONE.n22 SUNSAR_SAR8B_CV_0.DONE.n21 8.71144
R12461 SUNSAR_SAR8B_CV_0.DONE.n3 SUNSAR_SAR8B_CV_0.DONE.n2 8.39597
R12462 SUNSAR_SAR8B_CV_0.DONE.n19 SUNSAR_SAR8B_CV_0.DONE.n18 8.17291
R12463 SUNSAR_SAR8B_CV_0.DONE.n17 SUNSAR_SAR8B_CV_0.DONE.n16 8.17291
R12464 SUNSAR_SAR8B_CV_0.DONE.n15 SUNSAR_SAR8B_CV_0.DONE.n14 8.17291
R12465 SUNSAR_SAR8B_CV_0.DONE.n13 SUNSAR_SAR8B_CV_0.DONE.n12 8.17291
R12466 SUNSAR_SAR8B_CV_0.DONE.n11 SUNSAR_SAR8B_CV_0.DONE.n10 8.17291
R12467 SUNSAR_SAR8B_CV_0.DONE.n9 SUNSAR_SAR8B_CV_0.DONE.n8 8.17291
R12468 SUNSAR_SAR8B_CV_0.DONE.n7 SUNSAR_SAR8B_CV_0.DONE.n6 8.17291
R12469 SUNSAR_SAR8B_CV_0.DONE.n5 SUNSAR_SAR8B_CV_0.DONE.n4 8.17291
R12470 SUNSAR_SAR8B_CV_0.DONE.n1 tt_um_TT06_SAR_done_0.x3.MN0.G 6.82717
R12471 SUNSAR_SAR8B_CV_0.DONE.n21 SUNSAR_SAR8B_CV_0.DONE.n0 6.58575
R12472 SUNSAR_SAR8B_CV_0.DONE.n1 tt_um_TT06_SAR_done_0.x3.MN0.G 6.02403
R12473 SUNSAR_SAR8B_CV_0.DONE.n3 tt_um_TT06_SAR_done_0.DONE 0.177583
R12474 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.DONE.n3 0.138487
R12475 SUNSAR_SAR8B_CV_0.XA7.CP0.t13 SUNSAR_SAR8B_CV_0.XA7.CP0.t14 1060.4
R12476 SUNSAR_SAR8B_CV_0.XA7.CP0.t9 SUNSAR_SAR8B_CV_0.XA7.CP0.t11 1060.4
R12477 SUNSAR_SAR8B_CV_0.XA7.CP0.t15 SUNSAR_SAR8B_CV_0.XA7.CP0.t12 1060.4
R12478 SUNSAR_SAR8B_CV_0.XA7.CP0.t10 SUNSAR_SAR8B_CV_0.XA7.CP0.t8 1060.4
R12479 SUNSAR_SAR8B_CV_0.XA7.CP0.t14 SUNSAR_SAR8B_CV_0.XA7.CP0.n1 568.956
R12480 SUNSAR_SAR8B_CV_0.XA7.CP0.n2 SUNSAR_SAR8B_CV_0.XA7.CP0.t13 568.956
R12481 SUNSAR_SAR8B_CV_0.XA7.CP0.t11 SUNSAR_SAR8B_CV_0.XA7.CP0.n3 568.956
R12482 SUNSAR_SAR8B_CV_0.XA7.CP0.n4 SUNSAR_SAR8B_CV_0.XA7.CP0.t9 568.956
R12483 SUNSAR_SAR8B_CV_0.XA7.CP0.n7 SUNSAR_SAR8B_CV_0.XA7.CP0.t15 568.956
R12484 SUNSAR_SAR8B_CV_0.XA7.CP0.t12 SUNSAR_SAR8B_CV_0.XA7.CP0.n6 568.956
R12485 SUNSAR_SAR8B_CV_0.XA7.CP0.n5 SUNSAR_SAR8B_CV_0.XA7.CP0.t10 568.956
R12486 SUNSAR_SAR8B_CV_0.XA7.CP0.t8 SUNSAR_SAR8B_CV_0.XA7.CP0.n0 568.956
R12487 SUNSAR_SAR8B_CV_0.XA7.CP0.n12 SUNSAR_SAR8B_CV_0.XA7.CP0.n11 292.5
R12488 SUNSAR_SAR8B_CV_0.XA7.CP0.n15 SUNSAR_SAR8B_CV_0.XA7.CP0.n14 292.5
R12489 SUNSAR_SAR8B_CV_0.XA7.CP0.n9 SUNSAR_SAR8B_CV_0.XA7.CP0 197.272
R12490 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CP0.n10 112.829
R12491 SUNSAR_SAR8B_CV_0.XA7.CP0.n13 SUNSAR_SAR8B_CV_0.XA7.CP0.n12 111.059
R12492 SUNSAR_SAR8B_CV_0.XA7.CP0.n9 SUNSAR_SAR8B_CV_0.XA7.CP0.n8 92.5005
R12493 SUNSAR_SAR8B_CV_0.XA7.CP0.n16 SUNSAR_SAR8B_CV_0.XA7.CP0.n15 81.5064
R12494 SUNSAR_SAR8B_CV_0.XA7.CP0.n14 SUNSAR_SAR8B_CV_0.XA7.CP0.t2 63.8431
R12495 SUNSAR_SAR8B_CV_0.XA7.CP0.n14 SUNSAR_SAR8B_CV_0.XA7.CP0.t1 63.8431
R12496 SUNSAR_SAR8B_CV_0.XA7.CP0.n11 SUNSAR_SAR8B_CV_0.XA7.CP0.t4 63.8431
R12497 SUNSAR_SAR8B_CV_0.XA7.CP0.n11 SUNSAR_SAR8B_CV_0.XA7.CP0.t6 63.8431
R12498 SUNSAR_SAR8B_CV_0.XA7.CP0.n17 SUNSAR_SAR8B_CV_0.XA7.CP0.n13 53.4593
R12499 SUNSAR_SAR8B_CV_0.XA7.CP0.n10 SUNSAR_SAR8B_CV_0.XA7.CP0.t3 38.8894
R12500 SUNSAR_SAR8B_CV_0.XA7.CP0.n10 SUNSAR_SAR8B_CV_0.XA7.CP0.t7 38.8894
R12501 SUNSAR_SAR8B_CV_0.XA7.CP0.n8 SUNSAR_SAR8B_CV_0.XA7.CP0.t0 38.8894
R12502 SUNSAR_SAR8B_CV_0.XA7.CP0.n8 SUNSAR_SAR8B_CV_0.XA7.CP0.t5 38.8894
R12503 SUNSAR_SAR8B_CV_0.XA7.CP0.n17 SUNSAR_SAR8B_CV_0.XA7.CP0.n16 29.5534
R12504 SUNSAR_SAR8B_CV_0.XA7.CP0.n4 SUNSAR_SAR8B_CV_0.XA7.CP0.n1 20.3299
R12505 SUNSAR_SAR8B_CV_0.XA7.CP0.n1 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12506 SUNSAR_SAR8B_CV_0.XA7.CP0.n2 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12507 SUNSAR_SAR8B_CV_0.XA7.CP0.n3 SUNSAR_SAR8B_CV_0.XA7.CP0.n0 20.3299
R12508 SUNSAR_SAR8B_CV_0.XA7.CP0.n3 SUNSAR_SAR8B_CV_0.XA7.CP0.n2 20.3299
R12509 SUNSAR_SAR8B_CV_0.XA7.CP0.n3 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12510 SUNSAR_SAR8B_CV_0.XA7.CP0.n4 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12511 SUNSAR_SAR8B_CV_0.XA7.CP0.n6 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12512 SUNSAR_SAR8B_CV_0.XA7.CP0.n6 SUNSAR_SAR8B_CV_0.XA7.CP0.n5 20.3299
R12513 SUNSAR_SAR8B_CV_0.XA7.CP0.n5 SUNSAR_SAR8B_CV_0.XA7.CP0.n4 20.3299
R12514 SUNSAR_SAR8B_CV_0.XA7.CP0.n5 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12515 SUNSAR_SAR8B_CV_0.XA7.CP0.n0 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12516 SUNSAR_SAR8B_CV_0.XA7.CP0.n7 SUNSAR_SAR8B_CV_0.XA7.CP0.n0 20.3299
R12517 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CP0.n7 20.3299
R12518 SUNSAR_SAR8B_CV_0.XA7.CP0.n12 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12519 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CP0.n9 20.3299
R12520 SUNSAR_SAR8B_CV_0.XA7.CP0.n15 SUNSAR_SAR8B_CV_0.XA7.CP0 20.3299
R12521 SUNSAR_SAR8B_CV_0.XA7.CP0.n13 SUNSAR_SAR8B_CV_0.XA7.CP0 17.6946
R12522 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CP0.n17 17.6946
R12523 SUNSAR_SAR8B_CV_0.XA7.CP0.n16 SUNSAR_SAR8B_CV_0.XA7.CP0 10.3476
R12524 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n5 8084.31
R12525 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n4 2095.71
R12526 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t4 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t3 1060.4
R12527 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t2 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t5 1060.4
R12528 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n4 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n2 705.585
R12529 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t3 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 589.284
R12530 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t5 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 589.284
R12531 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n3 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t4 573.85
R12532 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n2 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t2 573.85
R12533 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t1 376.673
R12534 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n0 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.t0 131.389
R12535 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n1 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 121.977
R12536 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n3 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 12.9392
R12537 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n2 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 12.9392
R12538 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n5 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 12.8005
R12539 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n7 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n0 12.8005
R12540 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n4 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n3 10.82
R12541 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n7 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n6 9.39659
R12542 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n6 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n1 9.39269
R12543 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n7 7.52991
R12544 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n1 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n0 6.77697
R12545 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n5 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 6.4005
R12546 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n6 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 4.83062
R12547 SUNSAR_SAR8B_CV_0.XB1.CKN.t7 SUNSAR_SAR8B_CV_0.XB1.CKN.t5 1060.4
R12548 SUNSAR_SAR8B_CV_0.XB1.CKN.t6 SUNSAR_SAR8B_CV_0.XB1.CKN.t2 1060.4
R12549 SUNSAR_SAR8B_CV_0.XB1.CKN.t5 SUNSAR_SAR8B_CV_0.XB1.XA4.MP0.G 589.284
R12550 SUNSAR_SAR8B_CV_0.XB1.XA3.MP2.G SUNSAR_SAR8B_CV_0.XB1.CKN.t4 589.284
R12551 SUNSAR_SAR8B_CV_0.XB1.CKN.n7 SUNSAR_SAR8B_CV_0.XB1.CKN.t7 572.876
R12552 SUNSAR_SAR8B_CV_0.XB1.CKN.n3 SUNSAR_SAR8B_CV_0.XB1.CKN.t6 572.859
R12553 SUNSAR_SAR8B_CV_0.XB1.CKN.n1 SUNSAR_SAR8B_CV_0.XB1.CKN.t3 568.956
R12554 SUNSAR_SAR8B_CV_0.XB1.CKN.t2 SUNSAR_SAR8B_CV_0.XB1.CKN.n2 568.956
R12555 SUNSAR_SAR8B_CV_0.XB1.CKN.n0 SUNSAR_SAR8B_CV_0.XB1.CKN.t1 356.344
R12556 SUNSAR_SAR8B_CV_0.XB1.CKN.n8 SUNSAR_SAR8B_CV_0.XB1.CKN.t0 133.934
R12557 SUNSAR_SAR8B_CV_0.XB1.XA0.MN0.D SUNSAR_SAR8B_CV_0.XB1.CKN.n6 115.954
R12558 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA3.MP2.G 88.8476
R12559 SUNSAR_SAR8B_CV_0.XB1.CKN.n1 SUNSAR_SAR8B_CV_0.XB1.XA3.MN1.G 20.3299
R12560 SUNSAR_SAR8B_CV_0.XB1.CKN.n2 SUNSAR_SAR8B_CV_0.XB1.CKN.n1 20.3299
R12561 SUNSAR_SAR8B_CV_0.XB1.CKN.n2 SUNSAR_SAR8B_CV_0.XB1.XA3.MN0.G 20.3299
R12562 SUNSAR_SAR8B_CV_0.XB1.CKN.n8 SUNSAR_SAR8B_CV_0.XB1.CKN.n7 17.4212
R12563 SUNSAR_SAR8B_CV_0.XB1.CKN.n3 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.G 15.2303
R12564 SUNSAR_SAR8B_CV_0.XB1.CKN.n7 SUNSAR_SAR8B_CV_0.XB1.XA4.MN0.G 15.2129
R12565 SUNSAR_SAR8B_CV_0.XB1.CKN.n4 SUNSAR_SAR8B_CV_0.XB1.XA0.MP0.D 13.5534
R12566 SUNSAR_SAR8B_CV_0.XB1.CKN.n6 SUNSAR_SAR8B_CV_0.XB1.CKN.n0 12.8005
R12567 SUNSAR_SAR8B_CV_0.XB1.CKN.n6 SUNSAR_SAR8B_CV_0.XB1.CKN.n5 9.49168
R12568 SUNSAR_SAR8B_CV_0.XB1.CKN.n5 SUNSAR_SAR8B_CV_0.XB1.CKN.n4 9.3005
R12569 SUNSAR_SAR8B_CV_0.XB1.CKN.n4 SUNSAR_SAR8B_CV_0.XB1.CKN.n0 6.77697
R12570 SUNSAR_SAR8B_CV_0.XB1.CKN.n5 SUNSAR_SAR8B_CV_0.XB1.CKN.n3 6.43121
R12571 SUNSAR_SAR8B_CV_0.XB1.CKN.n9 SUNSAR_SAR8B_CV_0.XB1.CKN.n8 6.35381
R12572 SUNSAR_SAR8B_CV_0.XB1.CKN.n9 SUNSAR_SAR8B_CV_0.XB1.XA0.MN0.D 6.02403
R12573 SUNSAR_SAR8B_CV_0.XB1.XA0.MN0.D SUNSAR_SAR8B_CV_0.XB1.CKN.n9 4.01619
R12574 SUNSAR_SAR8B_CV_0.SARP.n87 SUNSAR_SAR8B_CV_0.SARP.t13 568.956
R12575 SUNSAR_SAR8B_CV_0.SARP.n83 SUNSAR_SAR8B_CV_0.SARP.t12 568.956
R12576 SUNSAR_SAR8B_CV_0.SARP.n84 SUNSAR_SAR8B_CV_0.SARP.t8 568.956
R12577 SUNSAR_SAR8B_CV_0.SARP.n85 SUNSAR_SAR8B_CV_0.SARP.t11 568.956
R12578 SUNSAR_SAR8B_CV_0.SARP.n86 SUNSAR_SAR8B_CV_0.SARP.t14 568.956
R12579 SUNSAR_SAR8B_CV_0.SARP.n81 SUNSAR_SAR8B_CV_0.SARP.t9 568.956
R12580 SUNSAR_SAR8B_CV_0.SARP.n77 SUNSAR_SAR8B_CV_0.SARP.t17 568.956
R12581 SUNSAR_SAR8B_CV_0.SARP.n78 SUNSAR_SAR8B_CV_0.SARP.t15 568.956
R12582 SUNSAR_SAR8B_CV_0.SARP.n79 SUNSAR_SAR8B_CV_0.SARP.t16 568.956
R12583 SUNSAR_SAR8B_CV_0.SARP.n80 SUNSAR_SAR8B_CV_0.SARP.t10 568.956
R12584 SUNSAR_SAR8B_CV_0.XB1.M1.S SUNSAR_SAR8B_CV_0.SARP.t2 151.719
R12585 SUNSAR_SAR8B_CV_0.XB1.M2.S SUNSAR_SAR8B_CV_0.SARP.t1 151.719
R12586 SUNSAR_SAR8B_CV_0.XB1.M3.S SUNSAR_SAR8B_CV_0.SARP.t3 151.719
R12587 SUNSAR_SAR8B_CV_0.SARP.n9 SUNSAR_SAR8B_CV_0.SARP.t6 131.389
R12588 SUNSAR_SAR8B_CV_0.SARP.n3 SUNSAR_SAR8B_CV_0.SARP.t4 131.389
R12589 SUNSAR_SAR8B_CV_0.SARP.n4 SUNSAR_SAR8B_CV_0.SARP.t5 131.389
R12590 SUNSAR_SAR8B_CV_0.SARP.n6 SUNSAR_SAR8B_CV_0.SARP.t7 131.389
R12591 SUNSAR_SAR8B_CV_0.SARP.n0 SUNSAR_SAR8B_CV_0.SARP.t0 131.389
R12592 SUNSAR_SAR8B_CV_0.SARP.n5 SUNSAR_SAR8B_CV_0.SARP.n3 91.4829
R12593 SUNSAR_SAR8B_CV_0.SARP.n8 SUNSAR_SAR8B_CV_0.SARP.n7 84.7064
R12594 SUNSAR_SAR8B_CV_0.SARP.n192 SUNSAR_SAR8B_CV_0.XB1.M1.S 71.1534
R12595 SUNSAR_SAR8B_CV_0.XB1.M4.S SUNSAR_SAR8B_CV_0.SARP.n193 71.1534
R12596 SUNSAR_SAR8B_CV_0.SARP.n7 SUNSAR_SAR8B_CV_0.SARP.n5 53.4593
R12597 SUNSAR_SAR8B_CV_0.SARP.n193 SUNSAR_SAR8B_CV_0.SARP.n192 53.4593
R12598 SUNSAR_SAR8B_CV_0.SARP.n5 SUNSAR_SAR8B_CV_0.SARP.n4 38.024
R12599 SUNSAR_SAR8B_CV_0.SARP.n7 SUNSAR_SAR8B_CV_0.SARP.n6 38.024
R12600 SUNSAR_SAR8B_CV_0.SARP.n121 SUNSAR_SAR8B_CV_0.SARP.n89 24.8589
R12601 SUNSAR_SAR8B_CV_0.SARP.n88 SUNSAR_SAR8B_CV_0.SARP.n87 22.1005
R12602 SUNSAR_SAR8B_CV_0.SARP.n3 SUNSAR_SAR8B_CV_0.XB2.M5.S 20.3299
R12603 SUNSAR_SAR8B_CV_0.SARP.n4 SUNSAR_SAR8B_CV_0.XB2.M6.S 20.3299
R12604 SUNSAR_SAR8B_CV_0.SARP.n6 SUNSAR_SAR8B_CV_0.XB2.M7.S 20.3299
R12605 SUNSAR_SAR8B_CV_0.SARP.n83 SUNSAR_SAR8B_CV_0.XA20.XA1.MN1.G 20.3299
R12606 SUNSAR_SAR8B_CV_0.SARP.n84 SUNSAR_SAR8B_CV_0.SARP.n83 20.3299
R12607 SUNSAR_SAR8B_CV_0.SARP.n84 SUNSAR_SAR8B_CV_0.XA20.XA1.MN2.G 20.3299
R12608 SUNSAR_SAR8B_CV_0.SARP.n85 SUNSAR_SAR8B_CV_0.SARP.n84 20.3299
R12609 SUNSAR_SAR8B_CV_0.SARP.n85 SUNSAR_SAR8B_CV_0.XA20.XA1.MN3.G 20.3299
R12610 SUNSAR_SAR8B_CV_0.SARP.n86 SUNSAR_SAR8B_CV_0.SARP.n85 20.3299
R12611 SUNSAR_SAR8B_CV_0.SARP.n86 SUNSAR_SAR8B_CV_0.XA20.XA1.MN4.G 20.3299
R12612 SUNSAR_SAR8B_CV_0.SARP.n87 SUNSAR_SAR8B_CV_0.SARP.n86 20.3299
R12613 SUNSAR_SAR8B_CV_0.SARP.n77 SUNSAR_SAR8B_CV_0.XA20.XA2.MN5.G 20.3299
R12614 SUNSAR_SAR8B_CV_0.SARP.n78 SUNSAR_SAR8B_CV_0.SARP.n77 20.3299
R12615 SUNSAR_SAR8B_CV_0.SARP.n78 SUNSAR_SAR8B_CV_0.XA20.XA2.MN4.G 20.3299
R12616 SUNSAR_SAR8B_CV_0.SARP.n79 SUNSAR_SAR8B_CV_0.SARP.n78 20.3299
R12617 SUNSAR_SAR8B_CV_0.SARP.n79 SUNSAR_SAR8B_CV_0.XA20.XA2.MN3.G 20.3299
R12618 SUNSAR_SAR8B_CV_0.SARP.n80 SUNSAR_SAR8B_CV_0.SARP.n79 20.3299
R12619 SUNSAR_SAR8B_CV_0.SARP.n80 SUNSAR_SAR8B_CV_0.XA20.XA2.MN2.G 20.3299
R12620 SUNSAR_SAR8B_CV_0.SARP.n81 SUNSAR_SAR8B_CV_0.SARP.n80 20.3299
R12621 SUNSAR_SAR8B_CV_0.SARP.n192 SUNSAR_SAR8B_CV_0.XB1.M2.S 17.6946
R12622 SUNSAR_SAR8B_CV_0.SARP.n193 SUNSAR_SAR8B_CV_0.XB1.M3.S 17.6946
R12623 SUNSAR_SAR8B_CV_0.SARP.n1 SUNSAR_SAR8B_CV_0.SARP.n0 16.077
R12624 SUNSAR_SAR8B_CV_0.SARP.n82 SUNSAR_SAR8B_CV_0.XA20.XA2.MN1.G 15.2303
R12625 SUNSAR_SAR8B_CV_0.SARP.n76 SUNSAR_SAR8B_CV_0.XA20.XA1.MN5.G 13.5534
R12626 SUNSAR_SAR8B_CV_0.SARP.n10 SUNSAR_SAR8B_CV_0.SARP.n9 12.8005
R12627 SUNSAR_SAR8B_CV_0.SARP.n191 SUNSAR_SAR8B_CV_0.SARP.n0 12.8005
R12628 SUNSAR_SAR8B_CV_0.SARP.n11 SUNSAR_SAR8B_CV_0.SARP.n8 9.39466
R12629 SUNSAR_SAR8B_CV_0.SARP.n11 SUNSAR_SAR8B_CV_0.SARP.n10 9.39462
R12630 SUNSAR_SAR8B_CV_0.SARP.n89 SUNSAR_SAR8B_CV_0.SARP.n76 9.36664
R12631 SUNSAR_SAR8B_CV_0.SARP.n191 SUNSAR_SAR8B_CV_0.SARP.n190 9.3005
R12632 SUNSAR_SAR8B_CV_0.SARP.n10 SUNSAR_SAR8B_CV_0.XB2.M8.S 7.52991
R12633 SUNSAR_SAR8B_CV_0.XB1.M4.S SUNSAR_SAR8B_CV_0.SARP.n191 7.52991
R12634 SUNSAR_SAR8B_CV_0.SARP.n88 SUNSAR_SAR8B_CV_0.SARP.n82 7.12974
R12635 SUNSAR_SAR8B_CV_0.SARP.n9 SUNSAR_SAR8B_CV_0.SARP.n8 6.77697
R12636 SUNSAR_SAR8B_CV_0.SARP.n87 SUNSAR_SAR8B_CV_0.SARP.n76 6.77697
R12637 SUNSAR_SAR8B_CV_0.SARP.n12 SUNSAR_SAR8B_CV_0.SARP.n11 5.97637
R12638 SUNSAR_SAR8B_CV_0.SARP.n2 SUNSAR_SAR8B_CV_0.SARP.n1 4.5005
R12639 SUNSAR_SAR8B_CV_0.SARP.n190 SUNSAR_SAR8B_CV_0.SARP.n189 4.5005
R12640 SUNSAR_SAR8B_CV_0.SARP.n82 SUNSAR_SAR8B_CV_0.SARP.n81 3.90429
R12641 SUNSAR_SAR8B_CV_0.SARP.n188 SUNSAR_SAR8B_CV_0.SARP.n187 3.7605
R12642 SUNSAR_SAR8B_CV_0.SARP.n12 SUNSAR_SAR8B_CV_0.SARP.n2 3.4105
R12643 SUNSAR_SAR8B_CV_0.SARP.n189 SUNSAR_SAR8B_CV_0.SARP.n188 3.4105
R12644 SUNSAR_SAR8B_CV_0.SARP.n90 SUNSAR_SAR8B_CV_0.SARP.n44 2.39524
R12645 SUNSAR_SAR8B_CV_0.SARP.n156 SUNSAR_SAR8B_CV_0.SARP.n44 2.39524
R12646 SUNSAR_SAR8B_CV_0.SARP.n187 SUNSAR_SAR8B_CV_0.SARP.n13 2.3035
R12647 SUNSAR_SAR8B_CV_0.SARP.n186 SUNSAR_SAR8B_CV_0.SARP.n14 2.3035
R12648 SUNSAR_SAR8B_CV_0.SARP.n185 SUNSAR_SAR8B_CV_0.SARP.n15 2.3035
R12649 SUNSAR_SAR8B_CV_0.SARP.n184 SUNSAR_SAR8B_CV_0.SARP.n16 2.3035
R12650 SUNSAR_SAR8B_CV_0.SARP.n183 SUNSAR_SAR8B_CV_0.SARP.n17 2.3035
R12651 SUNSAR_SAR8B_CV_0.SARP.n182 SUNSAR_SAR8B_CV_0.SARP.n18 2.3035
R12652 SUNSAR_SAR8B_CV_0.SARP.n181 SUNSAR_SAR8B_CV_0.SARP.n19 2.3035
R12653 SUNSAR_SAR8B_CV_0.SARP.n180 SUNSAR_SAR8B_CV_0.SARP.n20 2.3035
R12654 SUNSAR_SAR8B_CV_0.SARP.n179 SUNSAR_SAR8B_CV_0.SARP.n21 2.3035
R12655 SUNSAR_SAR8B_CV_0.SARP.n178 SUNSAR_SAR8B_CV_0.SARP.n22 2.3035
R12656 SUNSAR_SAR8B_CV_0.SARP.n177 SUNSAR_SAR8B_CV_0.SARP.n23 2.3035
R12657 SUNSAR_SAR8B_CV_0.SARP.n176 SUNSAR_SAR8B_CV_0.SARP.n24 2.3035
R12658 SUNSAR_SAR8B_CV_0.SARP.n175 SUNSAR_SAR8B_CV_0.SARP.n25 2.3035
R12659 SUNSAR_SAR8B_CV_0.SARP.n174 SUNSAR_SAR8B_CV_0.SARP.n26 2.3035
R12660 SUNSAR_SAR8B_CV_0.SARP.n173 SUNSAR_SAR8B_CV_0.SARP.n27 2.3035
R12661 SUNSAR_SAR8B_CV_0.SARP.n172 SUNSAR_SAR8B_CV_0.SARP.n28 2.3035
R12662 SUNSAR_SAR8B_CV_0.SARP.n171 SUNSAR_SAR8B_CV_0.SARP.n29 2.3035
R12663 SUNSAR_SAR8B_CV_0.SARP.n170 SUNSAR_SAR8B_CV_0.SARP.n30 2.3035
R12664 SUNSAR_SAR8B_CV_0.SARP.n169 SUNSAR_SAR8B_CV_0.SARP.n31 2.3035
R12665 SUNSAR_SAR8B_CV_0.SARP.n168 SUNSAR_SAR8B_CV_0.SARP.n32 2.3035
R12666 SUNSAR_SAR8B_CV_0.SARP.n167 SUNSAR_SAR8B_CV_0.SARP.n33 2.3035
R12667 SUNSAR_SAR8B_CV_0.SARP.n166 SUNSAR_SAR8B_CV_0.SARP.n34 2.3035
R12668 SUNSAR_SAR8B_CV_0.SARP.n165 SUNSAR_SAR8B_CV_0.SARP.n35 2.3035
R12669 SUNSAR_SAR8B_CV_0.SARP.n164 SUNSAR_SAR8B_CV_0.SARP.n36 2.3035
R12670 SUNSAR_SAR8B_CV_0.SARP.n163 SUNSAR_SAR8B_CV_0.SARP.n37 2.3035
R12671 SUNSAR_SAR8B_CV_0.SARP.n162 SUNSAR_SAR8B_CV_0.SARP.n38 2.3035
R12672 SUNSAR_SAR8B_CV_0.SARP.n161 SUNSAR_SAR8B_CV_0.SARP.n39 2.3035
R12673 SUNSAR_SAR8B_CV_0.SARP.n160 SUNSAR_SAR8B_CV_0.SARP.n40 2.3035
R12674 SUNSAR_SAR8B_CV_0.SARP.n159 SUNSAR_SAR8B_CV_0.SARP.n41 2.3035
R12675 SUNSAR_SAR8B_CV_0.SARP.n158 SUNSAR_SAR8B_CV_0.SARP.n42 2.3035
R12676 SUNSAR_SAR8B_CV_0.SARP.n157 SUNSAR_SAR8B_CV_0.SARP.n43 2.3035
R12677 SUNSAR_SAR8B_CV_0.SARP.n123 SUNSAR_SAR8B_CV_0.SARP.n13 2.3035
R12678 SUNSAR_SAR8B_CV_0.SARP.n124 SUNSAR_SAR8B_CV_0.SARP.n14 2.3035
R12679 SUNSAR_SAR8B_CV_0.SARP.n125 SUNSAR_SAR8B_CV_0.SARP.n15 2.3035
R12680 SUNSAR_SAR8B_CV_0.SARP.n126 SUNSAR_SAR8B_CV_0.SARP.n16 2.3035
R12681 SUNSAR_SAR8B_CV_0.SARP.n127 SUNSAR_SAR8B_CV_0.SARP.n17 2.3035
R12682 SUNSAR_SAR8B_CV_0.SARP.n128 SUNSAR_SAR8B_CV_0.SARP.n18 2.3035
R12683 SUNSAR_SAR8B_CV_0.SARP.n129 SUNSAR_SAR8B_CV_0.SARP.n19 2.3035
R12684 SUNSAR_SAR8B_CV_0.SARP.n130 SUNSAR_SAR8B_CV_0.SARP.n20 2.3035
R12685 SUNSAR_SAR8B_CV_0.SARP.n131 SUNSAR_SAR8B_CV_0.SARP.n21 2.3035
R12686 SUNSAR_SAR8B_CV_0.SARP.n132 SUNSAR_SAR8B_CV_0.SARP.n22 2.3035
R12687 SUNSAR_SAR8B_CV_0.SARP.n133 SUNSAR_SAR8B_CV_0.SARP.n23 2.3035
R12688 SUNSAR_SAR8B_CV_0.SARP.n134 SUNSAR_SAR8B_CV_0.SARP.n24 2.3035
R12689 SUNSAR_SAR8B_CV_0.SARP.n135 SUNSAR_SAR8B_CV_0.SARP.n25 2.3035
R12690 SUNSAR_SAR8B_CV_0.SARP.n136 SUNSAR_SAR8B_CV_0.SARP.n26 2.3035
R12691 SUNSAR_SAR8B_CV_0.SARP.n137 SUNSAR_SAR8B_CV_0.SARP.n27 2.3035
R12692 SUNSAR_SAR8B_CV_0.SARP.n138 SUNSAR_SAR8B_CV_0.SARP.n28 2.3035
R12693 SUNSAR_SAR8B_CV_0.SARP.n139 SUNSAR_SAR8B_CV_0.SARP.n29 2.3035
R12694 SUNSAR_SAR8B_CV_0.SARP.n140 SUNSAR_SAR8B_CV_0.SARP.n30 2.3035
R12695 SUNSAR_SAR8B_CV_0.SARP.n141 SUNSAR_SAR8B_CV_0.SARP.n31 2.3035
R12696 SUNSAR_SAR8B_CV_0.SARP.n142 SUNSAR_SAR8B_CV_0.SARP.n32 2.3035
R12697 SUNSAR_SAR8B_CV_0.SARP.n143 SUNSAR_SAR8B_CV_0.SARP.n33 2.3035
R12698 SUNSAR_SAR8B_CV_0.SARP.n144 SUNSAR_SAR8B_CV_0.SARP.n34 2.3035
R12699 SUNSAR_SAR8B_CV_0.SARP.n145 SUNSAR_SAR8B_CV_0.SARP.n35 2.3035
R12700 SUNSAR_SAR8B_CV_0.SARP.n146 SUNSAR_SAR8B_CV_0.SARP.n36 2.3035
R12701 SUNSAR_SAR8B_CV_0.SARP.n147 SUNSAR_SAR8B_CV_0.SARP.n37 2.3035
R12702 SUNSAR_SAR8B_CV_0.SARP.n148 SUNSAR_SAR8B_CV_0.SARP.n38 2.3035
R12703 SUNSAR_SAR8B_CV_0.SARP.n149 SUNSAR_SAR8B_CV_0.SARP.n39 2.3035
R12704 SUNSAR_SAR8B_CV_0.SARP.n150 SUNSAR_SAR8B_CV_0.SARP.n40 2.3035
R12705 SUNSAR_SAR8B_CV_0.SARP.n151 SUNSAR_SAR8B_CV_0.SARP.n41 2.3035
R12706 SUNSAR_SAR8B_CV_0.SARP.n152 SUNSAR_SAR8B_CV_0.SARP.n42 2.3035
R12707 SUNSAR_SAR8B_CV_0.SARP.n153 SUNSAR_SAR8B_CV_0.SARP.n43 2.3035
R12708 SUNSAR_SAR8B_CV_0.SARP.n123 SUNSAR_SAR8B_CV_0.SARP.n122 2.3035
R12709 SUNSAR_SAR8B_CV_0.SARP.n124 SUNSAR_SAR8B_CV_0.SARP.n75 2.3035
R12710 SUNSAR_SAR8B_CV_0.SARP.n125 SUNSAR_SAR8B_CV_0.SARP.n74 2.3035
R12711 SUNSAR_SAR8B_CV_0.SARP.n126 SUNSAR_SAR8B_CV_0.SARP.n73 2.3035
R12712 SUNSAR_SAR8B_CV_0.SARP.n127 SUNSAR_SAR8B_CV_0.SARP.n72 2.3035
R12713 SUNSAR_SAR8B_CV_0.SARP.n128 SUNSAR_SAR8B_CV_0.SARP.n71 2.3035
R12714 SUNSAR_SAR8B_CV_0.SARP.n129 SUNSAR_SAR8B_CV_0.SARP.n70 2.3035
R12715 SUNSAR_SAR8B_CV_0.SARP.n130 SUNSAR_SAR8B_CV_0.SARP.n69 2.3035
R12716 SUNSAR_SAR8B_CV_0.SARP.n131 SUNSAR_SAR8B_CV_0.SARP.n68 2.3035
R12717 SUNSAR_SAR8B_CV_0.SARP.n132 SUNSAR_SAR8B_CV_0.SARP.n67 2.3035
R12718 SUNSAR_SAR8B_CV_0.SARP.n133 SUNSAR_SAR8B_CV_0.SARP.n66 2.3035
R12719 SUNSAR_SAR8B_CV_0.SARP.n134 SUNSAR_SAR8B_CV_0.SARP.n65 2.3035
R12720 SUNSAR_SAR8B_CV_0.SARP.n135 SUNSAR_SAR8B_CV_0.SARP.n64 2.3035
R12721 SUNSAR_SAR8B_CV_0.SARP.n136 SUNSAR_SAR8B_CV_0.SARP.n63 2.3035
R12722 SUNSAR_SAR8B_CV_0.SARP.n137 SUNSAR_SAR8B_CV_0.SARP.n62 2.3035
R12723 SUNSAR_SAR8B_CV_0.SARP.n138 SUNSAR_SAR8B_CV_0.SARP.n61 2.3035
R12724 SUNSAR_SAR8B_CV_0.SARP.n139 SUNSAR_SAR8B_CV_0.SARP.n60 2.3035
R12725 SUNSAR_SAR8B_CV_0.SARP.n140 SUNSAR_SAR8B_CV_0.SARP.n59 2.3035
R12726 SUNSAR_SAR8B_CV_0.SARP.n141 SUNSAR_SAR8B_CV_0.SARP.n58 2.3035
R12727 SUNSAR_SAR8B_CV_0.SARP.n142 SUNSAR_SAR8B_CV_0.SARP.n57 2.3035
R12728 SUNSAR_SAR8B_CV_0.SARP.n143 SUNSAR_SAR8B_CV_0.SARP.n56 2.3035
R12729 SUNSAR_SAR8B_CV_0.SARP.n144 SUNSAR_SAR8B_CV_0.SARP.n55 2.3035
R12730 SUNSAR_SAR8B_CV_0.SARP.n145 SUNSAR_SAR8B_CV_0.SARP.n54 2.3035
R12731 SUNSAR_SAR8B_CV_0.SARP.n146 SUNSAR_SAR8B_CV_0.SARP.n53 2.3035
R12732 SUNSAR_SAR8B_CV_0.SARP.n147 SUNSAR_SAR8B_CV_0.SARP.n52 2.3035
R12733 SUNSAR_SAR8B_CV_0.SARP.n148 SUNSAR_SAR8B_CV_0.SARP.n51 2.3035
R12734 SUNSAR_SAR8B_CV_0.SARP.n149 SUNSAR_SAR8B_CV_0.SARP.n50 2.3035
R12735 SUNSAR_SAR8B_CV_0.SARP.n150 SUNSAR_SAR8B_CV_0.SARP.n49 2.3035
R12736 SUNSAR_SAR8B_CV_0.SARP.n151 SUNSAR_SAR8B_CV_0.SARP.n48 2.3035
R12737 SUNSAR_SAR8B_CV_0.SARP.n152 SUNSAR_SAR8B_CV_0.SARP.n47 2.3035
R12738 SUNSAR_SAR8B_CV_0.SARP.n153 SUNSAR_SAR8B_CV_0.SARP.n46 2.3035
R12739 SUNSAR_SAR8B_CV_0.SARP.n122 SUNSAR_SAR8B_CV_0.SARP.n121 2.3035
R12740 SUNSAR_SAR8B_CV_0.SARP.n91 SUNSAR_SAR8B_CV_0.SARP.n46 2.3035
R12741 SUNSAR_SAR8B_CV_0.SARP.n92 SUNSAR_SAR8B_CV_0.SARP.n47 2.3035
R12742 SUNSAR_SAR8B_CV_0.SARP.n93 SUNSAR_SAR8B_CV_0.SARP.n48 2.3035
R12743 SUNSAR_SAR8B_CV_0.SARP.n94 SUNSAR_SAR8B_CV_0.SARP.n49 2.3035
R12744 SUNSAR_SAR8B_CV_0.SARP.n95 SUNSAR_SAR8B_CV_0.SARP.n50 2.3035
R12745 SUNSAR_SAR8B_CV_0.SARP.n96 SUNSAR_SAR8B_CV_0.SARP.n51 2.3035
R12746 SUNSAR_SAR8B_CV_0.SARP.n97 SUNSAR_SAR8B_CV_0.SARP.n52 2.3035
R12747 SUNSAR_SAR8B_CV_0.SARP.n98 SUNSAR_SAR8B_CV_0.SARP.n53 2.3035
R12748 SUNSAR_SAR8B_CV_0.SARP.n99 SUNSAR_SAR8B_CV_0.SARP.n54 2.3035
R12749 SUNSAR_SAR8B_CV_0.SARP.n100 SUNSAR_SAR8B_CV_0.SARP.n55 2.3035
R12750 SUNSAR_SAR8B_CV_0.SARP.n101 SUNSAR_SAR8B_CV_0.SARP.n56 2.3035
R12751 SUNSAR_SAR8B_CV_0.SARP.n102 SUNSAR_SAR8B_CV_0.SARP.n57 2.3035
R12752 SUNSAR_SAR8B_CV_0.SARP.n103 SUNSAR_SAR8B_CV_0.SARP.n58 2.3035
R12753 SUNSAR_SAR8B_CV_0.SARP.n104 SUNSAR_SAR8B_CV_0.SARP.n59 2.3035
R12754 SUNSAR_SAR8B_CV_0.SARP.n105 SUNSAR_SAR8B_CV_0.SARP.n60 2.3035
R12755 SUNSAR_SAR8B_CV_0.SARP.n106 SUNSAR_SAR8B_CV_0.SARP.n61 2.3035
R12756 SUNSAR_SAR8B_CV_0.SARP.n107 SUNSAR_SAR8B_CV_0.SARP.n62 2.3035
R12757 SUNSAR_SAR8B_CV_0.SARP.n108 SUNSAR_SAR8B_CV_0.SARP.n63 2.3035
R12758 SUNSAR_SAR8B_CV_0.SARP.n109 SUNSAR_SAR8B_CV_0.SARP.n64 2.3035
R12759 SUNSAR_SAR8B_CV_0.SARP.n110 SUNSAR_SAR8B_CV_0.SARP.n65 2.3035
R12760 SUNSAR_SAR8B_CV_0.SARP.n111 SUNSAR_SAR8B_CV_0.SARP.n66 2.3035
R12761 SUNSAR_SAR8B_CV_0.SARP.n112 SUNSAR_SAR8B_CV_0.SARP.n67 2.3035
R12762 SUNSAR_SAR8B_CV_0.SARP.n113 SUNSAR_SAR8B_CV_0.SARP.n68 2.3035
R12763 SUNSAR_SAR8B_CV_0.SARP.n114 SUNSAR_SAR8B_CV_0.SARP.n69 2.3035
R12764 SUNSAR_SAR8B_CV_0.SARP.n115 SUNSAR_SAR8B_CV_0.SARP.n70 2.3035
R12765 SUNSAR_SAR8B_CV_0.SARP.n116 SUNSAR_SAR8B_CV_0.SARP.n71 2.3035
R12766 SUNSAR_SAR8B_CV_0.SARP.n117 SUNSAR_SAR8B_CV_0.SARP.n72 2.3035
R12767 SUNSAR_SAR8B_CV_0.SARP.n118 SUNSAR_SAR8B_CV_0.SARP.n73 2.3035
R12768 SUNSAR_SAR8B_CV_0.SARP.n119 SUNSAR_SAR8B_CV_0.SARP.n74 2.3035
R12769 SUNSAR_SAR8B_CV_0.SARP.n120 SUNSAR_SAR8B_CV_0.SARP.n75 2.3035
R12770 SUNSAR_SAR8B_CV_0.SARP.n154 SUNSAR_SAR8B_CV_0.SARP.n45 2.3035
R12771 SUNSAR_SAR8B_CV_0.SARP.n155 SUNSAR_SAR8B_CV_0.SARP.n154 2.3035
R12772 SUNSAR_SAR8B_CV_0.SARP.n91 SUNSAR_SAR8B_CV_0.SARP.n90 1.33497
R12773 SUNSAR_SAR8B_CV_0.SARP.n157 SUNSAR_SAR8B_CV_0.SARP.n156 1.33497
R12774 SUNSAR_SAR8B_CV_0.SARP.n189 SUNSAR_SAR8B_CV_0.SARP.n2 0.191676
R12775 SUNSAR_SAR8B_CV_0.SARP.n190 SUNSAR_SAR8B_CV_0.SARP.n1 0.191676
R12776 SUNSAR_SAR8B_CV_0.SARP.n120 SUNSAR_SAR8B_CV_0.SARP.n119 0.182971
R12777 SUNSAR_SAR8B_CV_0.SARP.n119 SUNSAR_SAR8B_CV_0.SARP.n118 0.182971
R12778 SUNSAR_SAR8B_CV_0.SARP.n118 SUNSAR_SAR8B_CV_0.SARP.n117 0.182971
R12779 SUNSAR_SAR8B_CV_0.SARP.n117 SUNSAR_SAR8B_CV_0.SARP.n116 0.182971
R12780 SUNSAR_SAR8B_CV_0.SARP.n116 SUNSAR_SAR8B_CV_0.SARP.n115 0.182971
R12781 SUNSAR_SAR8B_CV_0.SARP.n115 SUNSAR_SAR8B_CV_0.SARP.n114 0.182971
R12782 SUNSAR_SAR8B_CV_0.SARP.n114 SUNSAR_SAR8B_CV_0.SARP.n113 0.182971
R12783 SUNSAR_SAR8B_CV_0.SARP.n113 SUNSAR_SAR8B_CV_0.SARP.n112 0.182971
R12784 SUNSAR_SAR8B_CV_0.SARP.n112 SUNSAR_SAR8B_CV_0.SARP.n111 0.182971
R12785 SUNSAR_SAR8B_CV_0.SARP.n111 SUNSAR_SAR8B_CV_0.SARP.n110 0.182971
R12786 SUNSAR_SAR8B_CV_0.SARP.n110 SUNSAR_SAR8B_CV_0.SARP.n109 0.182971
R12787 SUNSAR_SAR8B_CV_0.SARP.n109 SUNSAR_SAR8B_CV_0.SARP.n108 0.182971
R12788 SUNSAR_SAR8B_CV_0.SARP.n108 SUNSAR_SAR8B_CV_0.SARP.n107 0.182971
R12789 SUNSAR_SAR8B_CV_0.SARP.n107 SUNSAR_SAR8B_CV_0.SARP.n106 0.182971
R12790 SUNSAR_SAR8B_CV_0.SARP.n106 SUNSAR_SAR8B_CV_0.SARP.n105 0.182971
R12791 SUNSAR_SAR8B_CV_0.SARP.n105 SUNSAR_SAR8B_CV_0.SARP.n104 0.182971
R12792 SUNSAR_SAR8B_CV_0.SARP.n104 SUNSAR_SAR8B_CV_0.SARP.n103 0.182971
R12793 SUNSAR_SAR8B_CV_0.SARP.n103 SUNSAR_SAR8B_CV_0.SARP.n102 0.182971
R12794 SUNSAR_SAR8B_CV_0.SARP.n102 SUNSAR_SAR8B_CV_0.SARP.n101 0.182971
R12795 SUNSAR_SAR8B_CV_0.SARP.n101 SUNSAR_SAR8B_CV_0.SARP.n100 0.182971
R12796 SUNSAR_SAR8B_CV_0.SARP.n100 SUNSAR_SAR8B_CV_0.SARP.n99 0.182971
R12797 SUNSAR_SAR8B_CV_0.SARP.n99 SUNSAR_SAR8B_CV_0.SARP.n98 0.182971
R12798 SUNSAR_SAR8B_CV_0.SARP.n98 SUNSAR_SAR8B_CV_0.SARP.n97 0.182971
R12799 SUNSAR_SAR8B_CV_0.SARP.n97 SUNSAR_SAR8B_CV_0.SARP.n96 0.182971
R12800 SUNSAR_SAR8B_CV_0.SARP.n96 SUNSAR_SAR8B_CV_0.SARP.n95 0.182971
R12801 SUNSAR_SAR8B_CV_0.SARP.n95 SUNSAR_SAR8B_CV_0.SARP.n94 0.182971
R12802 SUNSAR_SAR8B_CV_0.SARP.n94 SUNSAR_SAR8B_CV_0.SARP.n93 0.182971
R12803 SUNSAR_SAR8B_CV_0.SARP.n93 SUNSAR_SAR8B_CV_0.SARP.n92 0.182971
R12804 SUNSAR_SAR8B_CV_0.SARP.n92 SUNSAR_SAR8B_CV_0.SARP.n91 0.182971
R12805 SUNSAR_SAR8B_CV_0.SARP.n75 SUNSAR_SAR8B_CV_0.SARP.n74 0.182971
R12806 SUNSAR_SAR8B_CV_0.SARP.n74 SUNSAR_SAR8B_CV_0.SARP.n73 0.182971
R12807 SUNSAR_SAR8B_CV_0.SARP.n73 SUNSAR_SAR8B_CV_0.SARP.n72 0.182971
R12808 SUNSAR_SAR8B_CV_0.SARP.n72 SUNSAR_SAR8B_CV_0.SARP.n71 0.182971
R12809 SUNSAR_SAR8B_CV_0.SARP.n71 SUNSAR_SAR8B_CV_0.SARP.n70 0.182971
R12810 SUNSAR_SAR8B_CV_0.SARP.n70 SUNSAR_SAR8B_CV_0.SARP.n69 0.182971
R12811 SUNSAR_SAR8B_CV_0.SARP.n69 SUNSAR_SAR8B_CV_0.SARP.n68 0.182971
R12812 SUNSAR_SAR8B_CV_0.SARP.n68 SUNSAR_SAR8B_CV_0.SARP.n67 0.182971
R12813 SUNSAR_SAR8B_CV_0.SARP.n67 SUNSAR_SAR8B_CV_0.SARP.n66 0.182971
R12814 SUNSAR_SAR8B_CV_0.SARP.n66 SUNSAR_SAR8B_CV_0.SARP.n65 0.182971
R12815 SUNSAR_SAR8B_CV_0.SARP.n65 SUNSAR_SAR8B_CV_0.SARP.n64 0.182971
R12816 SUNSAR_SAR8B_CV_0.SARP.n64 SUNSAR_SAR8B_CV_0.SARP.n63 0.182971
R12817 SUNSAR_SAR8B_CV_0.SARP.n63 SUNSAR_SAR8B_CV_0.SARP.n62 0.182971
R12818 SUNSAR_SAR8B_CV_0.SARP.n62 SUNSAR_SAR8B_CV_0.SARP.n61 0.182971
R12819 SUNSAR_SAR8B_CV_0.SARP.n61 SUNSAR_SAR8B_CV_0.SARP.n60 0.182971
R12820 SUNSAR_SAR8B_CV_0.SARP.n60 SUNSAR_SAR8B_CV_0.SARP.n59 0.182971
R12821 SUNSAR_SAR8B_CV_0.SARP.n59 SUNSAR_SAR8B_CV_0.SARP.n58 0.182971
R12822 SUNSAR_SAR8B_CV_0.SARP.n58 SUNSAR_SAR8B_CV_0.SARP.n57 0.182971
R12823 SUNSAR_SAR8B_CV_0.SARP.n57 SUNSAR_SAR8B_CV_0.SARP.n56 0.182971
R12824 SUNSAR_SAR8B_CV_0.SARP.n56 SUNSAR_SAR8B_CV_0.SARP.n55 0.182971
R12825 SUNSAR_SAR8B_CV_0.SARP.n55 SUNSAR_SAR8B_CV_0.SARP.n54 0.182971
R12826 SUNSAR_SAR8B_CV_0.SARP.n54 SUNSAR_SAR8B_CV_0.SARP.n53 0.182971
R12827 SUNSAR_SAR8B_CV_0.SARP.n53 SUNSAR_SAR8B_CV_0.SARP.n52 0.182971
R12828 SUNSAR_SAR8B_CV_0.SARP.n52 SUNSAR_SAR8B_CV_0.SARP.n51 0.182971
R12829 SUNSAR_SAR8B_CV_0.SARP.n51 SUNSAR_SAR8B_CV_0.SARP.n50 0.182971
R12830 SUNSAR_SAR8B_CV_0.SARP.n50 SUNSAR_SAR8B_CV_0.SARP.n49 0.182971
R12831 SUNSAR_SAR8B_CV_0.SARP.n49 SUNSAR_SAR8B_CV_0.SARP.n48 0.182971
R12832 SUNSAR_SAR8B_CV_0.SARP.n48 SUNSAR_SAR8B_CV_0.SARP.n47 0.182971
R12833 SUNSAR_SAR8B_CV_0.SARP.n47 SUNSAR_SAR8B_CV_0.SARP.n46 0.182971
R12834 SUNSAR_SAR8B_CV_0.SARP.n46 SUNSAR_SAR8B_CV_0.SARP.n45 0.182971
R12835 SUNSAR_SAR8B_CV_0.SARP.n125 SUNSAR_SAR8B_CV_0.SARP.n124 0.182971
R12836 SUNSAR_SAR8B_CV_0.SARP.n126 SUNSAR_SAR8B_CV_0.SARP.n125 0.182971
R12837 SUNSAR_SAR8B_CV_0.SARP.n127 SUNSAR_SAR8B_CV_0.SARP.n126 0.182971
R12838 SUNSAR_SAR8B_CV_0.SARP.n128 SUNSAR_SAR8B_CV_0.SARP.n127 0.182971
R12839 SUNSAR_SAR8B_CV_0.SARP.n129 SUNSAR_SAR8B_CV_0.SARP.n128 0.182971
R12840 SUNSAR_SAR8B_CV_0.SARP.n130 SUNSAR_SAR8B_CV_0.SARP.n129 0.182971
R12841 SUNSAR_SAR8B_CV_0.SARP.n131 SUNSAR_SAR8B_CV_0.SARP.n130 0.182971
R12842 SUNSAR_SAR8B_CV_0.SARP.n132 SUNSAR_SAR8B_CV_0.SARP.n131 0.182971
R12843 SUNSAR_SAR8B_CV_0.SARP.n133 SUNSAR_SAR8B_CV_0.SARP.n132 0.182971
R12844 SUNSAR_SAR8B_CV_0.SARP.n134 SUNSAR_SAR8B_CV_0.SARP.n133 0.182971
R12845 SUNSAR_SAR8B_CV_0.SARP.n135 SUNSAR_SAR8B_CV_0.SARP.n134 0.182971
R12846 SUNSAR_SAR8B_CV_0.SARP.n136 SUNSAR_SAR8B_CV_0.SARP.n135 0.182971
R12847 SUNSAR_SAR8B_CV_0.SARP.n137 SUNSAR_SAR8B_CV_0.SARP.n136 0.182971
R12848 SUNSAR_SAR8B_CV_0.SARP.n138 SUNSAR_SAR8B_CV_0.SARP.n137 0.182971
R12849 SUNSAR_SAR8B_CV_0.SARP.n139 SUNSAR_SAR8B_CV_0.SARP.n138 0.182971
R12850 SUNSAR_SAR8B_CV_0.SARP.n140 SUNSAR_SAR8B_CV_0.SARP.n139 0.182971
R12851 SUNSAR_SAR8B_CV_0.SARP.n141 SUNSAR_SAR8B_CV_0.SARP.n140 0.182971
R12852 SUNSAR_SAR8B_CV_0.SARP.n142 SUNSAR_SAR8B_CV_0.SARP.n141 0.182971
R12853 SUNSAR_SAR8B_CV_0.SARP.n143 SUNSAR_SAR8B_CV_0.SARP.n142 0.182971
R12854 SUNSAR_SAR8B_CV_0.SARP.n144 SUNSAR_SAR8B_CV_0.SARP.n143 0.182971
R12855 SUNSAR_SAR8B_CV_0.SARP.n145 SUNSAR_SAR8B_CV_0.SARP.n144 0.182971
R12856 SUNSAR_SAR8B_CV_0.SARP.n146 SUNSAR_SAR8B_CV_0.SARP.n145 0.182971
R12857 SUNSAR_SAR8B_CV_0.SARP.n147 SUNSAR_SAR8B_CV_0.SARP.n146 0.182971
R12858 SUNSAR_SAR8B_CV_0.SARP.n148 SUNSAR_SAR8B_CV_0.SARP.n147 0.182971
R12859 SUNSAR_SAR8B_CV_0.SARP.n149 SUNSAR_SAR8B_CV_0.SARP.n148 0.182971
R12860 SUNSAR_SAR8B_CV_0.SARP.n150 SUNSAR_SAR8B_CV_0.SARP.n149 0.182971
R12861 SUNSAR_SAR8B_CV_0.SARP.n151 SUNSAR_SAR8B_CV_0.SARP.n150 0.182971
R12862 SUNSAR_SAR8B_CV_0.SARP.n152 SUNSAR_SAR8B_CV_0.SARP.n151 0.182971
R12863 SUNSAR_SAR8B_CV_0.SARP.n153 SUNSAR_SAR8B_CV_0.SARP.n152 0.182971
R12864 SUNSAR_SAR8B_CV_0.SARP.n154 SUNSAR_SAR8B_CV_0.SARP.n153 0.182971
R12865 SUNSAR_SAR8B_CV_0.SARP.n154 SUNSAR_SAR8B_CV_0.SARP.n44 0.182971
R12866 SUNSAR_SAR8B_CV_0.SARP.n15 SUNSAR_SAR8B_CV_0.SARP.n14 0.182971
R12867 SUNSAR_SAR8B_CV_0.SARP.n16 SUNSAR_SAR8B_CV_0.SARP.n15 0.182971
R12868 SUNSAR_SAR8B_CV_0.SARP.n17 SUNSAR_SAR8B_CV_0.SARP.n16 0.182971
R12869 SUNSAR_SAR8B_CV_0.SARP.n18 SUNSAR_SAR8B_CV_0.SARP.n17 0.182971
R12870 SUNSAR_SAR8B_CV_0.SARP.n19 SUNSAR_SAR8B_CV_0.SARP.n18 0.182971
R12871 SUNSAR_SAR8B_CV_0.SARP.n20 SUNSAR_SAR8B_CV_0.SARP.n19 0.182971
R12872 SUNSAR_SAR8B_CV_0.SARP.n21 SUNSAR_SAR8B_CV_0.SARP.n20 0.182971
R12873 SUNSAR_SAR8B_CV_0.SARP.n22 SUNSAR_SAR8B_CV_0.SARP.n21 0.182971
R12874 SUNSAR_SAR8B_CV_0.SARP.n23 SUNSAR_SAR8B_CV_0.SARP.n22 0.182971
R12875 SUNSAR_SAR8B_CV_0.SARP.n24 SUNSAR_SAR8B_CV_0.SARP.n23 0.182971
R12876 SUNSAR_SAR8B_CV_0.SARP.n25 SUNSAR_SAR8B_CV_0.SARP.n24 0.182971
R12877 SUNSAR_SAR8B_CV_0.SARP.n26 SUNSAR_SAR8B_CV_0.SARP.n25 0.182971
R12878 SUNSAR_SAR8B_CV_0.SARP.n27 SUNSAR_SAR8B_CV_0.SARP.n26 0.182971
R12879 SUNSAR_SAR8B_CV_0.SARP.n28 SUNSAR_SAR8B_CV_0.SARP.n27 0.182971
R12880 SUNSAR_SAR8B_CV_0.SARP.n29 SUNSAR_SAR8B_CV_0.SARP.n28 0.182971
R12881 SUNSAR_SAR8B_CV_0.SARP.n30 SUNSAR_SAR8B_CV_0.SARP.n29 0.182971
R12882 SUNSAR_SAR8B_CV_0.SARP.n31 SUNSAR_SAR8B_CV_0.SARP.n30 0.182971
R12883 SUNSAR_SAR8B_CV_0.SARP.n32 SUNSAR_SAR8B_CV_0.SARP.n31 0.182971
R12884 SUNSAR_SAR8B_CV_0.SARP.n33 SUNSAR_SAR8B_CV_0.SARP.n32 0.182971
R12885 SUNSAR_SAR8B_CV_0.SARP.n34 SUNSAR_SAR8B_CV_0.SARP.n33 0.182971
R12886 SUNSAR_SAR8B_CV_0.SARP.n35 SUNSAR_SAR8B_CV_0.SARP.n34 0.182971
R12887 SUNSAR_SAR8B_CV_0.SARP.n36 SUNSAR_SAR8B_CV_0.SARP.n35 0.182971
R12888 SUNSAR_SAR8B_CV_0.SARP.n37 SUNSAR_SAR8B_CV_0.SARP.n36 0.182971
R12889 SUNSAR_SAR8B_CV_0.SARP.n38 SUNSAR_SAR8B_CV_0.SARP.n37 0.182971
R12890 SUNSAR_SAR8B_CV_0.SARP.n39 SUNSAR_SAR8B_CV_0.SARP.n38 0.182971
R12891 SUNSAR_SAR8B_CV_0.SARP.n40 SUNSAR_SAR8B_CV_0.SARP.n39 0.182971
R12892 SUNSAR_SAR8B_CV_0.SARP.n41 SUNSAR_SAR8B_CV_0.SARP.n40 0.182971
R12893 SUNSAR_SAR8B_CV_0.SARP.n42 SUNSAR_SAR8B_CV_0.SARP.n41 0.182971
R12894 SUNSAR_SAR8B_CV_0.SARP.n43 SUNSAR_SAR8B_CV_0.SARP.n42 0.182971
R12895 SUNSAR_SAR8B_CV_0.SARP.n155 SUNSAR_SAR8B_CV_0.SARP.n43 0.182971
R12896 SUNSAR_SAR8B_CV_0.SARP.n186 SUNSAR_SAR8B_CV_0.SARP.n185 0.182971
R12897 SUNSAR_SAR8B_CV_0.SARP.n185 SUNSAR_SAR8B_CV_0.SARP.n184 0.182971
R12898 SUNSAR_SAR8B_CV_0.SARP.n184 SUNSAR_SAR8B_CV_0.SARP.n183 0.182971
R12899 SUNSAR_SAR8B_CV_0.SARP.n183 SUNSAR_SAR8B_CV_0.SARP.n182 0.182971
R12900 SUNSAR_SAR8B_CV_0.SARP.n182 SUNSAR_SAR8B_CV_0.SARP.n181 0.182971
R12901 SUNSAR_SAR8B_CV_0.SARP.n181 SUNSAR_SAR8B_CV_0.SARP.n180 0.182971
R12902 SUNSAR_SAR8B_CV_0.SARP.n180 SUNSAR_SAR8B_CV_0.SARP.n179 0.182971
R12903 SUNSAR_SAR8B_CV_0.SARP.n179 SUNSAR_SAR8B_CV_0.SARP.n178 0.182971
R12904 SUNSAR_SAR8B_CV_0.SARP.n178 SUNSAR_SAR8B_CV_0.SARP.n177 0.182971
R12905 SUNSAR_SAR8B_CV_0.SARP.n177 SUNSAR_SAR8B_CV_0.SARP.n176 0.182971
R12906 SUNSAR_SAR8B_CV_0.SARP.n176 SUNSAR_SAR8B_CV_0.SARP.n175 0.182971
R12907 SUNSAR_SAR8B_CV_0.SARP.n175 SUNSAR_SAR8B_CV_0.SARP.n174 0.182971
R12908 SUNSAR_SAR8B_CV_0.SARP.n174 SUNSAR_SAR8B_CV_0.SARP.n173 0.182971
R12909 SUNSAR_SAR8B_CV_0.SARP.n173 SUNSAR_SAR8B_CV_0.SARP.n172 0.182971
R12910 SUNSAR_SAR8B_CV_0.SARP.n172 SUNSAR_SAR8B_CV_0.SARP.n171 0.182971
R12911 SUNSAR_SAR8B_CV_0.SARP.n171 SUNSAR_SAR8B_CV_0.SARP.n170 0.182971
R12912 SUNSAR_SAR8B_CV_0.SARP.n170 SUNSAR_SAR8B_CV_0.SARP.n169 0.182971
R12913 SUNSAR_SAR8B_CV_0.SARP.n169 SUNSAR_SAR8B_CV_0.SARP.n168 0.182971
R12914 SUNSAR_SAR8B_CV_0.SARP.n168 SUNSAR_SAR8B_CV_0.SARP.n167 0.182971
R12915 SUNSAR_SAR8B_CV_0.SARP.n167 SUNSAR_SAR8B_CV_0.SARP.n166 0.182971
R12916 SUNSAR_SAR8B_CV_0.SARP.n166 SUNSAR_SAR8B_CV_0.SARP.n165 0.182971
R12917 SUNSAR_SAR8B_CV_0.SARP.n165 SUNSAR_SAR8B_CV_0.SARP.n164 0.182971
R12918 SUNSAR_SAR8B_CV_0.SARP.n164 SUNSAR_SAR8B_CV_0.SARP.n163 0.182971
R12919 SUNSAR_SAR8B_CV_0.SARP.n163 SUNSAR_SAR8B_CV_0.SARP.n162 0.182971
R12920 SUNSAR_SAR8B_CV_0.SARP.n162 SUNSAR_SAR8B_CV_0.SARP.n161 0.182971
R12921 SUNSAR_SAR8B_CV_0.SARP.n161 SUNSAR_SAR8B_CV_0.SARP.n160 0.182971
R12922 SUNSAR_SAR8B_CV_0.SARP.n160 SUNSAR_SAR8B_CV_0.SARP.n159 0.182971
R12923 SUNSAR_SAR8B_CV_0.SARP.n159 SUNSAR_SAR8B_CV_0.SARP.n158 0.182971
R12924 SUNSAR_SAR8B_CV_0.SARP.n158 SUNSAR_SAR8B_CV_0.SARP.n157 0.182971
R12925 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP SUNSAR_SAR8B_CV_0.SARP.n120 0.159471
R12926 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP SUNSAR_SAR8B_CV_0.SARP.n75 0.159471
R12927 SUNSAR_SAR8B_CV_0.SARP.n124 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.CTOP 0.159471
R12928 SUNSAR_SAR8B_CV_0.SARP.n14 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.CTOP 0.159471
R12929 SUNSAR_SAR8B_CV_0.XDAC1.XC1.CTOP SUNSAR_SAR8B_CV_0.SARP.n186 0.159471
R12930 SUNSAR_SAR8B_CV_0.SARP.n89 SUNSAR_SAR8B_CV_0.SARP.n88 0.124665
R12931 SUNSAR_SAR8B_CV_0.SARP.n90 SUNSAR_SAR8B_CV_0.SARP.n45 0.0855373
R12932 SUNSAR_SAR8B_CV_0.SARP.n156 SUNSAR_SAR8B_CV_0.SARP.n155 0.0855373
R12933 SUNSAR_SAR8B_CV_0.SARP.n188 SUNSAR_SAR8B_CV_0.SARP.n12 0.0723824
R12934 SUNSAR_SAR8B_CV_0.SARP.n187 SUNSAR_SAR8B_CV_0.XDAC1.XC1.CTOP 0.0475
R12935 SUNSAR_SAR8B_CV_0.SARP.n13 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.CTOP 0.0475
R12936 SUNSAR_SAR8B_CV_0.SARP.n123 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.CTOP 0.0475
R12937 SUNSAR_SAR8B_CV_0.SARP.n122 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP 0.0475
R12938 SUNSAR_SAR8B_CV_0.SARP.n121 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP 0.024
R12939 SUNSAR_SAR8B_CV_0.SARP.n122 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP 0.024
R12940 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.CTOP SUNSAR_SAR8B_CV_0.SARP.n123 0.024
R12941 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.CTOP SUNSAR_SAR8B_CV_0.SARP.n13 0.024
R12942 SUNSAR_SAR8B_CV_0.SARP.n187 SUNSAR_SAR8B_CV_0.XDAC1.XC1.CTOP 0.024
R12943 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t6 1060.4
R12944 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XF11.XA2.MN0.G 589.284
R12945 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t4 583.638
R12946 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t2 574.318
R12947 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t3 574.318
R12948 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t5 574.318
R12949 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t7 568.956
R12950 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t1 356.344
R12951 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.t0 131.389
R12952 SUNSAR_CAPT8B_CV_0.XF11.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n16 121.977
R12953 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n8 83.9534
R12954 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n4 16.077
R12955 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n3 12.8005
R12956 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n0 12.8005
R12957 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n12 12.8005
R12958 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.G 10.6968
R12959 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.G 10.6968
R12960 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.G 10.6968
R12961 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n15 9.49168
R12962 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n10 9.49168
R12963 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n2 9.3005
R12964 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n9 9.3005
R12965 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n14 9.3005
R12966 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n1 7.67644
R12967 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.G 7.52991
R12968 SUNSAR_CAPT8B_CV_0.XF11.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n11 7.52991
R12969 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XF11.XA1.MN0.D 7.52991
R12970 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n0 6.77697
R12971 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n12 6.77697
R12972 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n13 5.78673
R12973 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XF11.XA2.MP0.G 5.64756
R12974 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n6 4.28306
R12975 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n7 3.40124
R12976 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n5 1.79829
R12977 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n2 0.191676
R12978 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t2 1060.4
R12979 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XD09.XA2.MN0.G 589.284
R12980 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t3 583.638
R12981 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t6 574.318
R12982 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t7 574.318
R12983 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t5 574.318
R12984 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t4 568.956
R12985 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t1 356.344
R12986 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.t0 131.389
R12987 SUNSAR_CAPT8B_CV_0.XD09.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n16 121.977
R12988 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n8 83.9534
R12989 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n4 16.077
R12990 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n3 12.8005
R12991 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n0 12.8005
R12992 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n12 12.8005
R12993 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.G 10.6968
R12994 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.G 10.6968
R12995 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.G 10.6968
R12996 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n15 9.49168
R12997 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n10 9.49168
R12998 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n2 9.3005
R12999 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n9 9.3005
R13000 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n14 9.3005
R13001 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n1 7.67644
R13002 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.G 7.52991
R13003 SUNSAR_CAPT8B_CV_0.XD09.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n11 7.52991
R13004 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XD09.XA1.MN0.D 7.52991
R13005 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n0 6.77697
R13006 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n12 6.77697
R13007 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n13 5.78673
R13008 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XD09.XA2.MP0.G 5.64756
R13009 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n6 4.28306
R13010 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n7 3.40124
R13011 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n5 1.79829
R13012 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n2 0.191676
R13013 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t9 1060.4
R13014 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t5 1060.4
R13015 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t7 1060.4
R13016 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t8 1060.4
R13017 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n3 568.956
R13018 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t3 568.956
R13019 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n5 568.956
R13020 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t4 568.956
R13021 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t6 568.956
R13022 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n8 568.956
R13023 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t2 568.956
R13024 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n2 568.956
R13025 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.D SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t0 376.673
R13026 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.t1 131.389
R13027 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.D 121.977
R13028 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n3 20.3299
R13029 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA2.XA4.MP3.G 20.3299
R13030 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA2.XA4.MN3.G 20.3299
R13031 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n2 20.3299
R13032 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n4 20.3299
R13033 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA2.XA4.MN2.G 20.3299
R13034 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA2.XA4.MP2.G 20.3299
R13035 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA2.XA4.MP0.G 20.3299
R13036 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n7 20.3299
R13037 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n6 20.3299
R13038 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA2.XA4.MP1.G 20.3299
R13039 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA2.XA4.MN1.G 20.3299
R13040 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n2 20.3299
R13041 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n0 12.8005
R13042 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA2.XA4.MN0.G 10.6968
R13043 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n1 9.49168
R13044 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n10 9.47055
R13045 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n11 9.3005
R13046 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n12 7.52991
R13047 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n0 6.77697
R13048 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n9 5.36434
R13049 ua[1].n12 ua[1].t0 356.344
R13050 ua[1].n13 ua[1].t5 135.293
R13051 ua[1].n0 ua[1].t3 131.389
R13052 ua[1].n2 ua[1].t8 131.389
R13053 ua[1].n3 ua[1].t6 131.389
R13054 ua[1].n5 ua[1].t7 131.389
R13055 ua[1].n7 ua[1].t9 131.389
R13056 ua[1].n9 ua[1].t1 131.389
R13057 ua[1].n11 ua[1].t4 131.389
R13058 ua[1].n18 ua[1].t2 131.389
R13059 ua[1] ua[1].n12 128.754
R13060 ua[1].n4 ua[1].n2 91.4829
R13061 ua[1].n20 ua[1].n19 84.7064
R13062 ua[1].n6 ua[1].n4 53.4593
R13063 ua[1].n8 ua[1].n6 53.4593
R13064 ua[1].n10 ua[1].n8 53.4593
R13065 ua[1].n17 ua[1].n10 53.4593
R13066 ua[1].n19 ua[1].n17 53.4593
R13067 ua[1].n4 ua[1].n3 38.024
R13068 ua[1].n6 ua[1].n5 38.024
R13069 ua[1].n8 ua[1].n7 38.024
R13070 ua[1].n10 ua[1].n9 38.024
R13071 ua[1].n19 ua[1].n18 38.024
R13072 ua[1].n17 ua[1].n16 25.224
R13073 ua[1].n2 ua[1] 20.3299
R13074 ua[1].n3 ua[1] 20.3299
R13075 ua[1].n5 ua[1] 20.3299
R13076 ua[1].n7 ua[1] 20.3299
R13077 ua[1].n9 ua[1] 20.3299
R13078 ua[1].n12 ua[1] 20.3299
R13079 ua[1].n18 ua[1] 20.3299
R13080 ua[1].n13 ua[1] 15.2303
R13081 ua[1].n1 ua[1] 15.1836
R13082 ua[1].n14 ua[1] 13.5534
R13083 ua[1].n16 ua[1].n11 12.8005
R13084 ua[1].n22 ua[1].n0 12.8005
R13085 ua[1].n16 ua[1].n15 9.49168
R13086 ua[1].n21 ua[1].n20 9.3946
R13087 ua[1].n22 ua[1].n21 9.3946
R13088 ua[1].n15 ua[1].n14 9.3005
R13089 ua[1].n15 ua[1].n13 8.44592
R13090 ua[1] ua[1].n22 7.52991
R13091 ua[1].n14 ua[1].n11 6.77697
R13092 ua[1].n20 ua[1].n0 6.77697
R13093 ua[1].n21 ua[1].n1 2.2042
R13094 ua[1].n1 ua[1] 1.75093
R13095 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n19 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n6 8868.95
R13096 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t11 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t8 1060.4
R13097 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n20 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n19 665.066
R13098 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t8 SUNSAR_SAR8B_CV_0.XB2.TIE_L 589.284
R13099 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n6 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t11 574.383
R13100 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n11 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t6 568.956
R13101 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n8 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t9 568.956
R13102 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n9 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t3 568.956
R13103 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n10 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t2 568.956
R13104 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n3 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t7 568.956
R13105 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n0 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t4 568.956
R13106 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n1 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t5 568.956
R13107 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n2 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t10 568.956
R13108 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n25 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t0 136.817
R13109 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n14 SUNSAR_SAR8B_CV_0.XB1.TIE_L.t1 135.293
R13110 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n9 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n8 53.4593
R13111 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n10 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n9 53.4593
R13112 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n11 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n10 53.4593
R13113 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n1 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n0 53.4593
R13114 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n2 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n1 53.4593
R13115 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n3 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n2 53.4593
R13116 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n8 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13117 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n9 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13118 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n10 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13119 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n0 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13120 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n1 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13121 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n2 SUNSAR_SAR8B_CV_0.XB2.TIE_L 20.3299
R13122 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n14 SUNSAR_SAR8B_CV_0.XB2.TIE_L 15.2303
R13123 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n12 SUNSAR_SAR8B_CV_0.XB2.TIE_L 15.1965
R13124 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n4 SUNSAR_SAR8B_CV_0.XB2.TIE_L 10.6968
R13125 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n6 SUNSAR_SAR8B_CV_0.XB2.TIE_L 10.633
R13126 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.TIE_L.n25 10.633
R13127 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n19 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n18 9.45371
R13128 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n13 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n12 8.05861
R13129 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n5 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n4 6.63232
R13130 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n15 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n14 6.23268
R13131 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n4 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n3 5.36434
R13132 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n25 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n24 4.70885
R13133 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n16 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n15 4.5005
R13134 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n13 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n7 4.5005
R13135 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n22 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n5 4.5005
R13136 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n24 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n23 4.5005
R13137 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n12 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n11 3.93805
R13138 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n18 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n7 3.44644
R13139 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n23 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n20 3.44644
R13140 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n17 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n16 3.4105
R13141 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n22 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n21 3.4105
R13142 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n15 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n13 0.191676
R13143 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n16 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n7 0.191676
R13144 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n23 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n22 0.191676
R13145 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n24 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n5 0.191676
R13146 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n18 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n17 0.0364412
R13147 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n21 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n20 0.0364412
R13148 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n17 SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.0281471
R13149 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n21 SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.0281471
R13150 uo_out[3].t3 uo_out[3].t2 1060.4
R13151 uo_out[3].t2 uo_out[3] 589.284
R13152 uo_out[3].n0 uo_out[3].t3 574.383
R13153 uo_out[3].n1 uo_out[3].t1 361.707
R13154 uo_out[3].n3 uo_out[3].t0 131.389
R13155 uo_out[3].n2 uo_out[3] 118.966
R13156 uo_out[3] uo_out[3].n1 10.6968
R13157 uo_out[3].n0 uo_out[3] 10.633
R13158 uo_out[3].n4 uo_out[3] 10.5417
R13159 uo_out[3].n3 uo_out[3].n2 9.78874
R13160 uo_out[3].n4 uo_out[3].n3 9.78874
R13161 uo_out[3].n1 uo_out[3].n0 9.53185
R13162 uo_out[3].n5 uo_out[3].n2 9.39464
R13163 uo_out[3].n5 uo_out[3].n4 9.39464
R13164 uo_out[3].n6 uo_out[3] 9.15944
R13165 uo_out[3].n6 uo_out[3].n5 2.56815
R13166 uo_out[3] uo_out[3].n6 0.180647
R13167 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t2 1060.4
R13168 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XB07.XA2.MN0.G 589.284
R13169 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t3 583.638
R13170 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t7 574.318
R13171 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t6 574.318
R13172 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t5 574.318
R13173 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t4 568.956
R13174 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t1 356.344
R13175 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.t0 131.389
R13176 SUNSAR_CAPT8B_CV_0.XB07.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n16 121.977
R13177 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n8 83.9534
R13178 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n4 16.077
R13179 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n3 12.8005
R13180 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n0 12.8005
R13181 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n12 12.8005
R13182 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.G 10.6968
R13183 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.G 10.6968
R13184 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.G 10.6968
R13185 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n15 9.49168
R13186 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n10 9.49168
R13187 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n2 9.3005
R13188 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n9 9.3005
R13189 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n14 9.3005
R13190 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n1 7.67644
R13191 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.G 7.52991
R13192 SUNSAR_CAPT8B_CV_0.XB07.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n11 7.52991
R13193 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XB07.XA1.MN0.D 7.52991
R13194 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n0 6.77697
R13195 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n12 6.77697
R13196 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n13 5.78673
R13197 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XB07.XA2.MP0.G 5.64756
R13198 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n6 4.28306
R13199 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n7 3.40124
R13200 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n5 1.79829
R13201 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n2 0.191676
R13202 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t5 1060.4
R13203 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XE10.XA2.MN0.G 589.284
R13204 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t6 572.893
R13205 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t7 572.893
R13206 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t3 572.893
R13207 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t4 568.956
R13208 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t2 568.956
R13209 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t1 356.344
R13210 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.t0 135.293
R13211 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XE10.XA1.MN0.D 115.954
R13212 SUNSAR_CAPT8B_CV_0.XE10.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n13 85.0829
R13213 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n5 22.1005
R13214 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XE10.XA2.MP0.G 20.3299
R13215 SUNSAR_CAPT8B_CV_0.XE10.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n2 15.2303
R13216 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.G 15.1965
R13217 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.G 15.1965
R13218 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.G 15.1965
R13219 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.G 13.5534
R13220 SUNSAR_CAPT8B_CV_0.XE10.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n12 13.5534
R13221 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n0 12.8005
R13222 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n1 12.6805
R13223 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n3 9.49168
R13224 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n7 9.3005
R13225 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n11 9.3005
R13226 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n4 9.10273
R13227 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n6 6.77697
R13228 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n0 6.77697
R13229 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n9 5.70934
R13230 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n10 3.40124
R13231 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n8 1.79829
R13232 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n5 0.191676
R13233 SUNSAR_SAR8B_CV_0.XA3.ENO.t3 SUNSAR_SAR8B_CV_0.XA3.ENO.t4 1060.4
R13234 SUNSAR_SAR8B_CV_0.XA3.ENO.t5 SUNSAR_SAR8B_CV_0.XA3.ENO.t2 1060.4
R13235 SUNSAR_SAR8B_CV_0.XA3.ENO.t4 SUNSAR_SAR8B_CV_0.XA4.EN 589.284
R13236 SUNSAR_SAR8B_CV_0.XA3.ENO.t2 SUNSAR_SAR8B_CV_0.XA4.EN 589.284
R13237 SUNSAR_SAR8B_CV_0.XA3.ENO.n0 SUNSAR_SAR8B_CV_0.XA3.ENO.t3 583.638
R13238 SUNSAR_SAR8B_CV_0.XA3.ENO.n5 SUNSAR_SAR8B_CV_0.XA3.ENO.t8 574.383
R13239 SUNSAR_SAR8B_CV_0.XA3.ENO.n6 SUNSAR_SAR8B_CV_0.XA3.ENO.t6 574.383
R13240 SUNSAR_SAR8B_CV_0.XA3.ENO.n12 SUNSAR_SAR8B_CV_0.XA3.ENO.t5 572.893
R13241 SUNSAR_SAR8B_CV_0.XA3.ENO.n10 SUNSAR_SAR8B_CV_0.XA3.ENO.t7 568.956
R13242 SUNSAR_SAR8B_CV_0.XA3.ENO.n2 SUNSAR_SAR8B_CV_0.XA3.ENO.t1 356.344
R13243 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.ENO.n17 268.8
R13244 SUNSAR_SAR8B_CV_0.XA3.ENO.n1 SUNSAR_SAR8B_CV_0.XA3.ENO.t0 131.389
R13245 SUNSAR_SAR8B_CV_0.XA3.ENO.n1 SUNSAR_SAR8B_CV_0.XA3.ENO.n0 90.7299
R13246 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.ENO.n1 20.3299
R13247 SUNSAR_SAR8B_CV_0.XA3.ENO.n13 SUNSAR_SAR8B_CV_0.XA3.ENO.n12 20.0513
R13248 SUNSAR_SAR8B_CV_0.XA3.ENO.n11 SUNSAR_SAR8B_CV_0.XA3.ENO.n10 16.1445
R13249 SUNSAR_SAR8B_CV_0.XA3.ENO.n12 SUNSAR_SAR8B_CV_0.XA4.EN 15.1965
R13250 SUNSAR_SAR8B_CV_0.XA3.ENO.n3 SUNSAR_SAR8B_CV_0.XA4.EN 13.5534
R13251 SUNSAR_SAR8B_CV_0.XA3.ENO.n10 SUNSAR_SAR8B_CV_0.XA3.ENO.n9 12.8005
R13252 SUNSAR_SAR8B_CV_0.XA3.ENO.n17 SUNSAR_SAR8B_CV_0.XA3.ENO.n2 12.8005
R13253 SUNSAR_SAR8B_CV_0.XA3.ENO.n5 SUNSAR_SAR8B_CV_0.XA4.EN 10.633
R13254 SUNSAR_SAR8B_CV_0.XA3.ENO.n6 SUNSAR_SAR8B_CV_0.XA4.EN 10.633
R13255 SUNSAR_SAR8B_CV_0.XA3.ENO.n17 SUNSAR_SAR8B_CV_0.XA3.ENO.n16 9.35932
R13256 SUNSAR_SAR8B_CV_0.XA3.ENO.n9 SUNSAR_SAR8B_CV_0.XA3.ENO.n8 9.3005
R13257 SUNSAR_SAR8B_CV_0.XA3.ENO.n4 SUNSAR_SAR8B_CV_0.XA3.ENO.n3 9.3005
R13258 SUNSAR_SAR8B_CV_0.XA3.ENO.n9 SUNSAR_SAR8B_CV_0.XA4.EN 7.52991
R13259 SUNSAR_SAR8B_CV_0.XA3.ENO.n3 SUNSAR_SAR8B_CV_0.XA3.ENO.n2 6.77697
R13260 SUNSAR_SAR8B_CV_0.XA3.ENO.n0 SUNSAR_SAR8B_CV_0.XA4.EN 5.64756
R13261 SUNSAR_SAR8B_CV_0.XA3.ENO.n7 SUNSAR_SAR8B_CV_0.XA3.ENO.n5 5.35958
R13262 SUNSAR_SAR8B_CV_0.XA3.ENO.n14 SUNSAR_SAR8B_CV_0.XA3.ENO.n13 4.5005
R13263 SUNSAR_SAR8B_CV_0.XA3.ENO.n16 SUNSAR_SAR8B_CV_0.XA3.ENO.n15 4.5005
R13264 SUNSAR_SAR8B_CV_0.XA3.ENO.n15 SUNSAR_SAR8B_CV_0.XA4.EN 4.33874
R13265 SUNSAR_SAR8B_CV_0.XA3.ENO.n7 SUNSAR_SAR8B_CV_0.XA3.ENO.n6 4.19047
R13266 SUNSAR_SAR8B_CV_0.XA3.ENO.n8 SUNSAR_SAR8B_CV_0.XA3.ENO.n7 4.00418
R13267 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.ENO.n11 2.35274
R13268 SUNSAR_SAR8B_CV_0.XA3.ENO.n15 SUNSAR_SAR8B_CV_0.XA3.ENO.n14 0.191676
R13269 SUNSAR_SAR8B_CV_0.XA3.ENO.n16 SUNSAR_SAR8B_CV_0.XA3.ENO.n4 0.132853
R13270 SUNSAR_SAR8B_CV_0.XA3.ENO.n11 SUNSAR_SAR8B_CV_0.XA3.ENO.n8 0.123303
R13271 SUNSAR_SAR8B_CV_0.XA3.ENO.n14 SUNSAR_SAR8B_CV_0.XA4.EN 0.0740294
R13272 SUNSAR_SAR8B_CV_0.XA3.ENO.n13 SUNSAR_SAR8B_CV_0.XA3.ENO.n4 0.0593235
R13273 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n80 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n79 296.438
R13274 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n72 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n71 91.8472
R13275 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n71 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n68 91.8472
R13276 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n9 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n8 91.8472
R13277 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n8 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n5 91.8472
R13278 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n24 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n23 91.8472
R13279 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n23 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n20 91.8472
R13280 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n40 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n39 91.8472
R13281 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n39 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n36 91.8472
R13282 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n56 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n55 91.8472
R13283 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n55 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n52 91.8472
R13284 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n79 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.t1 63.8431
R13285 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n79 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.t0 63.8431
R13286 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n71 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n70 49.1805
R13287 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n8 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n7 49.1805
R13288 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n23 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n22 49.1805
R13289 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n39 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n38 49.1805
R13290 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n55 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n54 49.1805
R13291 SUNSAR_SAR8B_CV_0.XB1.XA4.MP0.D SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n80 15.1965
R13292 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n80 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n78 10.4602
R13293 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n76 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB0.A 3.99785
R13294 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n13 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB4.A 3.99785
R13295 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n28 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB3.A 3.99785
R13296 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n44 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB2.A 3.99785
R13297 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n60 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB1.A 3.99785
R13298 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n76 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n75 2.03137
R13299 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n13 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n12 2.03137
R13300 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n28 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n27 2.03137
R13301 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n44 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n43 2.03137
R13302 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n60 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n59 2.03137
R13303 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n75 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n74 2.03137
R13304 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n12 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n11 2.03137
R13305 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n27 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n26 2.03137
R13306 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n43 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n42 2.03137
R13307 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n59 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n58 2.03137
R13308 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n75 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n65 1.8747
R13309 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n12 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n2 1.8747
R13310 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n27 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n17 1.8747
R13311 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n43 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n33 1.8747
R13312 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n59 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n49 1.8747
R13313 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n73 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n72 1.5005
R13314 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n68 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n64 1.5005
R13315 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n70 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n69 1.5005
R13316 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n10 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n9 1.5005
R13317 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n5 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n1 1.5005
R13318 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n7 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n6 1.5005
R13319 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n25 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n24 1.5005
R13320 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n20 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n16 1.5005
R13321 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n22 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n21 1.5005
R13322 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n41 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n40 1.5005
R13323 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n36 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n32 1.5005
R13324 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n38 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n37 1.5005
R13325 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n57 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n56 1.5005
R13326 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n52 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n48 1.5005
R13327 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n54 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n53 1.5005
R13328 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n74 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n73 1.13717
R13329 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n69 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n65 1.13717
R13330 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n76 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n64 1.13717
R13331 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n11 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n10 1.13717
R13332 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n6 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n2 1.13717
R13333 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n13 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n1 1.13717
R13334 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n26 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n25 1.13717
R13335 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n21 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n17 1.13717
R13336 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n28 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n16 1.13717
R13337 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n42 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n41 1.13717
R13338 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n37 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n33 1.13717
R13339 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n44 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n32 1.13717
R13340 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n58 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n57 1.13717
R13341 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n53 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n49 1.13717
R13342 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n60 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n48 1.13717
R13343 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n73 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n66 0.867167
R13344 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n72 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n67 0.867167
R13345 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n68 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n67 0.867167
R13346 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n66 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n64 0.867167
R13347 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n10 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n3 0.867167
R13348 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n9 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n4 0.867167
R13349 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n5 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n4 0.867167
R13350 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n3 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n1 0.867167
R13351 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n25 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n18 0.867167
R13352 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n24 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n19 0.867167
R13353 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n20 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n19 0.867167
R13354 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n18 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n16 0.867167
R13355 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n41 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n34 0.867167
R13356 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n40 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n35 0.867167
R13357 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n36 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n35 0.867167
R13358 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n34 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n32 0.867167
R13359 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n57 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n50 0.867167
R13360 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n56 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n51 0.867167
R13361 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n52 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n51 0.867167
R13362 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n50 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n48 0.867167
R13363 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n30 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n14 0.70315
R13364 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n78 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n77 0.646474
R13365 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n46 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n30 0.617029
R13366 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n62 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n46 0.617029
R13367 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n70 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n67 0.4505
R13368 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n69 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n66 0.4505
R13369 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n7 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n4 0.4505
R13370 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n6 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n3 0.4505
R13371 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n22 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n19 0.4505
R13372 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n21 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n18 0.4505
R13373 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n38 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n35 0.4505
R13374 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n37 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n34 0.4505
R13375 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n54 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n51 0.4505
R13376 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n53 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n50 0.4505
R13377 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n74 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n63 0.326367
R13378 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n11 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n0 0.326367
R13379 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n26 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n15 0.326367
R13380 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n42 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n31 0.326367
R13381 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n58 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n47 0.326367
R13382 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n65 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n63 0.1697
R13383 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n77 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n76 0.1697
R13384 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n2 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n0 0.1697
R13385 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n14 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n13 0.1697
R13386 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n17 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n15 0.1697
R13387 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n29 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n28 0.1697
R13388 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n33 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n31 0.1697
R13389 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n45 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n44 0.1697
R13390 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n49 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n47 0.1697
R13391 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n61 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n60 0.1697
R13392 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n77 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n63 0.157167
R13393 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n14 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n0 0.157167
R13394 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n29 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n15 0.157167
R13395 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n45 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n31 0.157167
R13396 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n61 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n47 0.157167
R13397 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n30 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n29 0.0866206
R13398 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n46 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n45 0.0866206
R13399 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n62 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n61 0.0866206
R13400 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n78 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n62 0.0101765
R13401 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t3 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t5 1060.4
R13402 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t5 SUNSAR_CAPT8B_CV_0.XH13.XA2.MN0.G 589.284
R13403 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t3 583.638
R13404 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t6 574.318
R13405 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t4 574.318
R13406 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t7 574.318
R13407 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t2 568.956
R13408 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t1 356.344
R13409 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.t0 131.389
R13410 SUNSAR_CAPT8B_CV_0.XH13.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n16 121.977
R13411 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n8 83.9534
R13412 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n4 16.077
R13413 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n3 12.8005
R13414 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n0 12.8005
R13415 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n12 12.8005
R13416 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.G 10.6968
R13417 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.G 10.6968
R13418 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.G 10.6968
R13419 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n15 9.49168
R13420 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n10 9.49168
R13421 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n2 9.3005
R13422 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n9 9.3005
R13423 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n14 9.3005
R13424 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n1 7.67644
R13425 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.G 7.52991
R13426 SUNSAR_CAPT8B_CV_0.XH13.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n11 7.52991
R13427 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n14 SUNSAR_CAPT8B_CV_0.XH13.XA1.MN0.D 7.52991
R13428 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n0 6.77697
R13429 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n16 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n12 6.77697
R13430 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n15 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n13 5.78673
R13431 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XH13.XA2.MP0.G 5.64756
R13432 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n6 4.28306
R13433 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n7 3.40124
R13434 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n5 1.79829
R13435 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n2 0.191676
R13436 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t2 1060.4
R13437 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t5 1060.4
R13438 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t4 1060.4
R13439 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t8 1060.4
R13440 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n1 568.956
R13441 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t3 568.956
R13442 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n3 568.956
R13443 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t9 568.956
R13444 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t6 568.956
R13445 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n6 568.956
R13446 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t7 568.956
R13447 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n0 568.956
R13448 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t0 356.344
R13449 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.t1 135.293
R13450 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n10 128.754
R13451 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n1 20.3299
R13452 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA3.XA4.MP3.G 20.3299
R13453 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA3.XA4.MN3.G 20.3299
R13454 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n0 20.3299
R13455 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n2 20.3299
R13456 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA3.XA4.MN2.G 20.3299
R13457 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA3.XA4.MP2.G 20.3299
R13458 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA3.XA4.MP0.G 20.3299
R13459 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n5 20.3299
R13460 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n4 20.3299
R13461 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA3.XA4.MP1.G 20.3299
R13462 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA3.XA4.MN1.G 20.3299
R13463 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n0 20.3299
R13464 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.D 20.3299
R13465 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n8 16.3643
R13466 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n9 15.2303
R13467 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA3.XA4.MN0.G 15.1965
R13468 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n7 3.93805
R13469 SUNSAR_SAR8B_CV_0.XA3.CP0.t15 SUNSAR_SAR8B_CV_0.XA3.CP0.t13 1060.4
R13470 SUNSAR_SAR8B_CV_0.XA3.CP0.t11 SUNSAR_SAR8B_CV_0.XA3.CP0.t14 1060.4
R13471 SUNSAR_SAR8B_CV_0.XA3.CP0.t10 SUNSAR_SAR8B_CV_0.XA3.CP0.t12 1060.4
R13472 SUNSAR_SAR8B_CV_0.XA3.CP0.t9 SUNSAR_SAR8B_CV_0.XA3.CP0.t8 1060.4
R13473 SUNSAR_SAR8B_CV_0.XA3.CP0.t13 SUNSAR_SAR8B_CV_0.XA3.CP0.n1 568.956
R13474 SUNSAR_SAR8B_CV_0.XA3.CP0.n2 SUNSAR_SAR8B_CV_0.XA3.CP0.t15 568.956
R13475 SUNSAR_SAR8B_CV_0.XA3.CP0.t14 SUNSAR_SAR8B_CV_0.XA3.CP0.n3 568.956
R13476 SUNSAR_SAR8B_CV_0.XA3.CP0.n4 SUNSAR_SAR8B_CV_0.XA3.CP0.t11 568.956
R13477 SUNSAR_SAR8B_CV_0.XA3.CP0.n7 SUNSAR_SAR8B_CV_0.XA3.CP0.t10 568.956
R13478 SUNSAR_SAR8B_CV_0.XA3.CP0.t12 SUNSAR_SAR8B_CV_0.XA3.CP0.n6 568.956
R13479 SUNSAR_SAR8B_CV_0.XA3.CP0.n5 SUNSAR_SAR8B_CV_0.XA3.CP0.t9 568.956
R13480 SUNSAR_SAR8B_CV_0.XA3.CP0.t8 SUNSAR_SAR8B_CV_0.XA3.CP0.n0 568.956
R13481 SUNSAR_SAR8B_CV_0.XA3.CP0.n12 SUNSAR_SAR8B_CV_0.XA3.CP0.n11 292.5
R13482 SUNSAR_SAR8B_CV_0.XA3.CP0.n15 SUNSAR_SAR8B_CV_0.XA3.CP0.n14 292.5
R13483 SUNSAR_SAR8B_CV_0.XA3.CP0.n9 SUNSAR_SAR8B_CV_0.XA3.CP0 197.272
R13484 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.CP0.n10 112.829
R13485 SUNSAR_SAR8B_CV_0.XA3.CP0.n13 SUNSAR_SAR8B_CV_0.XA3.CP0.n12 111.059
R13486 SUNSAR_SAR8B_CV_0.XA3.CP0.n9 SUNSAR_SAR8B_CV_0.XA3.CP0.n8 92.5005
R13487 SUNSAR_SAR8B_CV_0.XA3.CP0.n16 SUNSAR_SAR8B_CV_0.XA3.CP0.n15 81.5064
R13488 SUNSAR_SAR8B_CV_0.XA3.CP0.n14 SUNSAR_SAR8B_CV_0.XA3.CP0.t4 63.8431
R13489 SUNSAR_SAR8B_CV_0.XA3.CP0.n14 SUNSAR_SAR8B_CV_0.XA3.CP0.t5 63.8431
R13490 SUNSAR_SAR8B_CV_0.XA3.CP0.n11 SUNSAR_SAR8B_CV_0.XA3.CP0.t7 63.8431
R13491 SUNSAR_SAR8B_CV_0.XA3.CP0.n11 SUNSAR_SAR8B_CV_0.XA3.CP0.t6 63.8431
R13492 SUNSAR_SAR8B_CV_0.XA3.CP0.n17 SUNSAR_SAR8B_CV_0.XA3.CP0.n13 53.4593
R13493 SUNSAR_SAR8B_CV_0.XA3.CP0.n10 SUNSAR_SAR8B_CV_0.XA3.CP0.t1 38.8894
R13494 SUNSAR_SAR8B_CV_0.XA3.CP0.n10 SUNSAR_SAR8B_CV_0.XA3.CP0.t2 38.8894
R13495 SUNSAR_SAR8B_CV_0.XA3.CP0.n8 SUNSAR_SAR8B_CV_0.XA3.CP0.t3 38.8894
R13496 SUNSAR_SAR8B_CV_0.XA3.CP0.n8 SUNSAR_SAR8B_CV_0.XA3.CP0.t0 38.8894
R13497 SUNSAR_SAR8B_CV_0.XA3.CP0.n17 SUNSAR_SAR8B_CV_0.XA3.CP0.n16 29.5534
R13498 SUNSAR_SAR8B_CV_0.XA3.CP0.n4 SUNSAR_SAR8B_CV_0.XA3.CP0.n1 20.3299
R13499 SUNSAR_SAR8B_CV_0.XA3.CP0.n1 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13500 SUNSAR_SAR8B_CV_0.XA3.CP0.n2 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13501 SUNSAR_SAR8B_CV_0.XA3.CP0.n3 SUNSAR_SAR8B_CV_0.XA3.CP0.n0 20.3299
R13502 SUNSAR_SAR8B_CV_0.XA3.CP0.n3 SUNSAR_SAR8B_CV_0.XA3.CP0.n2 20.3299
R13503 SUNSAR_SAR8B_CV_0.XA3.CP0.n3 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13504 SUNSAR_SAR8B_CV_0.XA3.CP0.n4 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13505 SUNSAR_SAR8B_CV_0.XA3.CP0.n6 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13506 SUNSAR_SAR8B_CV_0.XA3.CP0.n6 SUNSAR_SAR8B_CV_0.XA3.CP0.n5 20.3299
R13507 SUNSAR_SAR8B_CV_0.XA3.CP0.n5 SUNSAR_SAR8B_CV_0.XA3.CP0.n4 20.3299
R13508 SUNSAR_SAR8B_CV_0.XA3.CP0.n5 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13509 SUNSAR_SAR8B_CV_0.XA3.CP0.n0 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13510 SUNSAR_SAR8B_CV_0.XA3.CP0.n7 SUNSAR_SAR8B_CV_0.XA3.CP0.n0 20.3299
R13511 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.CP0.n7 20.3299
R13512 SUNSAR_SAR8B_CV_0.XA3.CP0.n12 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13513 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.CP0.n9 20.3299
R13514 SUNSAR_SAR8B_CV_0.XA3.CP0.n15 SUNSAR_SAR8B_CV_0.XA3.CP0 20.3299
R13515 SUNSAR_SAR8B_CV_0.XA3.CP0.n13 SUNSAR_SAR8B_CV_0.XA3.CP0 17.6946
R13516 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.CP0.n17 17.6946
R13517 SUNSAR_SAR8B_CV_0.XA3.CP0.n16 SUNSAR_SAR8B_CV_0.XA3.CP0 10.3476
R13518 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t29 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t30 1060.4
R13519 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t26 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t8 1060.4
R13520 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t9 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t12 1060.4
R13521 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t27 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t22 1060.4
R13522 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t16 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t24 1060.4
R13523 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t13 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t23 1060.4
R13524 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t31 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t17 1060.4
R13525 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t14 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t21 1060.4
R13526 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t30 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.G 589.284
R13527 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t8 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.G 589.284
R13528 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.G SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t26 589.284
R13529 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t12 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.G 589.284
R13530 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t22 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.G 589.284
R13531 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.G SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t27 589.284
R13532 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t24 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.G 589.284
R13533 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t23 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.G 589.284
R13534 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.G SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t13 589.284
R13535 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t17 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.G 589.284
R13536 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t21 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.G 589.284
R13537 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.G SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t14 589.284
R13538 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n2 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t20 574.351
R13539 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n8 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t10 574.351
R13540 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n14 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t28 574.351
R13541 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n20 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t15 574.351
R13542 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n30 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t19 568.956
R13543 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n28 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t29 568.956
R13544 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n5 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t18 568.956
R13545 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n4 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t9 568.956
R13546 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n11 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t11 568.956
R13547 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n10 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t16 568.956
R13548 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n17 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t25 568.956
R13549 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n16 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t31 568.956
R13550 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n29 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n28 454.024
R13551 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n6 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n4 454.024
R13552 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n12 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n10 454.024
R13553 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n18 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n16 454.024
R13554 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.G 420.142
R13555 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.G 420.142
R13556 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.G 420.142
R13557 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.G 420.142
R13558 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n0 312.829
R13559 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n35 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n1 297.897
R13560 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n37 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n36 92.5005
R13561 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n40 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n39 92.5005
R13562 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n38 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP0.D 90.7299
R13563 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP2.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n41 90.7299
R13564 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n0 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t3 63.8431
R13565 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n0 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t7 63.8431
R13566 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t4 63.8431
R13567 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n1 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t2 63.8431
R13568 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n41 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n38 53.4593
R13569 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n36 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t1 38.8894
R13570 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n36 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t5 38.8894
R13571 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n39 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t6 38.8894
R13572 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n39 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.t0 38.8894
R13573 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n38 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n37 38.024
R13574 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n41 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n40 38.024
R13575 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n28 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN1.G 20.3299
R13576 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n4 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN1.G 20.3299
R13577 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n10 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN1.G 20.3299
R13578 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n16 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN1.G 20.3299
R13579 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n37 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN0.D 20.3299
R13580 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n40 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN2.D 20.3299
R13581 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n21 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n20 14.4056
R13582 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n31 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n30 12.8005
R13583 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n5 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n3 12.8005
R13584 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n11 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n9 12.8005
R13585 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n17 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n15 12.8005
R13586 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n35 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n34 12.2843
R13587 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n2 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.G 10.664
R13588 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n8 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.G 10.664
R13589 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n14 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.G 10.664
R13590 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n20 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.G 10.664
R13591 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP0.D SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n35 10.664
R13592 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n7 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n6 9.39659
R13593 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n13 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n12 9.39659
R13594 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n19 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n18 9.39659
R13595 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n7 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n3 9.39269
R13596 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n13 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n9 9.39269
R13597 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n19 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n15 9.39269
R13598 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n33 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n29 9.3005
R13599 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n32 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n31 9.3005
R13600 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n27 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n26 8.19535
R13601 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n25 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n24 7.67697
R13602 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n23 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n22 7.67697
R13603 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n31 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN0.G 7.52991
R13604 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n3 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN0.G 7.52991
R13605 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n9 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN0.G 7.52991
R13606 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n15 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN0.G 7.52991
R13607 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n30 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n29 6.77697
R13608 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n6 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n5 6.77697
R13609 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n12 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n11 6.77697
R13610 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n18 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n17 6.77697
R13611 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n26 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n2 6.72914
R13612 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n24 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n8 6.72914
R13613 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n22 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n14 6.72914
R13614 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n34 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n33 4.5005
R13615 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n32 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n27 4.5005
R13616 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n25 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n7 2.76938
R13617 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n23 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n13 2.76938
R13618 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n21 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n19 2.76938
R13619 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n26 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n25 1.58874
R13620 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n24 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n23 1.58874
R13621 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n22 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n21 1.58874
R13622 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n33 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n32 0.191676
R13623 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n34 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n27 0.191676
R13624 uo_out[0].t3 uo_out[0].t2 1060.4
R13625 uo_out[0].t2 uo_out[0] 589.284
R13626 uo_out[0].n1 uo_out[0].t3 572.859
R13627 uo_out[0].n0 uo_out[0].t1 356.344
R13628 uo_out[0].n5 uo_out[0].t0 136.285
R13629 uo_out[0] uo_out[0].n4 115.954
R13630 uo_out[0].n1 uo_out[0] 15.2303
R13631 uo_out[0].n2 uo_out[0] 13.5534
R13632 uo_out[0].n5 uo_out[0] 12.939
R13633 uo_out[0].n4 uo_out[0].n0 12.8005
R13634 uo_out[0].n6 uo_out[0] 10.9838
R13635 uo_out[0].n4 uo_out[0].n3 9.49168
R13636 uo_out[0].n3 uo_out[0].n2 9.3005
R13637 uo_out[0].n6 uo_out[0].n5 7.24734
R13638 uo_out[0].n3 uo_out[0].n1 7.07827
R13639 uo_out[0].n2 uo_out[0].n0 6.77697
R13640 uo_out[0] uo_out[0].n6 0.199029
R13641 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t6 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t15 1060.4
R13642 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t10 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t13 1060.4
R13643 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t7 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t14 1060.4
R13644 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t9 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t12 1060.4
R13645 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t8 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t11 1060.4
R13646 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t15 SUNSAR_SAR8B_CV_0.XA20.XA3.MN6.G 589.284
R13647 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n4 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t16 568.956
R13648 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n2 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t6 568.956
R13649 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t5 568.956
R13650 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t13 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n6 568.956
R13651 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n7 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t10 568.956
R13652 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t14 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n8 568.956
R13653 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n9 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t7 568.956
R13654 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n12 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t9 568.956
R13655 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t12 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n11 568.956
R13656 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n10 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t8 568.956
R13657 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t11 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n5 568.956
R13658 SUNSAR_SAR8B_CV_0.XA20.XA2.MP3.D SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n0 312.829
R13659 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n13 SUNSAR_SAR8B_CV_0.XA20.XA3.MP4.G 308.329
R13660 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n15 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n14 292.5
R13661 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n15 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n13 273.695
R13662 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n1 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t3 131.389
R13663 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n16 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n1 131.388
R13664 SUNSAR_SAR8B_CV_0.XA20.XA2.MP3.D SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n16 71.1534
R13665 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n14 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t1 63.8431
R13666 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n14 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t2 63.8431
R13667 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n0 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t4 63.8431
R13668 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n0 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t0 63.8431
R13669 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n13 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP0.G 22.9652
R13670 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n1 SUNSAR_SAR8B_CV_0.XA20.XA2.MN6.D 20.3299
R13671 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n2 SUNSAR_SAR8B_CV_0.XA20.XA3.MP6.G 20.3299
R13672 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n2 20.3299
R13673 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n3 SUNSAR_SAR8B_CV_0.XA20.XA3.MP5.G 20.3299
R13674 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n4 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n3 20.3299
R13675 SUNSAR_SAR8B_CV_0.XA20.XA3.MP4.G SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n4 20.3299
R13676 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n9 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n6 20.3299
R13677 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n6 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN3.G 20.3299
R13678 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n7 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP3.G 20.3299
R13679 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n8 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n5 20.3299
R13680 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n8 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n7 20.3299
R13681 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n8 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP2.G 20.3299
R13682 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n9 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN2.G 20.3299
R13683 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n11 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN0.G 20.3299
R13684 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n11 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n10 20.3299
R13685 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n10 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n9 20.3299
R13686 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n10 SUNSAR_SAR8B_CV_0.XA20.XA3a.MN1.G 20.3299
R13687 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n5 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP1.G 20.3299
R13688 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n12 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n5 20.3299
R13689 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP0.G SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n12 20.3299
R13690 SUNSAR_SAR8B_CV_0.XA20.XA2.MP5.D SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n15 20.3299
R13691 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n16 SUNSAR_SAR8B_CV_0.XA20.XA2.MP5.D 17.6946
R13692 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t2 1060.4
R13693 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t4 1060.4
R13694 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t8 1060.4
R13695 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t9 1060.4
R13696 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n1 568.956
R13697 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t3 568.956
R13698 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n3 568.956
R13699 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t7 568.956
R13700 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t5 568.956
R13701 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n6 568.956
R13702 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t6 568.956
R13703 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n0 568.956
R13704 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t0 356.344
R13705 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.t1 131.389
R13706 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n9 128.754
R13707 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA2.XA2.MP0.G 97.8829
R13708 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n1 20.3299
R13709 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA2.XA2.MN3.G 20.3299
R13710 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA2.XA2.MP3.G 20.3299
R13711 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n0 20.3299
R13712 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n2 20.3299
R13713 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA2.XA2.MP2.G 20.3299
R13714 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA2.XA2.MN2.G 20.3299
R13715 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA2.XA2.MN0.G 20.3299
R13716 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n5 20.3299
R13717 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n4 20.3299
R13718 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA2.XA2.MN1.G 20.3299
R13719 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA2.XA2.MP1.G 20.3299
R13720 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n0 20.3299
R13721 SUNSAR_SAR8B_CV_0.XA2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n7 20.3299
R13722 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n8 20.3299
R13723 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.D 20.3299
R13724 SUNSAR_SAR8B_CV_0.D<6>.t10 SUNSAR_SAR8B_CV_0.D<6>.t9 1060.4
R13725 SUNSAR_SAR8B_CV_0.D<6>.t9 SUNSAR_SAR8B_CV_0.D<6> 589.284
R13726 SUNSAR_SAR8B_CV_0.D<6>.n16 SUNSAR_SAR8B_CV_0.D<6>.t10 573.85
R13727 SUNSAR_SAR8B_CV_0.D<6>.n4 SUNSAR_SAR8B_CV_0.D<6>.t8 568.956
R13728 SUNSAR_SAR8B_CV_0.D<6>.n3 SUNSAR_SAR8B_CV_0.D<6>.t11 568.956
R13729 SUNSAR_SAR8B_CV_0.D<6>.n2 SUNSAR_SAR8B_CV_0.D<6>.n1 292.5
R13730 SUNSAR_SAR8B_CV_0.D<6>.n11 SUNSAR_SAR8B_CV_0.D<6>.n10 292.5
R13731 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<6>.n9 112.829
R13732 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<6>.n0 112.829
R13733 SUNSAR_SAR8B_CV_0.D<6>.n12 SUNSAR_SAR8B_CV_0.D<6>.n11 111.059
R13734 SUNSAR_SAR8B_CV_0.D<6>.n24 SUNSAR_SAR8B_CV_0.D<6>.n8 89.224
R13735 SUNSAR_SAR8B_CV_0.D<6>.n1 SUNSAR_SAR8B_CV_0.D<6>.t6 63.8431
R13736 SUNSAR_SAR8B_CV_0.D<6>.n1 SUNSAR_SAR8B_CV_0.D<6>.t4 63.8431
R13737 SUNSAR_SAR8B_CV_0.D<6>.n10 SUNSAR_SAR8B_CV_0.D<6>.t5 63.8431
R13738 SUNSAR_SAR8B_CV_0.D<6>.n10 SUNSAR_SAR8B_CV_0.D<6>.t7 63.8431
R13739 SUNSAR_SAR8B_CV_0.D<6>.n13 SUNSAR_SAR8B_CV_0.D<6>.n12 48.7856
R13740 SUNSAR_SAR8B_CV_0.D<6>.n9 SUNSAR_SAR8B_CV_0.D<6>.t1 38.8894
R13741 SUNSAR_SAR8B_CV_0.D<6>.n9 SUNSAR_SAR8B_CV_0.D<6>.t0 38.8894
R13742 SUNSAR_SAR8B_CV_0.D<6>.n0 SUNSAR_SAR8B_CV_0.D<6>.t3 38.8894
R13743 SUNSAR_SAR8B_CV_0.D<6>.n0 SUNSAR_SAR8B_CV_0.D<6>.t2 38.8894
R13744 SUNSAR_SAR8B_CV_0.D<6>.n20 SUNSAR_SAR8B_CV_0.D<6>.n19 35.5626
R13745 SUNSAR_SAR8B_CV_0.D<6>.n3 SUNSAR_SAR8B_CV_0.D<6> 20.3299
R13746 SUNSAR_SAR8B_CV_0.D<6>.n4 SUNSAR_SAR8B_CV_0.D<6>.n3 20.3299
R13747 SUNSAR_SAR8B_CV_0.D<6>.n11 SUNSAR_SAR8B_CV_0.D<6> 20.3299
R13748 SUNSAR_SAR8B_CV_0.D<6>.n19 SUNSAR_SAR8B_CV_0.D<6> 20.2398
R13749 SUNSAR_SAR8B_CV_0.D<6>.n24 SUNSAR_SAR8B_CV_0.D<6>.n23 17.9961
R13750 SUNSAR_SAR8B_CV_0.D<6>.n12 SUNSAR_SAR8B_CV_0.D<6> 17.6946
R13751 SUNSAR_SAR8B_CV_0.D<6>.n18 SUNSAR_SAR8B_CV_0.D<6>.n17 16.9626
R13752 SUNSAR_SAR8B_CV_0.D<6>.n5 SUNSAR_SAR8B_CV_0.D<6> 15.2303
R13753 SUNSAR_SAR8B_CV_0.D<6>.n6 SUNSAR_SAR8B_CV_0.D<6> 13.5534
R13754 SUNSAR_SAR8B_CV_0.D<6>.n16 SUNSAR_SAR8B_CV_0.D<6> 12.939
R13755 SUNSAR_SAR8B_CV_0.D<6>.n8 SUNSAR_SAR8B_CV_0.D<6>.n2 12.8005
R13756 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<6>.n24 11.2946
R13757 SUNSAR_SAR8B_CV_0.D<6>.n7 SUNSAR_SAR8B_CV_0.D<6>.n5 11.2842
R13758 SUNSAR_SAR8B_CV_0.D<6>.n17 SUNSAR_SAR8B_CV_0.D<6>.n16 10.501
R13759 SUNSAR_SAR8B_CV_0.D<6>.n8 SUNSAR_SAR8B_CV_0.D<6>.n7 9.49168
R13760 SUNSAR_SAR8B_CV_0.D<6>.n7 SUNSAR_SAR8B_CV_0.D<6>.n6 9.3005
R13761 SUNSAR_SAR8B_CV_0.D<6>.n14 SUNSAR_SAR8B_CV_0.D<6>.n13 9.3005
R13762 SUNSAR_SAR8B_CV_0.D<6>.n24 SUNSAR_SAR8B_CV_0.D<6>.n13 8.11757
R13763 SUNSAR_SAR8B_CV_0.D<6>.n6 SUNSAR_SAR8B_CV_0.D<6>.n2 6.77697
R13764 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<6>.n20 5.55039
R13765 SUNSAR_SAR8B_CV_0.D<6>.n15 SUNSAR_SAR8B_CV_0.D<6>.n14 4.5005
R13766 SUNSAR_SAR8B_CV_0.D<6>.n23 SUNSAR_SAR8B_CV_0.D<6>.n22 4.5005
R13767 SUNSAR_SAR8B_CV_0.D<6>.n5 SUNSAR_SAR8B_CV_0.D<6>.n4 3.90429
R13768 SUNSAR_SAR8B_CV_0.D<6>.n18 SUNSAR_SAR8B_CV_0.D<6>.n15 3.4105
R13769 SUNSAR_SAR8B_CV_0.D<6>.n22 SUNSAR_SAR8B_CV_0.D<6>.n21 3.4105
R13770 SUNSAR_SAR8B_CV_0.D<6>.n22 SUNSAR_SAR8B_CV_0.D<6>.n15 0.191676
R13771 SUNSAR_SAR8B_CV_0.D<6>.n23 SUNSAR_SAR8B_CV_0.D<6>.n14 0.191676
R13772 SUNSAR_SAR8B_CV_0.D<6>.n17 SUNSAR_SAR8B_CV_0.D<6> 0.173294
R13773 SUNSAR_SAR8B_CV_0.D<6>.n19 SUNSAR_SAR8B_CV_0.D<6> 0.168144
R13774 SUNSAR_SAR8B_CV_0.D<6>.n21 SUNSAR_SAR8B_CV_0.D<6>.n18 0.0713406
R13775 SUNSAR_SAR8B_CV_0.D<6>.n21 SUNSAR_SAR8B_CV_0.D<6> 0.0277464
R13776 SUNSAR_SAR8B_CV_0.D<6>.n20 SUNSAR_SAR8B_CV_0.D<6> 0.00726261
R13777 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t9 568.956
R13778 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t8 568.956
R13779 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n3 292.5
R13780 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n9 292.5
R13781 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n12 197.272
R13782 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n2 112.829
R13783 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n6 112.829
R13784 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n4 111.059
R13785 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t6 63.8431
R13786 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t4 63.8431
R13787 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t7 63.8431
R13788 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t5 63.8431
R13789 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n7 59.1064
R13790 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n5 53.4593
R13791 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n8 51.9534
R13792 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t0 38.8894
R13793 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t2 38.8894
R13794 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t3 38.8894
R13795 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.t1 38.8894
R13796 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n1 38.5859
R13797 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 20.3299
R13798 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 20.3299
R13799 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n11 20.3299
R13800 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 20.3299
R13801 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n10 20.3299
R13802 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 17.6946
R13803 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 17.6946
R13804 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 12.325
R13805 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 12.323
R13806 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 10.3476
R13807 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n0 9.29776
R13808 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.168144
R13809 SUNSAR_SAR8B_CV_0.D<2>.t11 SUNSAR_SAR8B_CV_0.D<2>.t10 1060.4
R13810 SUNSAR_SAR8B_CV_0.D<2>.t10 SUNSAR_SAR8B_CV_0.D<2> 589.284
R13811 SUNSAR_SAR8B_CV_0.D<2>.n11 SUNSAR_SAR8B_CV_0.D<2>.t11 573.85
R13812 SUNSAR_SAR8B_CV_0.D<2>.n3 SUNSAR_SAR8B_CV_0.D<2>.t9 568.956
R13813 SUNSAR_SAR8B_CV_0.D<2>.n2 SUNSAR_SAR8B_CV_0.D<2>.t8 568.956
R13814 SUNSAR_SAR8B_CV_0.D<2>.n1 SUNSAR_SAR8B_CV_0.D<2>.n0 292.5
R13815 SUNSAR_SAR8B_CV_0.D<2>.n26 SUNSAR_SAR8B_CV_0.D<2>.n25 292.5
R13816 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<2>.n8 112.829
R13817 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<2>.n23 112.829
R13818 SUNSAR_SAR8B_CV_0.D<2>.n26 SUNSAR_SAR8B_CV_0.D<2>.n24 111.059
R13819 SUNSAR_SAR8B_CV_0.D<2>.n9 SUNSAR_SAR8B_CV_0.D<2>.n7 89.224
R13820 SUNSAR_SAR8B_CV_0.D<2>.n25 SUNSAR_SAR8B_CV_0.D<2>.t7 63.8431
R13821 SUNSAR_SAR8B_CV_0.D<2>.n25 SUNSAR_SAR8B_CV_0.D<2>.t5 63.8431
R13822 SUNSAR_SAR8B_CV_0.D<2>.n0 SUNSAR_SAR8B_CV_0.D<2>.t6 63.8431
R13823 SUNSAR_SAR8B_CV_0.D<2>.n0 SUNSAR_SAR8B_CV_0.D<2>.t4 63.8431
R13824 SUNSAR_SAR8B_CV_0.D<2>.n24 SUNSAR_SAR8B_CV_0.D<2>.n22 48.7856
R13825 SUNSAR_SAR8B_CV_0.D<2>.n8 SUNSAR_SAR8B_CV_0.D<2>.t1 38.8894
R13826 SUNSAR_SAR8B_CV_0.D<2>.n8 SUNSAR_SAR8B_CV_0.D<2>.t2 38.8894
R13827 SUNSAR_SAR8B_CV_0.D<2>.n23 SUNSAR_SAR8B_CV_0.D<2>.t0 38.8894
R13828 SUNSAR_SAR8B_CV_0.D<2>.n23 SUNSAR_SAR8B_CV_0.D<2>.t3 38.8894
R13829 SUNSAR_SAR8B_CV_0.D<2>.n17 SUNSAR_SAR8B_CV_0.D<2>.n16 31.1545
R13830 SUNSAR_SAR8B_CV_0.D<2>.n16 SUNSAR_SAR8B_CV_0.D<2> 22.3133
R13831 SUNSAR_SAR8B_CV_0.D<2>.n2 SUNSAR_SAR8B_CV_0.D<2> 20.3299
R13832 SUNSAR_SAR8B_CV_0.D<2>.n3 SUNSAR_SAR8B_CV_0.D<2>.n2 20.3299
R13833 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<2>.n26 20.3299
R13834 SUNSAR_SAR8B_CV_0.D<2>.n20 SUNSAR_SAR8B_CV_0.D<2>.n9 17.9961
R13835 SUNSAR_SAR8B_CV_0.D<2>.n24 SUNSAR_SAR8B_CV_0.D<2> 17.6946
R13836 SUNSAR_SAR8B_CV_0.D<2>.n15 SUNSAR_SAR8B_CV_0.D<2>.n14 17.0038
R13837 SUNSAR_SAR8B_CV_0.D<2>.n4 SUNSAR_SAR8B_CV_0.D<2> 15.2303
R13838 SUNSAR_SAR8B_CV_0.D<2>.n5 SUNSAR_SAR8B_CV_0.D<2> 13.5534
R13839 SUNSAR_SAR8B_CV_0.D<2>.n11 SUNSAR_SAR8B_CV_0.D<2> 12.939
R13840 SUNSAR_SAR8B_CV_0.D<2>.n7 SUNSAR_SAR8B_CV_0.D<2>.n1 12.8005
R13841 SUNSAR_SAR8B_CV_0.D<2>.n9 SUNSAR_SAR8B_CV_0.D<2> 11.2946
R13842 SUNSAR_SAR8B_CV_0.D<2>.n6 SUNSAR_SAR8B_CV_0.D<2>.n4 11.2842
R13843 SUNSAR_SAR8B_CV_0.D<2>.n12 SUNSAR_SAR8B_CV_0.D<2>.n11 10.4477
R13844 SUNSAR_SAR8B_CV_0.D<2>.n7 SUNSAR_SAR8B_CV_0.D<2>.n6 9.49168
R13845 SUNSAR_SAR8B_CV_0.D<2>.n6 SUNSAR_SAR8B_CV_0.D<2>.n5 9.3005
R13846 SUNSAR_SAR8B_CV_0.D<2>.n22 SUNSAR_SAR8B_CV_0.D<2>.n21 9.3005
R13847 SUNSAR_SAR8B_CV_0.D<2>.n22 SUNSAR_SAR8B_CV_0.D<2>.n9 8.11757
R13848 SUNSAR_SAR8B_CV_0.D<2>.n5 SUNSAR_SAR8B_CV_0.D<2>.n1 6.77697
R13849 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<2>.n17 5.03616
R13850 SUNSAR_SAR8B_CV_0.D<2>.n21 SUNSAR_SAR8B_CV_0.D<2>.n10 4.5005
R13851 SUNSAR_SAR8B_CV_0.D<2>.n20 SUNSAR_SAR8B_CV_0.D<2>.n19 4.5005
R13852 SUNSAR_SAR8B_CV_0.D<2>.n4 SUNSAR_SAR8B_CV_0.D<2>.n3 3.90429
R13853 SUNSAR_SAR8B_CV_0.D<2>.n15 SUNSAR_SAR8B_CV_0.D<2>.n10 3.4105
R13854 SUNSAR_SAR8B_CV_0.D<2>.n19 SUNSAR_SAR8B_CV_0.D<2>.n18 3.4105
R13855 SUNSAR_SAR8B_CV_0.D<2>.n12 SUNSAR_SAR8B_CV_0.D<2> 0.312734
R13856 SUNSAR_SAR8B_CV_0.D<2>.n19 SUNSAR_SAR8B_CV_0.D<2>.n10 0.191676
R13857 SUNSAR_SAR8B_CV_0.D<2>.n21 SUNSAR_SAR8B_CV_0.D<2>.n20 0.191676
R13858 SUNSAR_SAR8B_CV_0.D<2>.n16 SUNSAR_SAR8B_CV_0.D<2> 0.168144
R13859 SUNSAR_SAR8B_CV_0.D<2>.n13 SUNSAR_SAR8B_CV_0.D<2> 0.103441
R13860 SUNSAR_SAR8B_CV_0.D<2>.n13 SUNSAR_SAR8B_CV_0.D<2> 0.0848373
R13861 SUNSAR_SAR8B_CV_0.D<2>.n18 SUNSAR_SAR8B_CV_0.D<2>.n15 0.0713406
R13862 SUNSAR_SAR8B_CV_0.D<2>.n14 SUNSAR_SAR8B_CV_0.D<2>.n13 0.0577289
R13863 SUNSAR_SAR8B_CV_0.D<2>.n18 SUNSAR_SAR8B_CV_0.D<2> 0.0277464
R13864 SUNSAR_SAR8B_CV_0.D<2>.n14 SUNSAR_SAR8B_CV_0.D<2>.n12 0.0215843
R13865 SUNSAR_SAR8B_CV_0.D<2>.n17 SUNSAR_SAR8B_CV_0.D<2> 0.00726261
R13866 SUNSAR_SAR8B_CV_0.XA4.CN1.t13 SUNSAR_SAR8B_CV_0.XA4.CN1.t8 1060.4
R13867 SUNSAR_SAR8B_CV_0.XA4.CN1.t14 SUNSAR_SAR8B_CV_0.XA4.CN1.t9 1060.4
R13868 SUNSAR_SAR8B_CV_0.XA4.CN1.t11 SUNSAR_SAR8B_CV_0.XA4.CN1.t15 1060.4
R13869 SUNSAR_SAR8B_CV_0.XA4.CN1.t12 SUNSAR_SAR8B_CV_0.XA4.CN1.t10 1060.4
R13870 SUNSAR_SAR8B_CV_0.XA4.CN1.t8 SUNSAR_SAR8B_CV_0.XA4.CN1.n3 568.956
R13871 SUNSAR_SAR8B_CV_0.XA4.CN1.n4 SUNSAR_SAR8B_CV_0.XA4.CN1.t13 568.956
R13872 SUNSAR_SAR8B_CV_0.XA4.CN1.t9 SUNSAR_SAR8B_CV_0.XA4.CN1.n5 568.956
R13873 SUNSAR_SAR8B_CV_0.XA4.CN1.n6 SUNSAR_SAR8B_CV_0.XA4.CN1.t14 568.956
R13874 SUNSAR_SAR8B_CV_0.XA4.CN1.n9 SUNSAR_SAR8B_CV_0.XA4.CN1.t11 568.956
R13875 SUNSAR_SAR8B_CV_0.XA4.CN1.t15 SUNSAR_SAR8B_CV_0.XA4.CN1.n8 568.956
R13876 SUNSAR_SAR8B_CV_0.XA4.CN1.n7 SUNSAR_SAR8B_CV_0.XA4.CN1.t12 568.956
R13877 SUNSAR_SAR8B_CV_0.XA4.CN1.t10 SUNSAR_SAR8B_CV_0.XA4.CN1.n2 568.956
R13878 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.CN1.n1 312.829
R13879 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.CN1.n0 312.829
R13880 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.CN1.n12 184.471
R13881 SUNSAR_SAR8B_CV_0.XA4.CN1.n14 SUNSAR_SAR8B_CV_0.XA4.CN1.n13 92.5005
R13882 SUNSAR_SAR8B_CV_0.XA4.CN1.n17 SUNSAR_SAR8B_CV_0.XA4.CN1.n16 92.5005
R13883 SUNSAR_SAR8B_CV_0.XA4.CN1.n15 SUNSAR_SAR8B_CV_0.XA4.CN1 90.7299
R13884 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.CN1.n18 90.7299
R13885 SUNSAR_SAR8B_CV_0.XA4.CN1.n1 SUNSAR_SAR8B_CV_0.XA4.CN1.t5 63.8431
R13886 SUNSAR_SAR8B_CV_0.XA4.CN1.n1 SUNSAR_SAR8B_CV_0.XA4.CN1.t6 63.8431
R13887 SUNSAR_SAR8B_CV_0.XA4.CN1.n0 SUNSAR_SAR8B_CV_0.XA4.CN1.t2 63.8431
R13888 SUNSAR_SAR8B_CV_0.XA4.CN1.n0 SUNSAR_SAR8B_CV_0.XA4.CN1.t0 63.8431
R13889 SUNSAR_SAR8B_CV_0.XA4.CN1.n18 SUNSAR_SAR8B_CV_0.XA4.CN1.n15 53.4593
R13890 SUNSAR_SAR8B_CV_0.XA4.CN1.n16 SUNSAR_SAR8B_CV_0.XA4.CN1.t4 38.8894
R13891 SUNSAR_SAR8B_CV_0.XA4.CN1.n16 SUNSAR_SAR8B_CV_0.XA4.CN1.t7 38.8894
R13892 SUNSAR_SAR8B_CV_0.XA4.CN1.n13 SUNSAR_SAR8B_CV_0.XA4.CN1.t1 38.8894
R13893 SUNSAR_SAR8B_CV_0.XA4.CN1.n13 SUNSAR_SAR8B_CV_0.XA4.CN1.t3 38.8894
R13894 SUNSAR_SAR8B_CV_0.XA4.CN1.n15 SUNSAR_SAR8B_CV_0.XA4.CN1.n14 38.024
R13895 SUNSAR_SAR8B_CV_0.XA4.CN1.n18 SUNSAR_SAR8B_CV_0.XA4.CN1.n17 38.024
R13896 SUNSAR_SAR8B_CV_0.XA4.CN1.n6 SUNSAR_SAR8B_CV_0.XA4.CN1.n3 20.3299
R13897 SUNSAR_SAR8B_CV_0.XA4.CN1.n3 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13898 SUNSAR_SAR8B_CV_0.XA4.CN1.n4 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13899 SUNSAR_SAR8B_CV_0.XA4.CN1.n5 SUNSAR_SAR8B_CV_0.XA4.CN1.n2 20.3299
R13900 SUNSAR_SAR8B_CV_0.XA4.CN1.n5 SUNSAR_SAR8B_CV_0.XA4.CN1.n4 20.3299
R13901 SUNSAR_SAR8B_CV_0.XA4.CN1.n5 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13902 SUNSAR_SAR8B_CV_0.XA4.CN1.n6 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13903 SUNSAR_SAR8B_CV_0.XA4.CN1.n8 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13904 SUNSAR_SAR8B_CV_0.XA4.CN1.n8 SUNSAR_SAR8B_CV_0.XA4.CN1.n7 20.3299
R13905 SUNSAR_SAR8B_CV_0.XA4.CN1.n7 SUNSAR_SAR8B_CV_0.XA4.CN1.n6 20.3299
R13906 SUNSAR_SAR8B_CV_0.XA4.CN1.n7 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13907 SUNSAR_SAR8B_CV_0.XA4.CN1.n2 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13908 SUNSAR_SAR8B_CV_0.XA4.CN1.n9 SUNSAR_SAR8B_CV_0.XA4.CN1.n2 20.3299
R13909 SUNSAR_SAR8B_CV_0.XA4.CN1.n14 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13910 SUNSAR_SAR8B_CV_0.XA4.CN1.n17 SUNSAR_SAR8B_CV_0.XA4.CN1 20.3299
R13911 SUNSAR_SAR8B_CV_0.XA4.CN1.n10 SUNSAR_SAR8B_CV_0.XA4.CN1 13.5534
R13912 SUNSAR_SAR8B_CV_0.XA4.CN1.n12 SUNSAR_SAR8B_CV_0.XA4.CN1.n9 12.8005
R13913 SUNSAR_SAR8B_CV_0.XA4.CN1.n12 SUNSAR_SAR8B_CV_0.XA4.CN1.n11 9.39466
R13914 SUNSAR_SAR8B_CV_0.XA4.CN1.n11 SUNSAR_SAR8B_CV_0.XA4.CN1.n10 9.39462
R13915 SUNSAR_SAR8B_CV_0.XA4.CN1.n10 SUNSAR_SAR8B_CV_0.XA4.CN1.n9 6.77697
R13916 SUNSAR_SAR8B_CV_0.XA4.CN1.n11 SUNSAR_SAR8B_CV_0.XA4.CN1 3.95537
R13917 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t3 1060.4
R13918 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t9 1060.4
R13919 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t2 1060.4
R13920 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t4 1060.4
R13921 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n2 568.956
R13922 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t8 568.956
R13923 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n4 568.956
R13924 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t6 568.956
R13925 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t7 568.956
R13926 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n7 568.956
R13927 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t5 568.956
R13928 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n1 568.956
R13929 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t0 356.344
R13930 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.D SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.t1 151.719
R13931 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.D 128.754
R13932 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n8 97.8829
R13933 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n2 20.3299
R13934 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA3.XA2.MN3.G 20.3299
R13935 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA3.XA2.MP3.G 20.3299
R13936 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n1 20.3299
R13937 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n3 20.3299
R13938 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA3.XA2.MP2.G 20.3299
R13939 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA3.XA2.MN2.G 20.3299
R13940 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA3.XA2.MN0.G 20.3299
R13941 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n6 20.3299
R13942 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n5 20.3299
R13943 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA3.XA2.MN1.G 20.3299
R13944 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA3.XA2.MP1.G 20.3299
R13945 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n1 20.3299
R13946 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA3.XA2.MP0.G 20.3299
R13947 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n0 20.3299
R13948 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t9 568.956
R13949 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t8 568.956
R13950 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n0 312.829
R13951 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n5 292.5
R13952 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 197.272
R13953 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n8 92.5005
R13954 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n11 92.5005
R13955 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n13 90.7299
R13956 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t5 63.8431
R13957 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t7 63.8431
R13958 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t6 63.8431
R13959 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t4 63.8431
R13960 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n7 59.1064
R13961 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n10 53.4593
R13962 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t2 38.8894
R13963 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t1 38.8894
R13964 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t3 38.8894
R13965 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.t0 38.8894
R13966 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n9 38.024
R13967 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n13 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n12 38.024
R13968 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n2 32.2698
R13969 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 31.624
R13970 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 20.3299
R13971 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n3 20.3299
R13972 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n4 20.3299
R13973 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n6 20.3299
R13974 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 20.3299
R13975 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 20.3299
R13976 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 12.325
R13977 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 12.323
R13978 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 10.3476
R13979 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n1 9.64335
R13980 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.168144
R13981 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t4 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t8 1060.4
R13982 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t3 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t7 1060.4
R13983 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t5 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t6 1060.4
R13984 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t8 SUNSAR_SAR8B_CV_0.XA20.XA9.MP0.G 589.284
R13985 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t7 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.G 589.284
R13986 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t6 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.G 589.284
R13987 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n2 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t3 574.383
R13988 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n3 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t5 574.383
R13989 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n7 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t4 568.956
R13990 SUNSAR_SAR8B_CV_0.XA20.XA10.MP0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n0 312.829
R13991 SUNSAR_SAR8B_CV_0.XA20.XA10.MP0.D SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n11 142.306
R13992 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n1 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t1 131.389
R13993 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n0 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t0 63.8431
R13994 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n0 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.t2 63.8431
R13995 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n8 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n7 16.077
R13996 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n4 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n2 15.0655
R13997 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n7 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n6 12.8005
R13998 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n9 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n1 12.8005
R13999 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n2 SUNSAR_SAR8B_CV_0.XA20.XA1.MN0.G 10.633
R14000 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n3 SUNSAR_SAR8B_CV_0.XA20.XA4.MN0.G 10.633
R14001 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n11 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n10 9.49168
R14002 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n6 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n5 9.3005
R14003 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n10 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n9 9.3005
R14004 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n6 SUNSAR_SAR8B_CV_0.XA20.XA9.MN0.G 7.52991
R14005 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n9 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.D 7.52991
R14006 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n11 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n1 6.77697
R14007 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n4 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n3 4.19047
R14008 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n5 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n4 2.71006
R14009 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n10 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n8 1.61079
R14010 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n8 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n5 0.191676
R14011 SUNSAR_SAR8B_CV_0.XA1.ENO.t2 SUNSAR_SAR8B_CV_0.XA1.ENO.t8 1060.4
R14012 SUNSAR_SAR8B_CV_0.XA1.ENO.t7 SUNSAR_SAR8B_CV_0.XA1.ENO.t6 1060.4
R14013 SUNSAR_SAR8B_CV_0.XA1.ENO.t8 SUNSAR_SAR8B_CV_0.XA2.EN 589.284
R14014 SUNSAR_SAR8B_CV_0.XA1.ENO.t6 SUNSAR_SAR8B_CV_0.XA2.EN 589.284
R14015 SUNSAR_SAR8B_CV_0.XA1.ENO.n0 SUNSAR_SAR8B_CV_0.XA1.ENO.t2 583.638
R14016 SUNSAR_SAR8B_CV_0.XA1.ENO.n5 SUNSAR_SAR8B_CV_0.XA1.ENO.t5 574.383
R14017 SUNSAR_SAR8B_CV_0.XA1.ENO.n6 SUNSAR_SAR8B_CV_0.XA1.ENO.t3 574.383
R14018 SUNSAR_SAR8B_CV_0.XA1.ENO.n12 SUNSAR_SAR8B_CV_0.XA1.ENO.t7 572.893
R14019 SUNSAR_SAR8B_CV_0.XA1.ENO.n10 SUNSAR_SAR8B_CV_0.XA1.ENO.t4 568.956
R14020 SUNSAR_SAR8B_CV_0.XA1.ENO.n2 SUNSAR_SAR8B_CV_0.XA1.ENO.t1 356.344
R14021 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.ENO.n17 268.8
R14022 SUNSAR_SAR8B_CV_0.XA1.ENO.n1 SUNSAR_SAR8B_CV_0.XA1.ENO.t0 131.389
R14023 SUNSAR_SAR8B_CV_0.XA1.ENO.n1 SUNSAR_SAR8B_CV_0.XA1.ENO.n0 90.7299
R14024 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.ENO.n1 20.3299
R14025 SUNSAR_SAR8B_CV_0.XA1.ENO.n13 SUNSAR_SAR8B_CV_0.XA1.ENO.n12 20.0513
R14026 SUNSAR_SAR8B_CV_0.XA1.ENO.n11 SUNSAR_SAR8B_CV_0.XA1.ENO.n10 16.1445
R14027 SUNSAR_SAR8B_CV_0.XA1.ENO.n12 SUNSAR_SAR8B_CV_0.XA2.EN 15.1965
R14028 SUNSAR_SAR8B_CV_0.XA1.ENO.n3 SUNSAR_SAR8B_CV_0.XA2.EN 13.5534
R14029 SUNSAR_SAR8B_CV_0.XA1.ENO.n10 SUNSAR_SAR8B_CV_0.XA1.ENO.n9 12.8005
R14030 SUNSAR_SAR8B_CV_0.XA1.ENO.n17 SUNSAR_SAR8B_CV_0.XA1.ENO.n2 12.8005
R14031 SUNSAR_SAR8B_CV_0.XA1.ENO.n5 SUNSAR_SAR8B_CV_0.XA2.EN 10.633
R14032 SUNSAR_SAR8B_CV_0.XA1.ENO.n6 SUNSAR_SAR8B_CV_0.XA2.EN 10.633
R14033 SUNSAR_SAR8B_CV_0.XA1.ENO.n17 SUNSAR_SAR8B_CV_0.XA1.ENO.n16 9.35932
R14034 SUNSAR_SAR8B_CV_0.XA1.ENO.n9 SUNSAR_SAR8B_CV_0.XA1.ENO.n8 9.3005
R14035 SUNSAR_SAR8B_CV_0.XA1.ENO.n4 SUNSAR_SAR8B_CV_0.XA1.ENO.n3 9.3005
R14036 SUNSAR_SAR8B_CV_0.XA1.ENO.n9 SUNSAR_SAR8B_CV_0.XA2.EN 7.52991
R14037 SUNSAR_SAR8B_CV_0.XA1.ENO.n3 SUNSAR_SAR8B_CV_0.XA1.ENO.n2 6.77697
R14038 SUNSAR_SAR8B_CV_0.XA1.ENO.n0 SUNSAR_SAR8B_CV_0.XA2.EN 5.64756
R14039 SUNSAR_SAR8B_CV_0.XA1.ENO.n7 SUNSAR_SAR8B_CV_0.XA1.ENO.n5 5.35958
R14040 SUNSAR_SAR8B_CV_0.XA1.ENO.n14 SUNSAR_SAR8B_CV_0.XA1.ENO.n13 4.5005
R14041 SUNSAR_SAR8B_CV_0.XA1.ENO.n16 SUNSAR_SAR8B_CV_0.XA1.ENO.n15 4.5005
R14042 SUNSAR_SAR8B_CV_0.XA1.ENO.n15 SUNSAR_SAR8B_CV_0.XA2.EN 4.33874
R14043 SUNSAR_SAR8B_CV_0.XA1.ENO.n7 SUNSAR_SAR8B_CV_0.XA1.ENO.n6 4.19047
R14044 SUNSAR_SAR8B_CV_0.XA1.ENO.n8 SUNSAR_SAR8B_CV_0.XA1.ENO.n7 4.00418
R14045 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.ENO.n11 2.35274
R14046 SUNSAR_SAR8B_CV_0.XA1.ENO.n15 SUNSAR_SAR8B_CV_0.XA1.ENO.n14 0.191676
R14047 SUNSAR_SAR8B_CV_0.XA1.ENO.n16 SUNSAR_SAR8B_CV_0.XA1.ENO.n4 0.132853
R14048 SUNSAR_SAR8B_CV_0.XA1.ENO.n11 SUNSAR_SAR8B_CV_0.XA1.ENO.n8 0.123303
R14049 SUNSAR_SAR8B_CV_0.XA1.ENO.n14 SUNSAR_SAR8B_CV_0.XA2.EN 0.0740294
R14050 SUNSAR_SAR8B_CV_0.XA1.ENO.n13 SUNSAR_SAR8B_CV_0.XA1.ENO.n4 0.0593235
R14051 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t6 1060.4
R14052 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t2 1060.4
R14053 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t5 1060.4
R14054 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t7 1060.4
R14055 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n1 568.956
R14056 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t4 568.956
R14057 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n3 568.956
R14058 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t9 568.956
R14059 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t8 568.956
R14060 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n6 568.956
R14061 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t3 568.956
R14062 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n0 568.956
R14063 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t0 356.344
R14064 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.t1 131.389
R14065 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n9 128.754
R14066 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA6.XA2.MP0.G 97.8829
R14067 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n1 20.3299
R14068 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA6.XA2.MN3.G 20.3299
R14069 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA6.XA2.MP3.G 20.3299
R14070 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n0 20.3299
R14071 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n2 20.3299
R14072 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA6.XA2.MP2.G 20.3299
R14073 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA6.XA2.MN2.G 20.3299
R14074 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA6.XA2.MN0.G 20.3299
R14075 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n5 20.3299
R14076 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n4 20.3299
R14077 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA6.XA2.MN1.G 20.3299
R14078 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA6.XA2.MP1.G 20.3299
R14079 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n0 20.3299
R14080 SUNSAR_SAR8B_CV_0.XA6.XA2.MP0.G SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n7 20.3299
R14081 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n8 20.3299
R14082 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.D 20.3299
R14083 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t3 1060.4
R14084 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t9 1060.4
R14085 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t6 1060.4
R14086 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t7 1060.4
R14087 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n3 568.956
R14088 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t2 568.956
R14089 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n5 568.956
R14090 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t5 568.956
R14091 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t8 568.956
R14092 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n8 568.956
R14093 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t4 568.956
R14094 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n2 568.956
R14095 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.D SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t0 376.673
R14096 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.t1 131.389
R14097 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.D 121.977
R14098 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n3 20.3299
R14099 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA6.XA4.MP3.G 20.3299
R14100 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA6.XA4.MN3.G 20.3299
R14101 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n2 20.3299
R14102 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n4 20.3299
R14103 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA6.XA4.MN2.G 20.3299
R14104 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA6.XA4.MP2.G 20.3299
R14105 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA6.XA4.MP0.G 20.3299
R14106 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n7 20.3299
R14107 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n6 20.3299
R14108 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA6.XA4.MP1.G 20.3299
R14109 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA6.XA4.MN1.G 20.3299
R14110 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n2 20.3299
R14111 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n0 12.8005
R14112 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA6.XA4.MN0.G 10.6968
R14113 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n1 9.49168
R14114 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n11 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n10 9.47055
R14115 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n12 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n11 9.3005
R14116 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n12 7.52991
R14117 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n0 6.77697
R14118 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n9 5.36434
R14119 SUNSAR_SAR8B_CV_0.XA5.ENO.t7 SUNSAR_SAR8B_CV_0.XA5.ENO.t6 1060.4
R14120 SUNSAR_SAR8B_CV_0.XA5.ENO.t2 SUNSAR_SAR8B_CV_0.XA5.ENO.t4 1060.4
R14121 SUNSAR_SAR8B_CV_0.XA5.ENO.t6 SUNSAR_SAR8B_CV_0.XA6.EN 589.284
R14122 SUNSAR_SAR8B_CV_0.XA5.ENO.t4 SUNSAR_SAR8B_CV_0.XA6.EN 589.284
R14123 SUNSAR_SAR8B_CV_0.XA5.ENO.n1 SUNSAR_SAR8B_CV_0.XA5.ENO.t2 583.638
R14124 SUNSAR_SAR8B_CV_0.XA5.ENO.n6 SUNSAR_SAR8B_CV_0.XA5.ENO.t3 574.383
R14125 SUNSAR_SAR8B_CV_0.XA5.ENO.n7 SUNSAR_SAR8B_CV_0.XA5.ENO.t8 574.383
R14126 SUNSAR_SAR8B_CV_0.XA5.ENO.n5 SUNSAR_SAR8B_CV_0.XA5.ENO.t7 572.893
R14127 SUNSAR_SAR8B_CV_0.XA5.ENO.n11 SUNSAR_SAR8B_CV_0.XA5.ENO.t5 568.956
R14128 SUNSAR_SAR8B_CV_0.XA5.ENO.n0 SUNSAR_SAR8B_CV_0.XA5.ENO.t0 356.344
R14129 SUNSAR_SAR8B_CV_0.XA5.ENO.n3 SUNSAR_SAR8B_CV_0.XA6.EN 268.8
R14130 SUNSAR_SAR8B_CV_0.XA5.ENO.n2 SUNSAR_SAR8B_CV_0.XA5.ENO.t1 131.389
R14131 SUNSAR_SAR8B_CV_0.XA5.ENO.n2 SUNSAR_SAR8B_CV_0.XA5.ENO.n1 90.7299
R14132 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.ENO.n2 20.3299
R14133 SUNSAR_SAR8B_CV_0.XA5.ENO.n15 SUNSAR_SAR8B_CV_0.XA5.ENO.n5 20.0513
R14134 SUNSAR_SAR8B_CV_0.XA5.ENO.n12 SUNSAR_SAR8B_CV_0.XA5.ENO.n11 16.1445
R14135 SUNSAR_SAR8B_CV_0.XA5.ENO.n5 SUNSAR_SAR8B_CV_0.XA6.EN 15.1965
R14136 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.ENO.n17 13.5534
R14137 SUNSAR_SAR8B_CV_0.XA5.ENO.n11 SUNSAR_SAR8B_CV_0.XA5.ENO.n10 12.8005
R14138 SUNSAR_SAR8B_CV_0.XA5.ENO.n3 SUNSAR_SAR8B_CV_0.XA5.ENO.n0 12.8005
R14139 SUNSAR_SAR8B_CV_0.XA5.ENO.n6 SUNSAR_SAR8B_CV_0.XA6.EN 10.633
R14140 SUNSAR_SAR8B_CV_0.XA5.ENO.n7 SUNSAR_SAR8B_CV_0.XA6.EN 10.633
R14141 SUNSAR_SAR8B_CV_0.XA5.ENO.n4 SUNSAR_SAR8B_CV_0.XA5.ENO.n3 9.35932
R14142 SUNSAR_SAR8B_CV_0.XA5.ENO.n10 SUNSAR_SAR8B_CV_0.XA5.ENO.n9 9.3005
R14143 SUNSAR_SAR8B_CV_0.XA5.ENO.n17 SUNSAR_SAR8B_CV_0.XA5.ENO.n16 9.3005
R14144 SUNSAR_SAR8B_CV_0.XA5.ENO.n10 SUNSAR_SAR8B_CV_0.XA6.EN 7.52991
R14145 SUNSAR_SAR8B_CV_0.XA5.ENO.n17 SUNSAR_SAR8B_CV_0.XA5.ENO.n0 6.77697
R14146 SUNSAR_SAR8B_CV_0.XA5.ENO.n1 SUNSAR_SAR8B_CV_0.XA6.EN 5.64756
R14147 SUNSAR_SAR8B_CV_0.XA5.ENO.n8 SUNSAR_SAR8B_CV_0.XA5.ENO.n6 5.35958
R14148 SUNSAR_SAR8B_CV_0.XA5.ENO.n15 SUNSAR_SAR8B_CV_0.XA5.ENO.n14 4.5005
R14149 SUNSAR_SAR8B_CV_0.XA5.ENO.n13 SUNSAR_SAR8B_CV_0.XA5.ENO.n4 4.5005
R14150 SUNSAR_SAR8B_CV_0.XA5.ENO.n13 SUNSAR_SAR8B_CV_0.XA6.EN 4.33874
R14151 SUNSAR_SAR8B_CV_0.XA5.ENO.n8 SUNSAR_SAR8B_CV_0.XA5.ENO.n7 4.19047
R14152 SUNSAR_SAR8B_CV_0.XA5.ENO.n9 SUNSAR_SAR8B_CV_0.XA5.ENO.n8 4.00418
R14153 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.ENO.n12 2.35274
R14154 SUNSAR_SAR8B_CV_0.XA5.ENO.n14 SUNSAR_SAR8B_CV_0.XA5.ENO.n13 0.191676
R14155 SUNSAR_SAR8B_CV_0.XA5.ENO.n16 SUNSAR_SAR8B_CV_0.XA5.ENO.n4 0.132853
R14156 SUNSAR_SAR8B_CV_0.XA5.ENO.n12 SUNSAR_SAR8B_CV_0.XA5.ENO.n9 0.123303
R14157 SUNSAR_SAR8B_CV_0.XA5.ENO.n14 SUNSAR_SAR8B_CV_0.XA6.EN 0.0740294
R14158 SUNSAR_SAR8B_CV_0.XA5.ENO.n16 SUNSAR_SAR8B_CV_0.XA5.ENO.n15 0.0593235
R14159 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t7 1060.4
R14160 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XC08.XA2.MN0.G 589.284
R14161 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t2 572.893
R14162 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t3 572.893
R14163 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t5 572.893
R14164 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t4 568.956
R14165 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t6 568.956
R14166 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t1 356.344
R14167 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.t0 135.293
R14168 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XC08.XA1.MN0.D 115.954
R14169 SUNSAR_CAPT8B_CV_0.XC08.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n13 85.0829
R14170 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n5 22.1005
R14171 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XC08.XA2.MP0.G 20.3299
R14172 SUNSAR_CAPT8B_CV_0.XC08.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n2 15.2303
R14173 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.G 15.1965
R14174 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.G 15.1965
R14175 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.G 15.1965
R14176 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.G 13.5534
R14177 SUNSAR_CAPT8B_CV_0.XC08.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n12 13.5534
R14178 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n0 12.8005
R14179 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n1 12.6805
R14180 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n3 9.49168
R14181 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n7 9.3005
R14182 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n11 9.3005
R14183 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n4 9.10273
R14184 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n6 6.77697
R14185 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n0 6.77697
R14186 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n9 5.70934
R14187 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n10 3.40124
R14188 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n8 1.79829
R14189 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n5 0.191676
R14190 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t6 1060.4
R14191 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t9 1060.4
R14192 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t3 1060.4
R14193 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t2 1060.4
R14194 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n1 568.956
R14195 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t5 568.956
R14196 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n3 568.956
R14197 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t8 568.956
R14198 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t7 568.956
R14199 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n6 568.956
R14200 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t4 568.956
R14201 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n0 568.956
R14202 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t0 356.344
R14203 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.t1 135.293
R14204 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n10 128.754
R14205 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n1 20.3299
R14206 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA7.XA4.MP3.G 20.3299
R14207 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA7.XA4.MN3.G 20.3299
R14208 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n0 20.3299
R14209 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n2 20.3299
R14210 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA7.XA4.MN2.G 20.3299
R14211 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA7.XA4.MP2.G 20.3299
R14212 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA7.XA4.MP0.G 20.3299
R14213 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n5 20.3299
R14214 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n4 20.3299
R14215 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA7.XA4.MP1.G 20.3299
R14216 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA7.XA4.MN1.G 20.3299
R14217 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n0 20.3299
R14218 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.D 20.3299
R14219 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n8 16.3643
R14220 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n9 15.2303
R14221 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA7.XA4.MN0.G 15.1965
R14222 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n7 3.93805
R14223 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n1 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n0 292.5
R14224 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n3 SUNSAR_SAR8B_CV_0.XB1.XA3.MN1.D 115.954
R14225 SUNSAR_SAR8B_CV_0.XB1.XA3.MN1.D SUNSAR_SAR8B_CV_0.XB1.XA3.B.n2 112.829
R14226 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n20 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n19 80.3272
R14227 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n19 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n15 80.3272
R14228 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n29 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n28 80.3272
R14229 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n28 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n27 80.3272
R14230 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n45 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n44 80.3272
R14231 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n44 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n43 80.3272
R14232 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n61 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n60 80.3272
R14233 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n60 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n59 80.3272
R14234 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n80 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n79 80.3272
R14235 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n79 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n78 80.3272
R14236 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n0 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t2 63.8431
R14237 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n0 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t0 63.8431
R14238 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n2 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t3 38.8894
R14239 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n2 SUNSAR_SAR8B_CV_0.XB1.XA3.B.t1 38.8894
R14240 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n19 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n18 37.6605
R14241 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n31 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n28 37.6605
R14242 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n47 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n44 37.6605
R14243 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n63 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n60 37.6605
R14244 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n79 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n7 37.6605
R14245 SUNSAR_SAR8B_CV_0.XB1.XA3.MP1_DMY.D SUNSAR_SAR8B_CV_0.XB1.XA3.B.n84 13.5534
R14246 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n3 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n1 12.8005
R14247 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n83 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n82 9.93976
R14248 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n83 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n3 9.39659
R14249 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n84 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n83 9.39269
R14250 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n84 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n1 6.77697
R14251 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n22 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n10 1.98907
R14252 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n13 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n10 1.98907
R14253 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n37 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n36 1.98907
R14254 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n36 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n35 1.98907
R14255 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n53 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n52 1.98907
R14256 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n52 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n51 1.98907
R14257 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n69 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n68 1.98907
R14258 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n68 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n67 1.98907
R14259 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n8 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n4 1.98907
R14260 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n76 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n8 1.98907
R14261 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n16 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n10 1.8324
R14262 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n36 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n26 1.8324
R14263 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n52 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n42 1.8324
R14264 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n68 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n58 1.8324
R14265 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n74 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n8 1.8324
R14266 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n21 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n20 1.5005
R14267 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n15 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n14 1.5005
R14268 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n18 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n17 1.5005
R14269 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n29 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n25 1.5005
R14270 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n34 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n27 1.5005
R14271 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n32 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n31 1.5005
R14272 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n45 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n41 1.5005
R14273 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n50 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n43 1.5005
R14274 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n48 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n47 1.5005
R14275 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n61 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n57 1.5005
R14276 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n66 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n59 1.5005
R14277 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n64 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n63 1.5005
R14278 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n78 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n77 1.5005
R14279 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n73 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n7 1.5005
R14280 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n81 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n80 1.5005
R14281 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n14 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n13 1.13717
R14282 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n17 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n16 1.13717
R14283 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n22 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n21 1.13717
R14284 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n35 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n34 1.13717
R14285 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n32 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n26 1.13717
R14286 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n37 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n25 1.13717
R14287 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n51 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n50 1.13717
R14288 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n48 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n42 1.13717
R14289 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n53 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n41 1.13717
R14290 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n67 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n66 1.13717
R14291 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n64 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n58 1.13717
R14292 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n69 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n57 1.13717
R14293 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n77 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n76 1.13717
R14294 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n74 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n73 1.13717
R14295 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n21 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n11 0.754667
R14296 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n20 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n12 0.754667
R14297 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n15 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n12 0.754667
R14298 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n14 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n11 0.754667
R14299 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n33 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n25 0.754667
R14300 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n30 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n29 0.754667
R14301 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n30 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n27 0.754667
R14302 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n34 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n33 0.754667
R14303 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n49 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n41 0.754667
R14304 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n46 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n45 0.754667
R14305 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n46 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n43 0.754667
R14306 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n50 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n49 0.754667
R14307 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n65 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n57 0.754667
R14308 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n62 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n61 0.754667
R14309 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n62 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n59 0.754667
R14310 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n66 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n65 0.754667
R14311 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n77 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n5 0.754667
R14312 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n80 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n6 0.754667
R14313 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n78 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n6 0.754667
R14314 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n81 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n5 0.754667
R14315 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n82 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n81 0.694488
R14316 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n39 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB4.B 0.682
R14317 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB0.B SUNSAR_SAR8B_CV_0.XB1.XA3.B.n71 0.682
R14318 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n55 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n39 0.617029
R14319 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n71 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n55 0.617029
R14320 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n82 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n4 0.369799
R14321 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n18 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n12 0.338
R14322 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n17 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n11 0.338
R14323 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n31 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n30 0.338
R14324 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n33 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n32 0.338
R14325 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n47 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n46 0.338
R14326 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n49 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n48 0.338
R14327 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n63 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n62 0.338
R14328 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n65 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n64 0.338
R14329 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n7 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n6 0.338
R14330 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n73 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n5 0.338
R14331 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n13 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n9 0.284067
R14332 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n35 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n24 0.284067
R14333 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n51 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n40 0.284067
R14334 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n67 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n56 0.284067
R14335 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n76 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n75 0.284067
R14336 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n75 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n72 0.157167
R14337 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n23 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n9 0.157167
R14338 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n38 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n24 0.157167
R14339 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n54 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n40 0.157167
R14340 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n70 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n56 0.157167
R14341 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n16 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n9 0.1274
R14342 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n23 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n22 0.1274
R14343 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n26 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n24 0.1274
R14344 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n38 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n37 0.1274
R14345 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n42 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n40 0.1274
R14346 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n54 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n53 0.1274
R14347 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n58 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n56 0.1274
R14348 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n70 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n69 0.1274
R14349 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n72 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n4 0.1274
R14350 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n75 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n74 0.1274
R14351 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n39 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB3.B 0.0654706
R14352 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n55 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB2.B 0.0654706
R14353 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n71 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB1.B 0.0654706
R14354 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB4.B SUNSAR_SAR8B_CV_0.XB1.XA3.B.n23 0.02165
R14355 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB3.B SUNSAR_SAR8B_CV_0.XB1.XA3.B.n38 0.02165
R14356 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB2.B SUNSAR_SAR8B_CV_0.XB1.XA3.B.n54 0.02165
R14357 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB1.B SUNSAR_SAR8B_CV_0.XB1.XA3.B.n70 0.02165
R14358 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n72 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB0.B 0.02165
R14359 uo_out[5].t2 uo_out[5].t3 1060.4
R14360 uo_out[5].t3 uo_out[5] 589.284
R14361 uo_out[5].n0 uo_out[5].t2 574.383
R14362 uo_out[5].n1 uo_out[5].t1 361.707
R14363 uo_out[5].n3 uo_out[5].t0 131.389
R14364 uo_out[5].n2 uo_out[5] 118.966
R14365 uo_out[5].n6 uo_out[5] 12.3444
R14366 uo_out[5] uo_out[5].n1 10.6968
R14367 uo_out[5].n0 uo_out[5] 10.633
R14368 uo_out[5].n4 uo_out[5] 10.5417
R14369 uo_out[5].n3 uo_out[5].n2 9.78874
R14370 uo_out[5].n4 uo_out[5].n3 9.78874
R14371 uo_out[5].n1 uo_out[5].n0 9.53185
R14372 uo_out[5].n5 uo_out[5].n2 9.39464
R14373 uo_out[5].n5 uo_out[5].n4 9.39464
R14374 uo_out[5].n6 uo_out[5].n5 2.56815
R14375 uo_out[5] uo_out[5].n6 0.180647
R14376 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t9 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t14 1060.4
R14377 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t11 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t13 1060.4
R14378 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t7 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t8 1060.4
R14379 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t16 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t12 1060.4
R14380 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t5 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t6 1060.4
R14381 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t14 SUNSAR_SAR8B_CV_0.XA20.XA2.MN6.G 589.284
R14382 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t10 568.956
R14383 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n2 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t9 568.956
R14384 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n1 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t15 568.956
R14385 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t13 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n6 568.956
R14386 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n7 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t11 568.956
R14387 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t8 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n8 568.956
R14388 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n9 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t7 568.956
R14389 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n12 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t16 568.956
R14390 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t12 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n11 568.956
R14391 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n10 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t5 568.956
R14392 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t6 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n5 568.956
R14393 SUNSAR_SAR8B_CV_0.XA20.XA3.MP5.D SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n17 312.829
R14394 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n15 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n0 297.865
R14395 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n16 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t4 131.389
R14396 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n18 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n16 131.388
R14397 SUNSAR_SAR8B_CV_0.XA20.XA3.MP3.D SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n18 71.1534
R14398 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n17 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t2 63.8431
R14399 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n17 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t3 63.8431
R14400 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n0 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t1 63.8431
R14401 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n0 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t0 63.8431
R14402 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n2 SUNSAR_SAR8B_CV_0.XA20.XA2.MP6.G 20.3299
R14403 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n1 SUNSAR_SAR8B_CV_0.XA20.XA2.MP4.G 20.3299
R14404 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n1 20.3299
R14405 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n3 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n2 20.3299
R14406 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n9 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n6 20.3299
R14407 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n6 SUNSAR_SAR8B_CV_0.XA20.XA2a.MN3.G 20.3299
R14408 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n7 SUNSAR_SAR8B_CV_0.XA20.XA2a.MP3.G 20.3299
R14409 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n8 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n5 20.3299
R14410 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n8 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n7 20.3299
R14411 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n8 SUNSAR_SAR8B_CV_0.XA20.XA2a.MP2.G 20.3299
R14412 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n9 SUNSAR_SAR8B_CV_0.XA20.XA2a.MN2.G 20.3299
R14413 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n11 SUNSAR_SAR8B_CV_0.XA20.XA2a.MN0.G 20.3299
R14414 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n11 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n10 20.3299
R14415 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n10 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n9 20.3299
R14416 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n10 SUNSAR_SAR8B_CV_0.XA20.XA2a.MN1.G 20.3299
R14417 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n5 SUNSAR_SAR8B_CV_0.XA20.XA2a.MP1.G 20.3299
R14418 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n12 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n5 20.3299
R14419 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n16 SUNSAR_SAR8B_CV_0.XA20.XA3.MN6.D 20.3299
R14420 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n18 SUNSAR_SAR8B_CV_0.XA20.XA3.MP5.D 17.6946
R14421 SUNSAR_SAR8B_CV_0.XA20.XA3.MP3.D SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n15 10.6968
R14422 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n4 SUNSAR_SAR8B_CV_0.XA20.XA2.MP5.G 10.633
R14423 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n13 SUNSAR_SAR8B_CV_0.XA20.XA2a.MP0.G 10.633
R14424 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n15 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n14 8.5257
R14425 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n4 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n3 5.42812
R14426 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n13 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n12 5.42812
R14427 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n14 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n4 5.08753
R14428 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n14 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n13 4.24194
R14429 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t6 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t7 1060.4
R14430 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t7 SUNSAR_CAPT8B_CV_0.XI14.XA2.MN0.G 589.284
R14431 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t3 572.893
R14432 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t4 572.893
R14433 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t2 572.893
R14434 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t5 568.956
R14435 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t6 568.956
R14436 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t1 356.344
R14437 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.t0 135.293
R14438 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XI14.XA1.MN0.D 115.954
R14439 SUNSAR_CAPT8B_CV_0.XI14.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n13 85.0829
R14440 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n5 22.1005
R14441 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XI14.XA2.MP0.G 20.3299
R14442 SUNSAR_CAPT8B_CV_0.XI14.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n2 15.2303
R14443 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.G 15.1965
R14444 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.G 15.1965
R14445 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.G 15.1965
R14446 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.G 13.5534
R14447 SUNSAR_CAPT8B_CV_0.XI14.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n12 13.5534
R14448 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n0 12.8005
R14449 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n1 12.6805
R14450 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n3 9.49168
R14451 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n7 9.3005
R14452 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n11 9.3005
R14453 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n4 9.10273
R14454 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n6 6.77697
R14455 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n0 6.77697
R14456 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n9 5.70934
R14457 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n10 3.40124
R14458 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n8 1.79829
R14459 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n5 0.191676
R14460 SUNSAR_SAR8B_CV_0.XA5.CP0.t8 SUNSAR_SAR8B_CV_0.XA5.CP0.t10 1060.4
R14461 SUNSAR_SAR8B_CV_0.XA5.CP0.t15 SUNSAR_SAR8B_CV_0.XA5.CP0.t9 1060.4
R14462 SUNSAR_SAR8B_CV_0.XA5.CP0.t13 SUNSAR_SAR8B_CV_0.XA5.CP0.t14 1060.4
R14463 SUNSAR_SAR8B_CV_0.XA5.CP0.t11 SUNSAR_SAR8B_CV_0.XA5.CP0.t12 1060.4
R14464 SUNSAR_SAR8B_CV_0.XA5.CP0.t10 SUNSAR_SAR8B_CV_0.XA5.CP0.n1 568.956
R14465 SUNSAR_SAR8B_CV_0.XA5.CP0.n2 SUNSAR_SAR8B_CV_0.XA5.CP0.t8 568.956
R14466 SUNSAR_SAR8B_CV_0.XA5.CP0.t9 SUNSAR_SAR8B_CV_0.XA5.CP0.n3 568.956
R14467 SUNSAR_SAR8B_CV_0.XA5.CP0.n4 SUNSAR_SAR8B_CV_0.XA5.CP0.t15 568.956
R14468 SUNSAR_SAR8B_CV_0.XA5.CP0.n7 SUNSAR_SAR8B_CV_0.XA5.CP0.t13 568.956
R14469 SUNSAR_SAR8B_CV_0.XA5.CP0.t14 SUNSAR_SAR8B_CV_0.XA5.CP0.n6 568.956
R14470 SUNSAR_SAR8B_CV_0.XA5.CP0.n5 SUNSAR_SAR8B_CV_0.XA5.CP0.t11 568.956
R14471 SUNSAR_SAR8B_CV_0.XA5.CP0.t12 SUNSAR_SAR8B_CV_0.XA5.CP0.n0 568.956
R14472 SUNSAR_SAR8B_CV_0.XA5.CP0.n11 SUNSAR_SAR8B_CV_0.XA5.CP0.n10 292.5
R14473 SUNSAR_SAR8B_CV_0.XA5.CP0.n17 SUNSAR_SAR8B_CV_0.XA5.CP0.n16 292.5
R14474 SUNSAR_SAR8B_CV_0.XA5.CP0.n9 SUNSAR_SAR8B_CV_0.XA5.CP0 197.272
R14475 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.CP0.n14 112.829
R14476 SUNSAR_SAR8B_CV_0.XA5.CP0.n17 SUNSAR_SAR8B_CV_0.XA5.CP0.n15 111.059
R14477 SUNSAR_SAR8B_CV_0.XA5.CP0.n9 SUNSAR_SAR8B_CV_0.XA5.CP0.n8 92.5005
R14478 SUNSAR_SAR8B_CV_0.XA5.CP0.n12 SUNSAR_SAR8B_CV_0.XA5.CP0.n11 81.5064
R14479 SUNSAR_SAR8B_CV_0.XA5.CP0.n16 SUNSAR_SAR8B_CV_0.XA5.CP0.t2 63.8431
R14480 SUNSAR_SAR8B_CV_0.XA5.CP0.n16 SUNSAR_SAR8B_CV_0.XA5.CP0.t6 63.8431
R14481 SUNSAR_SAR8B_CV_0.XA5.CP0.n10 SUNSAR_SAR8B_CV_0.XA5.CP0.t5 63.8431
R14482 SUNSAR_SAR8B_CV_0.XA5.CP0.n10 SUNSAR_SAR8B_CV_0.XA5.CP0.t4 63.8431
R14483 SUNSAR_SAR8B_CV_0.XA5.CP0.n15 SUNSAR_SAR8B_CV_0.XA5.CP0.n13 53.4593
R14484 SUNSAR_SAR8B_CV_0.XA5.CP0.n8 SUNSAR_SAR8B_CV_0.XA5.CP0.t3 38.8894
R14485 SUNSAR_SAR8B_CV_0.XA5.CP0.n8 SUNSAR_SAR8B_CV_0.XA5.CP0.t7 38.8894
R14486 SUNSAR_SAR8B_CV_0.XA5.CP0.n14 SUNSAR_SAR8B_CV_0.XA5.CP0.t1 38.8894
R14487 SUNSAR_SAR8B_CV_0.XA5.CP0.n14 SUNSAR_SAR8B_CV_0.XA5.CP0.t0 38.8894
R14488 SUNSAR_SAR8B_CV_0.XA5.CP0.n13 SUNSAR_SAR8B_CV_0.XA5.CP0.n12 29.5534
R14489 SUNSAR_SAR8B_CV_0.XA5.CP0.n4 SUNSAR_SAR8B_CV_0.XA5.CP0.n1 20.3299
R14490 SUNSAR_SAR8B_CV_0.XA5.CP0.n1 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14491 SUNSAR_SAR8B_CV_0.XA5.CP0.n2 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14492 SUNSAR_SAR8B_CV_0.XA5.CP0.n3 SUNSAR_SAR8B_CV_0.XA5.CP0.n0 20.3299
R14493 SUNSAR_SAR8B_CV_0.XA5.CP0.n3 SUNSAR_SAR8B_CV_0.XA5.CP0.n2 20.3299
R14494 SUNSAR_SAR8B_CV_0.XA5.CP0.n3 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14495 SUNSAR_SAR8B_CV_0.XA5.CP0.n4 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14496 SUNSAR_SAR8B_CV_0.XA5.CP0.n6 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14497 SUNSAR_SAR8B_CV_0.XA5.CP0.n6 SUNSAR_SAR8B_CV_0.XA5.CP0.n5 20.3299
R14498 SUNSAR_SAR8B_CV_0.XA5.CP0.n5 SUNSAR_SAR8B_CV_0.XA5.CP0.n4 20.3299
R14499 SUNSAR_SAR8B_CV_0.XA5.CP0.n5 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14500 SUNSAR_SAR8B_CV_0.XA5.CP0.n0 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14501 SUNSAR_SAR8B_CV_0.XA5.CP0.n7 SUNSAR_SAR8B_CV_0.XA5.CP0.n0 20.3299
R14502 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.CP0.n7 20.3299
R14503 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.CP0.n9 20.3299
R14504 SUNSAR_SAR8B_CV_0.XA5.CP0.n11 SUNSAR_SAR8B_CV_0.XA5.CP0 20.3299
R14505 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.CP0.n17 20.3299
R14506 SUNSAR_SAR8B_CV_0.XA5.CP0.n13 SUNSAR_SAR8B_CV_0.XA5.CP0 17.6946
R14507 SUNSAR_SAR8B_CV_0.XA5.CP0.n15 SUNSAR_SAR8B_CV_0.XA5.CP0 17.6946
R14508 SUNSAR_SAR8B_CV_0.XA5.CP0.n12 SUNSAR_SAR8B_CV_0.XA5.CP0 10.3476
R14509 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t9 568.956
R14510 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t8 568.956
R14511 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n3 292.5
R14512 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n9 292.5
R14513 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n12 197.272
R14514 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n2 112.829
R14515 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n6 112.829
R14516 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n4 111.059
R14517 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t5 63.8431
R14518 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n9 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t7 63.8431
R14519 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t4 63.8431
R14520 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n3 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t6 63.8431
R14521 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n7 59.1064
R14522 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n5 53.4593
R14523 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n10 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n8 51.9534
R14524 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t2 38.8894
R14525 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n2 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t1 38.8894
R14526 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t0 38.8894
R14527 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n6 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.t3 38.8894
R14528 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n1 37.1229
R14529 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 20.3299
R14530 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n11 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 20.3299
R14531 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n11 20.3299
R14532 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n12 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 20.3299
R14533 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n10 20.3299
R14534 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n5 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 17.6946
R14535 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n7 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 17.6946
R14536 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 12.325
R14537 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 12.323
R14538 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n8 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 10.3476
R14539 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n0 9.98893
R14540 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n1 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.168144
R14541 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t4 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t6 1060.4
R14542 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t9 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t2 1060.4
R14543 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t8 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t5 1060.4
R14544 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t3 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t7 1060.4
R14545 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n1 568.956
R14546 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t4 568.956
R14547 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t2 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n3 568.956
R14548 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t9 568.956
R14549 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t8 568.956
R14550 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n6 568.956
R14551 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t3 568.956
R14552 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n0 568.956
R14553 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t0 356.344
R14554 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.t1 131.389
R14555 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n9 128.754
R14556 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n8 SUNSAR_SAR8B_CV_0.XA4.XA2.MP0.G 97.8829
R14557 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n1 20.3299
R14558 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n1 SUNSAR_SAR8B_CV_0.XA4.XA2.MN3.G 20.3299
R14559 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n2 SUNSAR_SAR8B_CV_0.XA4.XA2.MP3.G 20.3299
R14560 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n0 20.3299
R14561 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n2 20.3299
R14562 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n3 SUNSAR_SAR8B_CV_0.XA4.XA2.MP2.G 20.3299
R14563 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n4 SUNSAR_SAR8B_CV_0.XA4.XA2.MN2.G 20.3299
R14564 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA4.XA2.MN0.G 20.3299
R14565 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n6 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n5 20.3299
R14566 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n4 20.3299
R14567 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n5 SUNSAR_SAR8B_CV_0.XA4.XA2.MN1.G 20.3299
R14568 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n0 SUNSAR_SAR8B_CV_0.XA4.XA2.MP1.G 20.3299
R14569 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n7 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n0 20.3299
R14570 SUNSAR_SAR8B_CV_0.XA4.XA2.MP0.G SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n7 20.3299
R14571 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.D SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n8 20.3299
R14572 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n9 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.D 20.3299
R14573 ua[0] ua[0].t9 376.673
R14574 ua[0] ua[0].t1 151.719
R14575 ua[0] ua[0].t2 151.719
R14576 ua[0] ua[0].t0 151.719
R14577 ua[0] ua[0].t3 151.719
R14578 ua[0] ua[0].t5 151.719
R14579 ua[0] ua[0].t8 151.719
R14580 ua[0].n16 ua[0].t6 136.754
R14581 ua[0].n0 ua[0].t7 131.389
R14582 ua[0].n13 ua[0].t4 131.389
R14583 ua[0].n12 ua[0] 121.977
R14584 ua[0].n8 ua[0] 71.1534
R14585 ua[0] ua[0].n18 71.1534
R14586 ua[0].n9 ua[0].n8 53.4593
R14587 ua[0].n10 ua[0].n9 53.4593
R14588 ua[0].n11 ua[0].n10 53.4593
R14589 ua[0].n17 ua[0].n11 53.4593
R14590 ua[0].n18 ua[0].n17 53.4593
R14591 ua[0].n1 ua[0].n0 22.1005
R14592 ua[0].n8 ua[0] 17.6946
R14593 ua[0].n9 ua[0] 17.6946
R14594 ua[0].n10 ua[0] 17.6946
R14595 ua[0].n11 ua[0] 17.6946
R14596 ua[0].n17 ua[0] 17.6946
R14597 ua[0].n18 ua[0] 17.6946
R14598 ua[0].n2 ua[0] 16.016
R14599 ua[0] ua[0].n7 13.5534
R14600 ua[0].n14 ua[0].n13 12.8005
R14601 ua[0] ua[0].n16 10.6968
R14602 ua[0].n15 ua[0].n12 9.49168
R14603 ua[0].n15 ua[0].n14 9.3005
R14604 ua[0].n7 ua[0].n6 9.3005
R14605 ua[0].n14 ua[0] 7.52991
R14606 ua[0].n16 ua[0].n15 6.95585
R14607 ua[0].n13 ua[0].n12 6.77697
R14608 ua[0].n7 ua[0].n0 6.77697
R14609 ua[0].n6 ua[0].n5 4.5005
R14610 ua[0].n3 ua[0].n1 4.5005
R14611 ua[0].n4 ua[0].n3 3.48238
R14612 ua[0].n5 ua[0].n4 3.4105
R14613 ua[0].n6 ua[0].n1 0.191676
R14614 ua[0].n5 ua[0].n2 0.0813824
R14615 ua[0].n4 ua[0] 0.0281471
R14616 ua[0].n3 ua[0].n2 0.00767963
R14617 uio_oe[0].n2 uio_oe[0] 1529.78
R14618 uio_oe[0].n1 uio_oe[0].t0 356.344
R14619 uio_oe[0].n1 uio_oe[0].n0 14.3064
R14620 uio_oe[0].n2 uio_oe[0].n1 8.50847
R14621 uio_oe[0].n0 uio_oe[0] 6.82717
R14622 uio_oe[0].n0 uio_oe[0] 6.02403
R14623 uio_oe[0] uio_oe[0].n2 0.448417
R14624 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t4 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t2 1060.4
R14625 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t2 SUNSAR_CAPT8B_CV_0.XG12.XA2.MN0.G 589.284
R14626 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t3 572.893
R14627 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t5 572.893
R14628 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t7 572.893
R14629 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t6 568.956
R14630 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t4 568.956
R14631 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n0 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t1 356.344
R14632 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.t0 135.293
R14633 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XG12.XA1.MN0.D 115.954
R14634 SUNSAR_CAPT8B_CV_0.XG12.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n13 85.0829
R14635 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n6 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n5 22.1005
R14636 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n13 SUNSAR_CAPT8B_CV_0.XG12.XA2.MP0.G 20.3299
R14637 SUNSAR_CAPT8B_CV_0.XG12.XA1.MN0.D SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n2 15.2303
R14638 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n1 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.G 15.1965
R14639 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n4 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.G 15.1965
R14640 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n9 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.G 15.1965
R14641 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.G 13.5534
R14642 SUNSAR_CAPT8B_CV_0.XG12.XA1.MP0.D SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n12 13.5534
R14643 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n3 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n0 12.8005
R14644 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n2 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n1 12.6805
R14645 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n3 9.49168
R14646 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n7 9.3005
R14647 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n11 9.3005
R14648 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n5 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n4 9.10273
R14649 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n7 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n6 6.77697
R14650 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n12 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n0 6.77697
R14651 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n9 5.70934
R14652 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n11 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n10 3.40124
R14653 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n10 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n8 1.79829
R14654 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n8 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n5 0.191676
R14655 uio_out[0].n3 uio_out[0] 3295.43
R14656 uio_out[0] uio_out[0].t1 379.384
R14657 uio_out[0].n2 uio_out[0] 140.198
R14658 uio_out[0].n1 uio_out[0].t0 131.389
R14659 uio_out[0].n1 uio_out[0].n0 14.3064
R14660 uio_out[0].n0 uio_out[0] 6.82717
R14661 uio_out[0].n3 uio_out[0].n2 6.3217
R14662 uio_out[0].n0 uio_out[0] 6.02403
R14663 uio_out[0].n2 uio_out[0].n1 3.01226
R14664 uio_out[0] uio_out[0].n3 0.140083
R14665 SUNSAR_SAR8B_CV_0.D<0>.t11 SUNSAR_SAR8B_CV_0.D<0>.t8 1060.4
R14666 SUNSAR_SAR8B_CV_0.D<0>.t8 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.G 589.284
R14667 SUNSAR_SAR8B_CV_0.D<0>.n11 SUNSAR_SAR8B_CV_0.D<0>.t11 573.85
R14668 SUNSAR_SAR8B_CV_0.D<0>.n3 SUNSAR_SAR8B_CV_0.D<0>.t9 568.956
R14669 SUNSAR_SAR8B_CV_0.D<0>.n2 SUNSAR_SAR8B_CV_0.D<0>.t10 568.956
R14670 SUNSAR_SAR8B_CV_0.D<0>.n1 SUNSAR_SAR8B_CV_0.D<0>.n0 292.5
R14671 SUNSAR_SAR8B_CV_0.D<0>.n22 SUNSAR_SAR8B_CV_0.D<0>.n21 292.5
R14672 SUNSAR_SAR8B_CV_0.XA7.XA3.MN0.D SUNSAR_SAR8B_CV_0.D<0>.n8 112.829
R14673 SUNSAR_SAR8B_CV_0.XA7.XA3.MN2.D SUNSAR_SAR8B_CV_0.D<0>.n19 112.829
R14674 SUNSAR_SAR8B_CV_0.D<0>.n22 SUNSAR_SAR8B_CV_0.D<0>.n20 111.059
R14675 SUNSAR_SAR8B_CV_0.D<0>.n9 SUNSAR_SAR8B_CV_0.D<0>.n7 89.224
R14676 SUNSAR_SAR8B_CV_0.D<0>.n21 SUNSAR_SAR8B_CV_0.D<0>.t4 63.8431
R14677 SUNSAR_SAR8B_CV_0.D<0>.n21 SUNSAR_SAR8B_CV_0.D<0>.t5 63.8431
R14678 SUNSAR_SAR8B_CV_0.D<0>.n0 SUNSAR_SAR8B_CV_0.D<0>.t6 63.8431
R14679 SUNSAR_SAR8B_CV_0.D<0>.n0 SUNSAR_SAR8B_CV_0.D<0>.t7 63.8431
R14680 SUNSAR_SAR8B_CV_0.D<0>.n20 SUNSAR_SAR8B_CV_0.D<0>.n18 48.7856
R14681 SUNSAR_SAR8B_CV_0.D<0>.n8 SUNSAR_SAR8B_CV_0.D<0>.t1 38.8894
R14682 SUNSAR_SAR8B_CV_0.D<0>.n8 SUNSAR_SAR8B_CV_0.D<0>.t0 38.8894
R14683 SUNSAR_SAR8B_CV_0.D<0>.n19 SUNSAR_SAR8B_CV_0.D<0>.t3 38.8894
R14684 SUNSAR_SAR8B_CV_0.D<0>.n19 SUNSAR_SAR8B_CV_0.D<0>.t2 38.8894
R14685 SUNSAR_SAR8B_CV_0.D<0>.n2 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.G 20.3299
R14686 SUNSAR_SAR8B_CV_0.D<0>.n3 SUNSAR_SAR8B_CV_0.D<0>.n2 20.3299
R14687 SUNSAR_SAR8B_CV_0.XA7.XA3.MP2.D SUNSAR_SAR8B_CV_0.D<0>.n22 20.3299
R14688 SUNSAR_SAR8B_CV_0.D<0>.n16 SUNSAR_SAR8B_CV_0.D<0>.n9 17.9961
R14689 SUNSAR_SAR8B_CV_0.D<0>.n20 SUNSAR_SAR8B_CV_0.XA7.XA3.MN2.D 17.6946
R14690 SUNSAR_SAR8B_CV_0.D<0>.n4 SUNSAR_SAR8B_CV_0.XA7.XA6.MP2.G 15.2303
R14691 SUNSAR_SAR8B_CV_0.D<0>.n5 SUNSAR_SAR8B_CV_0.XA7.XA3.MP0.D 13.5534
R14692 SUNSAR_SAR8B_CV_0.D<0>.n11 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN0.G 12.939
R14693 SUNSAR_SAR8B_CV_0.D<0>.n7 SUNSAR_SAR8B_CV_0.D<0>.n1 12.8005
R14694 SUNSAR_SAR8B_CV_0.D<0>.n9 SUNSAR_SAR8B_CV_0.XA7.XA3.MN0.D 11.2946
R14695 SUNSAR_SAR8B_CV_0.D<0>.n6 SUNSAR_SAR8B_CV_0.D<0>.n4 11.2842
R14696 SUNSAR_SAR8B_CV_0.D<0>.n12 SUNSAR_SAR8B_CV_0.D<0>.n11 10.501
R14697 SUNSAR_SAR8B_CV_0.D<0>.n7 SUNSAR_SAR8B_CV_0.D<0>.n6 9.49168
R14698 SUNSAR_SAR8B_CV_0.D<0>.n13 SUNSAR_SAR8B_CV_0.D<0>.n12 9.36597
R14699 SUNSAR_SAR8B_CV_0.D<0>.n6 SUNSAR_SAR8B_CV_0.D<0>.n5 9.3005
R14700 SUNSAR_SAR8B_CV_0.D<0>.n18 SUNSAR_SAR8B_CV_0.D<0>.n17 9.3005
R14701 SUNSAR_SAR8B_CV_0.D<0>.n18 SUNSAR_SAR8B_CV_0.D<0>.n9 8.11757
R14702 SUNSAR_SAR8B_CV_0.D<0>.n5 SUNSAR_SAR8B_CV_0.D<0>.n1 6.77697
R14703 SUNSAR_SAR8B_CV_0.D<0>.n17 SUNSAR_SAR8B_CV_0.D<0>.n10 4.5005
R14704 SUNSAR_SAR8B_CV_0.D<0>.n16 SUNSAR_SAR8B_CV_0.D<0>.n15 4.5005
R14705 SUNSAR_SAR8B_CV_0.D<0>.n4 SUNSAR_SAR8B_CV_0.D<0>.n3 3.90429
R14706 SUNSAR_SAR8B_CV_0.D<0>.n13 SUNSAR_SAR8B_CV_0.D<0>.n10 3.4105
R14707 SUNSAR_SAR8B_CV_0.D<0>.n15 SUNSAR_SAR8B_CV_0.D<0>.n14 3.4105
R14708 SUNSAR_SAR8B_CV_0.D<0>.n15 SUNSAR_SAR8B_CV_0.D<0>.n10 0.191676
R14709 SUNSAR_SAR8B_CV_0.D<0>.n17 SUNSAR_SAR8B_CV_0.D<0>.n16 0.191676
R14710 SUNSAR_SAR8B_CV_0.D<0>.n12 SUNSAR_CAPT8B_CV_0.D<0> 0.173294
R14711 SUNSAR_SAR8B_CV_0.D<0>.n14 SUNSAR_SAR8B_CV_0.D<0>.n13 0.0713406
R14712 SUNSAR_SAR8B_CV_0.D<0>.n14 SUNSAR_SAR8B_CV_0.XA7.CP1 0.0277464
R14713 uo_out[7].t2 uo_out[7].t3 1060.4
R14714 uo_out[7].t3 uo_out[7] 589.284
R14715 uo_out[7].n0 uo_out[7].t2 574.383
R14716 uo_out[7].n1 uo_out[7].t1 361.707
R14717 uo_out[7].n3 uo_out[7].t0 131.389
R14718 uo_out[7].n2 uo_out[7] 118.966
R14719 uo_out[7].n6 uo_out[7] 14.887
R14720 uo_out[7] uo_out[7].n1 10.6968
R14721 uo_out[7].n0 uo_out[7] 10.633
R14722 uo_out[7].n4 uo_out[7] 10.5417
R14723 uo_out[7].n3 uo_out[7].n2 9.78874
R14724 uo_out[7].n4 uo_out[7].n3 9.78874
R14725 uo_out[7].n1 uo_out[7].n0 9.53185
R14726 uo_out[7].n5 uo_out[7].n2 9.39464
R14727 uo_out[7].n5 uo_out[7].n4 9.39464
R14728 uo_out[7].n6 uo_out[7].n5 2.54977
R14729 uo_out[7] uo_out[7].n6 0.199029
R14730 SUNSAR_SAR8B_CV_0.XB2.CKN.t6 SUNSAR_SAR8B_CV_0.XB2.CKN.t4 1060.4
R14731 SUNSAR_SAR8B_CV_0.XB2.CKN.t2 SUNSAR_SAR8B_CV_0.XB2.CKN.t7 1060.4
R14732 SUNSAR_SAR8B_CV_0.XB2.CKN.t4 SUNSAR_SAR8B_CV_0.XB2.XA4.MP0.G 589.284
R14733 SUNSAR_SAR8B_CV_0.XB2.CKN.n11 SUNSAR_SAR8B_CV_0.XB2.CKN.t6 574.351
R14734 SUNSAR_SAR8B_CV_0.XB2.CKN.n3 SUNSAR_SAR8B_CV_0.XB2.CKN.t3 568.956
R14735 SUNSAR_SAR8B_CV_0.XB2.CKN.t7 SUNSAR_SAR8B_CV_0.XB2.CKN.n4 568.956
R14736 SUNSAR_SAR8B_CV_0.XB2.CKN.n5 SUNSAR_SAR8B_CV_0.XB2.CKN.t2 568.956
R14737 SUNSAR_SAR8B_CV_0.XB2.CKN.n1 SUNSAR_SAR8B_CV_0.XB2.CKN.t5 568.956
R14738 SUNSAR_SAR8B_CV_0.XB2.CKN.n8 SUNSAR_SAR8B_CV_0.XB2.CKN.t1 361.707
R14739 SUNSAR_SAR8B_CV_0.XB2.CKN.n0 SUNSAR_SAR8B_CV_0.XB2.CKN.t0 131.389
R14740 SUNSAR_SAR8B_CV_0.XB2.CKN.n2 SUNSAR_SAR8B_CV_0.XB2.CKN.n1 122.73
R14741 SUNSAR_SAR8B_CV_0.XB2.CKN.n9 SUNSAR_SAR8B_CV_0.XB2.XA0.MP0.D 114.448
R14742 SUNSAR_SAR8B_CV_0.XB2.CKN.n9 SUNSAR_SAR8B_CV_0.XB2.XA0.MN0.D 34.6358
R14743 SUNSAR_SAR8B_CV_0.XB2.CKN.n3 SUNSAR_SAR8B_CV_0.XB2.XA3.MN1.G 20.3299
R14744 SUNSAR_SAR8B_CV_0.XB2.CKN.n4 SUNSAR_SAR8B_CV_0.XB2.CKN.n3 20.3299
R14745 SUNSAR_SAR8B_CV_0.XB2.CKN.n4 SUNSAR_SAR8B_CV_0.XB2.XA3.MN0.G 20.3299
R14746 SUNSAR_SAR8B_CV_0.XB2.CKN.n1 SUNSAR_SAR8B_CV_0.XB2.XA3.MP2.G 20.3299
R14747 SUNSAR_SAR8B_CV_0.XB2.CKN.n6 SUNSAR_SAR8B_CV_0.XB2.CKN.n5 12.8005
R14748 SUNSAR_SAR8B_CV_0.XB2.XA0.MP0.D SUNSAR_SAR8B_CV_0.XB2.CKN.n8 10.6968
R14749 SUNSAR_SAR8B_CV_0.XB2.CKN.n11 SUNSAR_SAR8B_CV_0.XB2.XA4.MN0.G 10.6653
R14750 SUNSAR_SAR8B_CV_0.XB2.CKN.n12 SUNSAR_SAR8B_CV_0.XB2.CKN.n11 10.6568
R14751 SUNSAR_SAR8B_CV_0.XB2.CKN.n7 SUNSAR_SAR8B_CV_0.XB2.CKN.n2 9.49168
R14752 SUNSAR_SAR8B_CV_0.XB2.CKN.n12 SUNSAR_SAR8B_CV_0.XB2.CKN.n10 9.39659
R14753 SUNSAR_SAR8B_CV_0.XB2.CKN.n13 SUNSAR_SAR8B_CV_0.XB2.CKN.n12 9.39269
R14754 SUNSAR_SAR8B_CV_0.XB2.CKN.n7 SUNSAR_SAR8B_CV_0.XB2.CKN.n6 9.3005
R14755 SUNSAR_SAR8B_CV_0.XB2.CKN.n13 SUNSAR_SAR8B_CV_0.XB2.CKN.n0 8.53383
R14756 SUNSAR_SAR8B_CV_0.XB2.CKN.n6 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.G 7.52991
R14757 SUNSAR_SAR8B_CV_0.XB2.CKN.n5 SUNSAR_SAR8B_CV_0.XB2.CKN.n2 6.77697
R14758 SUNSAR_SAR8B_CV_0.XB2.CKN.n10 SUNSAR_SAR8B_CV_0.XB2.CKN.n9 5.02011
R14759 SUNSAR_SAR8B_CV_0.XB2.XA0.MN0.D SUNSAR_SAR8B_CV_0.XB2.CKN.n13 5.02011
R14760 SUNSAR_SAR8B_CV_0.XB2.CKN.n8 SUNSAR_SAR8B_CV_0.XB2.CKN.n7 4.94114
R14761 SUNSAR_SAR8B_CV_0.XB2.CKN.n10 SUNSAR_SAR8B_CV_0.XB2.CKN.n0 4.51815
R14762 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t4 1060.4
R14763 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t8 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t2 1060.4
R14764 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t9 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t6 1060.4
R14765 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t5 1060.4
R14766 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n1 568.956
R14767 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t3 568.956
R14768 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t2 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n3 568.956
R14769 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t8 568.956
R14770 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t9 568.956
R14771 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n6 568.956
R14772 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t7 568.956
R14773 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n0 568.956
R14774 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t0 356.344
R14775 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.t1 135.293
R14776 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n10 128.754
R14777 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n1 20.3299
R14778 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n1 SUNSAR_SAR8B_CV_0.XA5.XA4.MP3.G 20.3299
R14779 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n2 SUNSAR_SAR8B_CV_0.XA5.XA4.MN3.G 20.3299
R14780 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n0 20.3299
R14781 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n2 20.3299
R14782 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n3 SUNSAR_SAR8B_CV_0.XA5.XA4.MN2.G 20.3299
R14783 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n4 SUNSAR_SAR8B_CV_0.XA5.XA4.MP2.G 20.3299
R14784 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA5.XA4.MP0.G 20.3299
R14785 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n6 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n5 20.3299
R14786 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n4 20.3299
R14787 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n5 SUNSAR_SAR8B_CV_0.XA5.XA4.MP1.G 20.3299
R14788 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n0 SUNSAR_SAR8B_CV_0.XA5.XA4.MN1.G 20.3299
R14789 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n7 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n0 20.3299
R14790 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n10 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.D 20.3299
R14791 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n9 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n8 16.3643
R14792 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.D SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n9 15.2303
R14793 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA5.XA4.MN0.G 15.1965
R14794 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n8 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n7 3.93805
R14795 uo_out[6].t3 uo_out[6].t2 1060.4
R14796 uo_out[6].t2 uo_out[6] 589.284
R14797 uo_out[6].n1 uo_out[6].t3 572.859
R14798 uo_out[6].n0 uo_out[6].t1 356.344
R14799 uo_out[6].n5 uo_out[6].t0 136.285
R14800 uo_out[6] uo_out[6].n4 115.954
R14801 uo_out[6].n1 uo_out[6] 15.2303
R14802 uo_out[6].n2 uo_out[6] 13.5534
R14803 uo_out[6].n5 uo_out[6] 12.939
R14804 uo_out[6].n4 uo_out[6].n0 12.8005
R14805 uo_out[6].n6 uo_out[6] 12.6596
R14806 uo_out[6].n4 uo_out[6].n3 9.49168
R14807 uo_out[6].n3 uo_out[6].n2 9.3005
R14808 uo_out[6].n6 uo_out[6].n5 7.24734
R14809 uo_out[6].n3 uo_out[6].n1 7.07827
R14810 uo_out[6].n2 uo_out[6].n0 6.77697
R14811 uo_out[6] uo_out[6].n6 0.199029
R14812 ui_in[0].t1 ui_in[0].t0 1060.4
R14813 ui_in[0].t0 ui_in[0] 589.284
R14814 ui_in[0].n0 ui_in[0].t1 572.875
R14815 ui_in[0].n0 ui_in[0] 15.2133
R14816 ui_in[0] ui_in[0].n0 10.3815
R14817 SUNSAR_SAR8B_CV_0.XA7.ENO.t5 SUNSAR_SAR8B_CV_0.XA7.ENO.t4 1060.4
R14818 SUNSAR_SAR8B_CV_0.XA7.ENO.t2 SUNSAR_SAR8B_CV_0.XA7.ENO.t3 1060.4
R14819 SUNSAR_SAR8B_CV_0.XA7.ENO.t4 SUNSAR_SAR8B_CV_0.XA7.ENO 589.284
R14820 SUNSAR_SAR8B_CV_0.XA7.ENO.t3 SUNSAR_SAR8B_CV_0.XA7.ENO 589.284
R14821 SUNSAR_SAR8B_CV_0.XA7.ENO.n1 SUNSAR_SAR8B_CV_0.XA7.ENO.t2 583.638
R14822 SUNSAR_SAR8B_CV_0.XA7.ENO.n5 SUNSAR_SAR8B_CV_0.XA7.ENO.t5 572.893
R14823 SUNSAR_SAR8B_CV_0.XA7.ENO.n0 SUNSAR_SAR8B_CV_0.XA7.ENO.t0 356.344
R14824 SUNSAR_SAR8B_CV_0.XA7.ENO.n3 SUNSAR_SAR8B_CV_0.XA7.ENO 268.8
R14825 SUNSAR_SAR8B_CV_0.XA7.ENO.n2 SUNSAR_SAR8B_CV_0.XA7.ENO.t1 131.389
R14826 SUNSAR_SAR8B_CV_0.XA7.ENO.n2 SUNSAR_SAR8B_CV_0.XA7.ENO.n1 90.7299
R14827 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.ENO.n2 20.3299
R14828 SUNSAR_SAR8B_CV_0.XA7.ENO.n7 SUNSAR_SAR8B_CV_0.XA7.ENO.n5 20.0513
R14829 SUNSAR_SAR8B_CV_0.XA7.ENO.n5 SUNSAR_SAR8B_CV_0.XA7.ENO 15.1965
R14830 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.ENO.n9 13.5534
R14831 SUNSAR_SAR8B_CV_0.XA7.ENO.n3 SUNSAR_SAR8B_CV_0.XA7.ENO.n0 12.8005
R14832 SUNSAR_SAR8B_CV_0.XA7.ENO.n4 SUNSAR_SAR8B_CV_0.XA7.ENO.n3 9.35932
R14833 SUNSAR_SAR8B_CV_0.XA7.ENO.n9 SUNSAR_SAR8B_CV_0.XA7.ENO.n8 9.3005
R14834 SUNSAR_SAR8B_CV_0.XA7.ENO.n9 SUNSAR_SAR8B_CV_0.XA7.ENO.n0 6.77697
R14835 SUNSAR_SAR8B_CV_0.XA7.ENO.n1 SUNSAR_SAR8B_CV_0.XA7.ENO 5.64756
R14836 SUNSAR_SAR8B_CV_0.XA7.ENO.n6 SUNSAR_SAR8B_CV_0.XA7.ENO.n4 4.69168
R14837 SUNSAR_SAR8B_CV_0.XA7.ENO.n7 SUNSAR_SAR8B_CV_0.XA7.ENO.n6 4.5005
R14838 SUNSAR_SAR8B_CV_0.XA7.ENO.n8 SUNSAR_SAR8B_CV_0.XA7.ENO.n4 0.132853
R14839 SUNSAR_SAR8B_CV_0.XA7.ENO.n6 SUNSAR_SAR8B_CV_0.XA7.ENO 0.0740294
R14840 SUNSAR_SAR8B_CV_0.XA7.ENO.n8 SUNSAR_SAR8B_CV_0.XA7.ENO.n7 0.0593235
R14841 uo_out[1].t2 uo_out[1].t3 1060.4
R14842 uo_out[1].t3 uo_out[1] 589.284
R14843 uo_out[1].n0 uo_out[1].t2 574.383
R14844 uo_out[1].n1 uo_out[1].t1 361.707
R14845 uo_out[1].n3 uo_out[1].t0 131.389
R14846 uo_out[1].n2 uo_out[1] 118.966
R14847 uo_out[1] uo_out[1].n1 10.6968
R14848 uo_out[1].n0 uo_out[1] 10.633
R14849 uo_out[1].n4 uo_out[1] 10.5417
R14850 uo_out[1].n3 uo_out[1].n2 9.78874
R14851 uo_out[1].n4 uo_out[1].n3 9.78874
R14852 uo_out[1].n1 uo_out[1].n0 9.53185
R14853 uo_out[1].n5 uo_out[1].n2 9.39464
R14854 uo_out[1].n5 uo_out[1].n4 9.39464
R14855 uo_out[1].n6 uo_out[1] 8.67651
R14856 uo_out[1].n6 uo_out[1].n5 2.56815
R14857 uo_out[1] uo_out[1].n6 0.180647
R14858 uo_out[2].t3 uo_out[2].t2 1060.4
R14859 uo_out[2].t2 uo_out[2] 589.284
R14860 uo_out[2].n1 uo_out[2].t3 572.859
R14861 uo_out[2].n0 uo_out[2].t1 356.344
R14862 uo_out[2].n5 uo_out[2].t0 136.285
R14863 uo_out[2] uo_out[2].n4 115.954
R14864 uo_out[2].n1 uo_out[2] 15.2303
R14865 uo_out[2].n2 uo_out[2] 13.5534
R14866 uo_out[2].n5 uo_out[2] 12.939
R14867 uo_out[2].n4 uo_out[2].n0 12.8005
R14868 uo_out[2].n4 uo_out[2].n3 9.49168
R14869 uo_out[2].n3 uo_out[2].n2 9.3005
R14870 uo_out[2].n6 uo_out[2] 7.74629
R14871 uo_out[2].n6 uo_out[2].n5 7.25101
R14872 uo_out[2].n3 uo_out[2].n1 7.07827
R14873 uo_out[2].n2 uo_out[2].n0 6.77697
R14874 uo_out[2] uo_out[2].n6 0.195353
R14875 uo_out[4].t3 uo_out[4].t2 1060.4
R14876 uo_out[4].t2 uo_out[4] 589.284
R14877 uo_out[4].n1 uo_out[4].t3 572.859
R14878 uo_out[4].n0 uo_out[4].t1 356.344
R14879 uo_out[4].n5 uo_out[4].t0 136.285
R14880 uo_out[4] uo_out[4].n4 115.954
R14881 uo_out[4].n1 uo_out[4] 15.2303
R14882 uo_out[4].n2 uo_out[4] 13.5534
R14883 uo_out[4].n5 uo_out[4] 12.939
R14884 uo_out[4].n4 uo_out[4].n0 12.8005
R14885 uo_out[4].n6 uo_out[4] 10.1297
R14886 uo_out[4].n4 uo_out[4].n3 9.49168
R14887 uo_out[4].n3 uo_out[4].n2 9.3005
R14888 uo_out[4].n6 uo_out[4].n5 7.24734
R14889 uo_out[4].n3 uo_out[4].n1 7.07827
R14890 uo_out[4].n2 uo_out[4].n0 6.77697
R14891 uo_out[4] uo_out[4].n6 0.199029
R14892 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n80 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n0 297.865
R14893 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n73 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n72 91.8472
R14894 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n72 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n69 91.8472
R14895 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n10 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n9 91.8472
R14896 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n9 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n6 91.8472
R14897 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n25 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n24 91.8472
R14898 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n24 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n21 91.8472
R14899 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n41 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n40 91.8472
R14900 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n40 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n37 91.8472
R14901 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n57 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n56 91.8472
R14902 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n56 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n53 91.8472
R14903 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n0 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.t0 63.8431
R14904 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n0 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.t1 63.8431
R14905 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n72 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n71 49.1805
R14906 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n9 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n8 49.1805
R14907 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n24 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n23 49.1805
R14908 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n40 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n39 49.1805
R14909 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n56 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n55 49.1805
R14910 SUNSAR_SAR8B_CV_0.XB2.XA4.MP0.D SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n80 10.6968
R14911 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n80 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n79 9.0349
R14912 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n77 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n76 2.03137
R14913 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n14 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n13 2.03137
R14914 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n29 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n28 2.03137
R14915 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n45 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n44 2.03137
R14916 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n61 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n60 2.03137
R14917 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n76 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n75 2.03137
R14918 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n13 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n12 2.03137
R14919 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n28 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n27 2.03137
R14920 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n44 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n43 2.03137
R14921 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n60 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n59 2.03137
R14922 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n76 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n66 1.8747
R14923 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n13 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n3 1.8747
R14924 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n28 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n18 1.8747
R14925 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n44 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n34 1.8747
R14926 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n60 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n50 1.8747
R14927 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n74 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n73 1.5005
R14928 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n69 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n65 1.5005
R14929 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n71 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n70 1.5005
R14930 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n11 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n10 1.5005
R14931 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n6 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n2 1.5005
R14932 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n8 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n7 1.5005
R14933 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n26 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n25 1.5005
R14934 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n21 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n17 1.5005
R14935 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n23 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n22 1.5005
R14936 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n42 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n41 1.5005
R14937 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n37 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n33 1.5005
R14938 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n39 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n38 1.5005
R14939 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n58 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n57 1.5005
R14940 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n53 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n49 1.5005
R14941 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n55 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n54 1.5005
R14942 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n75 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n74 1.13717
R14943 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n70 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n66 1.13717
R14944 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n77 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n65 1.13717
R14945 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n12 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n11 1.13717
R14946 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n7 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n3 1.13717
R14947 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n14 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n2 1.13717
R14948 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n27 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n26 1.13717
R14949 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n22 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n18 1.13717
R14950 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n29 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n17 1.13717
R14951 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n43 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n42 1.13717
R14952 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n38 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n34 1.13717
R14953 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n45 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n33 1.13717
R14954 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n59 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n58 1.13717
R14955 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n54 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n50 1.13717
R14956 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n61 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n49 1.13717
R14957 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n74 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n67 0.867167
R14958 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n73 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n68 0.867167
R14959 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n69 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n68 0.867167
R14960 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n67 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n65 0.867167
R14961 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n11 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n4 0.867167
R14962 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n10 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n5 0.867167
R14963 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n6 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n5 0.867167
R14964 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n4 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n2 0.867167
R14965 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n26 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n19 0.867167
R14966 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n25 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n20 0.867167
R14967 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n21 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n20 0.867167
R14968 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n19 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n17 0.867167
R14969 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n42 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n35 0.867167
R14970 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n41 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n36 0.867167
R14971 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n37 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n36 0.867167
R14972 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n35 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n33 0.867167
R14973 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n58 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n51 0.867167
R14974 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n57 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n52 0.867167
R14975 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n53 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n52 0.867167
R14976 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n51 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n49 0.867167
R14977 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n31 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB4.A 0.682
R14978 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n79 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB0.A 0.625324
R14979 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n47 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n31 0.617029
R14980 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n63 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n47 0.617029
R14981 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n71 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n68 0.4505
R14982 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n70 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n67 0.4505
R14983 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n8 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n5 0.4505
R14984 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n7 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n4 0.4505
R14985 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n23 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n20 0.4505
R14986 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n22 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n19 0.4505
R14987 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n39 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n36 0.4505
R14988 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n38 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n35 0.4505
R14989 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n55 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n52 0.4505
R14990 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n54 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n51 0.4505
R14991 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n75 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n64 0.326367
R14992 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n12 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n1 0.326367
R14993 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n27 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n16 0.326367
R14994 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n43 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n32 0.326367
R14995 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n59 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n48 0.326367
R14996 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n66 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n64 0.1697
R14997 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n78 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n77 0.1697
R14998 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n3 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n1 0.1697
R14999 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n15 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n14 0.1697
R15000 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n18 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n16 0.1697
R15001 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n30 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n29 0.1697
R15002 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n34 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n32 0.1697
R15003 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n46 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n45 0.1697
R15004 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n50 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n48 0.1697
R15005 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n62 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n61 0.1697
R15006 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n78 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n64 0.157167
R15007 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n15 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n1 0.157167
R15008 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n30 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n16 0.157167
R15009 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n46 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n32 0.157167
R15010 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n62 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n48 0.157167
R15011 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n31 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB3.A 0.0654706
R15012 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n47 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB2.A 0.0654706
R15013 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n63 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB1.A 0.0654706
R15014 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB0.A SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n78 0.02165
R15015 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB4.A SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n15 0.02165
R15016 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB3.A SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n30 0.02165
R15017 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB2.A SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n46 0.02165
R15018 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n62 0.02165
R15019 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n79 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n63 0.0101765
C0 VPWR a_8802_36300# 0.399161f
C1 VPWR a_3762_37180# 0.473713f
C2 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C3 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.375196f
C4 SUNSAR_SAR8B_CV_0.XA0.XA12.A a_2610_36828# 0.10248f
C5 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.158152f
C6 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.XA7.CN 0.306905f
C7 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S 0.106927f
C8 VPWR a_18902_41000# 0.388256f
C9 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.432466f
C10 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.301665f
C11 uio_oe[0] uio_out[0] 1.55761f
C12 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 1.06002f
C13 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.55251f
C14 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C15 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_4390# 0.15559f
C16 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.15651f
C17 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C18 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.587991f
C19 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S 0.138148f
C20 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C21 VPWR a_5150_41880# 0.395781f
C22 VPWR a_5130_32956# 0.436368f
C23 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA6.A 1.63909f
C24 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<3> 0.297504f
C25 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C26 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S 0.112858f
C27 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_4390# 0.15559f
C28 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.30776f
C29 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.220689f
C30 VPWR a_5130_27148# 0.470364f
C31 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA7.CN 1.77562f
C32 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C33 VPWR a_5130_35420# 0.39968f
C34 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA20.CPO 0.255261f
C35 clk uio_out[0] 0.120689f
C36 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 1.06875f
C37 VPWR a_3782_41880# 0.395781f
C38 VPWR a_5130_36300# 0.398846f
C39 VPWR a_3762_32956# 0.436368f
C40 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S 0.104609f
C41 VPWR a_20250_37532# 0.454392f
C42 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C43 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.59087f
C44 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.29297f
C45 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_SAR8B_CV_0.D<2> 0.241356f
C46 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S 0.112858f
C47 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.128204f
C48 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.383512f
C49 VPWR a_3762_27148# 0.471462f
C50 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.22339f
C51 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S 0.106927f
C52 VPWR a_15230_41000# 0.388156f
C53 VPWR a_3762_35420# 0.39968f
C54 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.267238f
C55 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S 0.137646f
C56 uo_out[0] uio_out[0] 0.201579f
C57 clk uio_oe[0] 0.260056f
C58 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.164325f
C59 VPWR a_3762_36300# 0.399161f
C60 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.440586f
C61 SUNSAR_SAR8B_CV_0.XA0.XA11.A a_2610_36300# 0.13253f
C62 VPWR a_18882_37532# 0.458267f
C63 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C64 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.2622f
C65 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.377598f
C66 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.224309f
C67 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.308722f
C68 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_6282_35420# 0.160931f
C69 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.419738f
C70 VPWR a_13862_41000# 0.388256f
C71 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C72 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 1.05322f
C73 clk ui_in[0] 0.169609f
C74 uo_out[0] uio_oe[0] 0.670799f
C75 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.118162f
C76 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.A 0.744161f
C77 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 54.2165f
C78 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA6.A 1.63909f
C79 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<4> 0.297602f
C80 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.88588f
C81 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 3.09787f
C82 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.363295f
C83 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 1.77562f
C84 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_5130_35420# 0.133834f
C85 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C86 VPWR SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.106794f
C87 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S 0.138148f
C88 uo_out[1] uio_oe[0] 0.432144f
C89 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C90 VPWR SUNSAR_CAPT8B_CV_0.XA5.B 1.20019f
C91 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C92 VPWR a_23922_36652# 0.449853f
C93 VPWR a_23922_33132# 0.415713f
C94 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S 0.104609f
C95 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.665006f
C96 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.431984f
C97 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.151329f
C98 VPWR a_20250_27500# 0.382397f
C99 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.293159f
C100 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.527529f
C101 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.419738f
C102 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.432466f
C103 VPWR SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.658328f
C104 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 1.06875f
C105 uo_out[2] uio_oe[0] 0.267754f
C106 VPWR a_16542_4566# 0.413433f
C107 VPWR a_15210_37532# 0.459479f
C108 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.07164f
C109 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.B 0.545186f
C110 VPWR a_20250_34716# 0.396749f
C111 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.337652f
C112 VPWR a_18882_27500# 0.382189f
C113 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA4.CEIN 0.432008f
C114 VPWR SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.765792f
C115 VPWR a_10190_41000# 0.388175f
C116 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C117 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.62595f
C118 VPWR a_20250_31196# 0.437f
C119 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S 0.137646f
C120 uo_out[3] uio_oe[0] 0.212351f
C121 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C122 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.106927f
C123 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C124 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.718455f
C125 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 2.66621f
C126 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA6.A 1.63909f
C127 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.142061f
C128 VPWR a_13842_37532# 0.458324f
C129 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<5> 0.297941f
C130 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.316693f
C131 VPWR a_18882_34716# 0.399819f
C132 VPWR a_23922_29964# 0.429137f
C133 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.158152f
C134 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_3762_35420# 0.133834f
C135 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_2768# 0.172147f
C136 VPWR a_8822_41000# 0.388256f
C137 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.A 1.20972f
C138 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C139 VPWR a_18882_31196# 0.44007f
C140 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 1.05322f
C141 uo_out[4] uio_oe[0] 0.550054f
C142 uo_out[5] uio_out[0] 0.109219f
C143 uo_out[1] uo_out[0] 0.355472f
C144 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.106927f
C145 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S 0.101562f
C146 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 2.64055f
C147 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 6.86675f
C148 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.665006f
C149 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.42393f
C150 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.126806f
C151 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.1501f
C152 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_SAR8B_CV_0.D<3> 0.241356f
C153 VPWR a_20270_43816# 0.391817f
C154 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_2610_35420# 0.160931f
C155 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C156 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_42408# 0.100131f
C157 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.924613f
C158 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S 0.138148f
C159 VPWR ua[0] 0.51729f
C160 uo_out[5] uio_oe[0] 1.55329f
C161 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.119314f
C162 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L 1.05246f
C163 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 2.64054f
C164 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C165 uio_out[0] tt_um_TT06_SAR_done_0.x3.MP1.G 0.165429f
C166 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.375196f
C167 VPWR a_15210_27500# 0.382397f
C168 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.220689f
C169 VPWR a_18902_43816# 0.391817f
C170 ua[0] SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.247314f
C171 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.432466f
C172 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.A 1.22023f
C173 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 1.06875f
C174 VPWR ua[1] 0.225132f
C175 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.725614f
C176 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.704356f
C177 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 2.64055f
C178 VPWR a_9990_4566# 0.413433f
C179 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA6.A 1.63909f
C180 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C181 VPWR a_10170_37532# 0.459599f
C182 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<6> 0.298165f
C183 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.363295f
C184 VPWR a_15210_34716# 0.399819f
C185 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S 0.108436f
C186 VPWR a_13842_27500# 0.382189f
C187 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.527529f
C188 VPWR a_5150_41000# 0.388161f
C189 VPWR a_15210_31196# 0.44007f
C190 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S 0.137646f
C191 uo_out[7] uio_oe[0] 0.43252f
C192 VPWR uio_out[0] 0.408488f
C193 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C194 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.106927f
C195 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.722887f
C196 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 2.64054f
C197 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.452478f
C198 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43816# 0.129239f
C199 VPWR a_8802_37532# 0.458443f
C200 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.26537f
C201 VPWR a_13842_34716# 0.399819f
C202 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.279205f
C203 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.377598f
C204 VPWR a_3782_41000# 0.388256f
C205 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_3728# 0.172147f
C206 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.449584f
C207 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C208 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.930839f
C209 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C210 VPWR a_13842_31196# 0.44007f
C211 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 1.05322f
C212 uo_out[3] uo_out[2] 0.109993f
C213 VPWR uio_oe[0] 1.67769f
C214 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.106927f
C215 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.101979f
C216 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.7271f
C217 VPWR a_20250_29612# 0.398044f
C218 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1615f
C219 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.232115f
C220 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN 0.144331f
C221 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C222 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.268769f
C223 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_4742# 0.156331f
C224 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.383512f
C225 VPWR a_15230_43816# 0.391817f
C226 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.22339f
C227 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S 0.138148f
C228 VPWR ui_in[0] 1.85366f
C229 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.437693f
C230 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.426291f
C231 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.119314f
C232 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.15234f
C233 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.72582f
C234 VPWR a_18882_29612# 0.397362f
C235 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA6.A 1.63909f
C236 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<7> 0.294651f
C237 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.316693f
C238 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_4742# 0.156331f
C239 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.36754f
C240 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S 0.104609f
C241 VPWR a_10170_27500# 0.382397f
C242 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.293159f
C243 VPWR a_13862_43816# 0.391817f
C244 VPWR a_23942_41352# 0.376408f
C245 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.449584f
C246 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.165965f
C247 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.A 1.2202f
C248 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C249 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.138433f
C250 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 1.06875f
C251 VPWR clk 0.644902f
C252 uo_out[4] uo_out[3] 0.854997f
C253 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.725614f
C254 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.340491f
C255 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 2.72889f
C256 VPWR SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.519052f
C257 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.726497f
C258 VPWR a_5130_37532# 0.459538f
C259 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_41880# 0.100592f
C260 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.126806f
C261 VPWR a_10170_34716# 0.399819f
C262 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA2.CEIN 0.432008f
C263 VPWR a_8802_27500# 0.382189f
C264 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.93081f
C265 VPWR a_10170_31196# 0.44007f
C266 VPWR a_23922_28556# 0.499441f
C267 VPWR uo_out[0] 1.02382f
C268 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.106927f
C269 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.437693f
C270 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.722887f
C271 VPWR a_16542_4918# 0.470354f
C272 clk SUNSAR_CAPT8B_CV_0.XA6.A 0.206733f
C273 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43816# 0.127669f
C274 VPWR a_3762_37532# 0.458382f
C275 VPWR a_8802_34716# 0.399819f
C276 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.158152f
C277 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_4688# 0.172147f
C278 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.432466f
C279 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.A 1.22023f
C280 VPWR a_8802_31196# 0.44007f
C281 VPWR uo_out[1] 1.02322f
C282 uo_out[5] uo_out[4] 1.16093f
C283 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.106927f
C284 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.101979f
C285 VPWR a_20250_33836# 0.407174f
C286 VPWR a_15210_29612# 0.397362f
C287 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6519f
C288 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA6.A 1.63909f
C289 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_SAR8B_CV_0.D<4> 0.241356f
C290 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.363295f
C291 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.175967f
C292 VPWR a_10190_43816# 0.391817f
C293 VPWR a_20270_41352# 0.394053f
C294 uo_out[6] uo_out[4] 0.843602f
C295 VPWR uo_out[2] 1.02322f
C296 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.119314f
C297 VPWR a_18882_33836# 0.409601f
C298 ua[0] SUNSAR_SAR8B_CV_0.SARN 1.02347f
C299 VPWR a_13842_29612# 0.397362f
C300 VPWR SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.519052f
C301 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN 0.144331f
C302 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_21402_35068# 0.129098f
C303 SUNSAR_CAPT8B_CV_0.XG12.QN a_16382_43816# 0.129239f
C304 VPWR a_28727_39955# 0.355584f
C305 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.271482f
C306 VPWR a_5130_27500# 0.382397f
C307 VPWR a_8822_43816# 0.391817f
C308 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.527529f
C309 VPWR a_18902_41352# 0.394053f
C310 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.930839f
C311 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.107567f
C312 VPWR a_20250_28556# 0.406628f
C313 uo_out[7] uo_out[4] 0.121648f
C314 uo_out[6] uo_out[5] 0.327382f
C315 VPWR uo_out[3] 1.25759f
C316 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.725614f
C317 ua[1] SUNSAR_SAR8B_CV_0.SARN 0.806872f
C318 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H 0.452478f
C319 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.441867f
C320 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C321 VPWR a_5130_34716# 0.399819f
C322 VPWR a_3762_27500# 0.382189f
C323 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN 0.24816f
C324 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.109613f
C325 VPWR a_5130_31196# 0.44007f
C326 VPWR a_18882_28556# 0.406628f
C327 VPWR uo_out[4] 1.03021f
C328 uo_out[7] uo_out[5] 1.57818f
C329 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.106927f
C330 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.722887f
C331 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.11641f
C332 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA6.A 1.63909f
C333 VPWR a_28727_40307# 0.410063f
C334 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.671839f
C335 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.301485f
C336 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.316693f
C337 VPWR a_3762_34716# 0.399819f
C338 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.375025f
C339 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S 0.104609f
C340 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.40569f
C341 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_5648# 0.172147f
C342 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.432466f
C343 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.A 1.2202f
C344 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.109137f
C345 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.CPO 0.131536f
C346 VPWR a_3762_31196# 0.44007f
C347 uo_out[7] uo_out[6] 2.38922f
C348 VPWR uo_out[5] 1.02721f
C349 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.106927f
C350 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.101979f
C351 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.143675f
C352 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.152052f
C353 VPWR a_15210_33836# 0.409601f
C354 VPWR a_10170_29612# 0.397362f
C355 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.55251f
C356 VPWR a_9990_4918# 0.468783f
C357 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN 0.144331f
C358 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.441867f
C359 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.126806f
C360 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.271482f
C361 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN 0.248827f
C362 VPWR a_5150_43816# 0.391817f
C363 VPWR a_15230_41352# 0.394053f
C364 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.16676f
C365 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_42408# 0.100131f
C366 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.93081f
C367 VPWR uo_out[6] 1.34623f
C368 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C369 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.119314f
C370 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.144778f
C371 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.180903f
C372 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.339883f
C373 VPWR a_13842_33836# 0.409601f
C374 VPWR a_8802_29612# 0.397362f
C375 SUNSAR_CAPT8B_CV_0.XF11.QN a_12710_43816# 0.127669f
C376 VPWR tt_um_TT06_SAR_done_0.x3.MP1.G 0.695784f
C377 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_5094# 0.160184f
C378 VPWR a_20250_27852# 0.358413f
C379 VPWR a_3782_43816# 0.391817f
C380 VPWR a_13862_41352# 0.394053f
C381 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C382 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.45828f
C383 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C384 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.A 1.22023f
C385 VPWR a_15210_28556# 0.406628f
C386 VPWR uo_out[7] 1.27659f
C387 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.327152f
C388 VPWR a_23942_42408# 0.3915f
C389 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.728421f
C390 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.139471f
C391 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.B 0.297144f
C392 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.293873f
C393 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA6.A 1.63909f
C394 uio_oe[0] TIE_L1 0.902557f
C395 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_17730_35068# 0.127528f
C396 VPWR a_28727_40659# 0.39147f
C397 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_5094# 0.160184f
C398 SUNSAR_SAR8B_CV_0.XA7.EN a_17730_28556# 0.132757f
C399 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_SAR8B_CV_0.D<5> 0.241356f
C400 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.363295f
C401 VPWR a_23922_34892# 0.395601f
C402 VPWR a_18882_27852# 0.358599f
C403 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN 0.249322f
C404 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.527529f
C405 clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.438597f
C406 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.109613f
C407 VPWR a_23922_31724# 0.412398f
C408 VPWR a_13842_28556# 0.406628f
C409 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.55251f
C410 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C411 VPWR SUNSAR_SAR8B_CV_0.XB2.TIE_L 7.37316f
C412 VPWR a_16542_5270# 0.489055f
C413 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43816# 0.129239f
C414 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.791379f
C415 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.301485f
C416 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S 0.104609f
C417 VPWR SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 11.7505f
C418 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_6608# 0.172147f
C419 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.930839f
C420 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.110962f
C421 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.TIE_L 4.28648f
C422 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.154232f
C423 VPWR a_10170_33836# 0.409601f
C424 VPWR a_5130_29612# 0.397362f
C425 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 3.55251f
C426 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.787331f
C427 VPWR SUNSAR_CAPT8B_CV_0.XA6.A 1.18734f
C428 VPWR tt_um_TT06_SAR_done_0.x4.MP0.G 0.511762f
C429 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B 0.254583f
C430 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_28556# 0.135353f
C431 VPWR SUNSAR_SAR8B_CV_0.XA7.ENO 4.77251f
C432 VPWR a_23942_43992# 0.388156f
C433 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN 0.267395f
C434 VPWR a_10190_41352# 0.394053f
C435 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C436 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 2.62711f
C437 VPWR a_20270_42408# 0.391292f
C438 VPWR a_20250_36828# 0.392512f
C439 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.3401f
C440 VPWR a_8802_33836# 0.409601f
C441 VPWR a_3762_29612# 0.397362f
C442 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN 0.144331f
C443 VPWR a_28727_41011# 0.468616f
C444 VPWR SUNSAR_SAR8B_CV_0.XA7.EN 5.54203f
C445 VPWR a_15210_27852# 0.358413f
C446 VPWR a_8822_41352# 0.394053f
C447 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.432466f
C448 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.A 1.2202f
C449 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C450 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 2.62329f
C451 VPWR a_10170_28556# 0.406628f
C452 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.327909f
C453 VPWR a_18902_42408# 0.391292f
C454 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.B 0.342913f
C455 VPWR a_18882_36828# 0.395703f
C456 VPWR a_9990_5270# 0.490626f
C457 VPWR a_20270_43288# 0.394205f
C458 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.419738f
C459 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_41880# 0.100592f
C460 VPWR SUNSAR_SAR8B_CV_0.XA6.EN 4.84607f
C461 VPWR a_13842_27852# 0.358599f
C462 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN 0.248612f
C463 VPWR SUNSAR_CAPT8B_CV_0.XI14.QN 0.901631f
C464 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.240612f
C465 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.744161f
C466 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.93081f
C467 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 2.62342f
C468 VPWR a_8802_28556# 0.406628f
C469 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 54.2165f
C470 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.793076f
C471 VPWR SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G 0.808658f
C472 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.381914f
C473 VPWR a_18902_43288# 0.394205f
C474 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_16362_35068# 0.129098f
C475 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C476 VPWR a_28727_41363# 0.440399f
C477 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.301485f
C478 VPWR SUNSAR_SAR8B_CV_0.XA5.EN 5.52623f
C479 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.271482f
C480 VPWR SUNSAR_CAPT8B_CV_0.XH13.QN 0.901622f
C481 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C482 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.A 1.22398f
C483 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 2.62342f
C484 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_22790_43640# 0.127669f
C485 VPWR a_5130_33836# 0.409601f
C486 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 54.2173f
C487 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_2982# 0.158066f
C488 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN 0.144331f
C489 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.419738f
C490 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C491 SUNSAR_SAR8B_CV_0.XA5.EN a_12690_28556# 0.132757f
C492 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_5446# 0.102604f
C493 VPWR SUNSAR_SAR8B_CV_0.XA4.EN 4.84607f
C494 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN 0.248535f
C495 VPWR SUNSAR_CAPT8B_CV_0.XG12.QN 0.901622f
C496 VPWR a_5150_41352# 0.394053f
C497 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 2.62342f
C498 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C499 VPWR a_15230_42408# 0.391292f
C500 VPWR a_15210_36828# 0.395582f
C501 VPWR a_3762_33836# 0.409601f
C502 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C503 VPWR a_23942_40296# 0.453754f
C504 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_5446# 0.101033f
C505 VPWR SUNSAR_SAR8B_CV_0.XA3.EN 5.52623f
C506 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S 0.104609f
C507 VPWR a_10170_27852# 0.358413f
C508 VPWR SUNSAR_CAPT8B_CV_0.XF11.QN 0.901622f
C509 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.527529f
C510 VPWR a_3782_41352# 0.394053f
C511 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C512 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.432466f
C513 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.94014f
C514 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.62393f
C515 VPWR a_5130_28556# 0.406628f
C516 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.327152f
C517 VPWR a_13862_42408# 0.391292f
C518 VPWR a_13842_36828# 0.395703f
C519 VPWR a_16542_5622# 0.472384f
C520 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C521 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38576f
C522 VPWR a_15230_43288# 0.394205f
C523 uo_out[5] TIE_L1 0.275794f
C524 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_SAR8B_CV_0.D<6> 0.241356f
C525 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_20270_42760# 0.111734f
C526 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_28556# 0.135353f
C527 VPWR SUNSAR_SAR8B_CV_0.XA2.EN 4.84607f
C528 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.271482f
C529 VPWR a_8802_27852# 0.358599f
C530 VPWR SUNSAR_CAPT8B_CV_0.XE10.QN 0.901622f
C531 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN 0.258218f
C532 VPWR a_23922_35948# 0.390687f
C533 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.62403f
C534 VPWR a_3762_28556# 0.406628f
C535 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 6.86675f
C536 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C537 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA6.EN 1.2771f
C538 VPWR SUNSAR_SAR8B_CV_0.SARN 0.132799f
C539 VPWR a_13862_43288# 0.394205f
C540 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN 0.538639f
C541 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.301485f
C542 VPWR SUNSAR_SAR8B_CV_0.XA1.EN 5.52718f
C543 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.474658f
C544 VPWR SUNSAR_CAPT8B_CV_0.XD09.QN 0.901622f
C545 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.412143f
C546 VPWR SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.635621f
C547 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C548 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.162703f
C549 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.152052f
C550 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 6.86675f
C551 VPWR a_16542_5974# 0.449888f
C552 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.303978f
C553 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_2982# 0.158066f
C554 uo_out[7] TIE_L1 0.206895f
C555 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_12690_35068# 0.127528f
C556 VPWR a_20270_40296# 0.455248f
C557 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.791351f
C558 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C559 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN 0.263255f
C560 VPWR SUNSAR_CAPT8B_CV_0.XC08.QN 0.901622f
C561 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.744161f
C562 VPWR a_20250_32076# 0.433941f
C563 VPWR a_10190_42408# 0.391292f
C564 VPWR a_10170_36828# 0.396003f
C565 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.339883f
C566 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.206292f
C567 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.57155f
C568 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.13078f
C569 VPWR TIE_L1 0.114647f
C570 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN 0.144331f
C571 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C572 VPWR a_18902_40296# 0.457343f
C573 VPWR a_20250_35068# 0.391458f
C574 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S 0.104609f
C575 VPWR a_5130_27852# 0.358413f
C576 VPWR SUNSAR_CAPT8B_CV_0.XB07.QN 0.901622f
C577 VPWR a_20250_35948# 0.414756f
C578 VPWR a_18882_32076# 0.436368f
C579 VPWR a_20250_28908# 0.395394f
C580 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.327909f
C581 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C582 VPWR a_8822_42408# 0.391292f
C583 VPWR a_8802_36828# 0.396052f
C584 VPWR SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.405511f
C585 VPWR SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G 0.808658f
C586 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3334# 0.163985f
C587 VPWR a_10190_43288# 0.394205f
C588 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.449584f
C589 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_18902_42760# 0.113305f
C590 VPWR a_18882_35068# 0.394528f
C591 SUNSAR_SAR8B_CV_0.XA3.EN a_7650_28556# 0.132757f
C592 VPWR a_3762_27852# 0.358599f
C593 VPWR SUNSAR_CAPT8B_CV_0.XA2.MP0.G 0.667429f
C594 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.527529f
C595 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S 0.106927f
C596 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C597 VPWR a_18882_35948# 0.417826f
C598 VPWR a_18882_28908# 0.395394f
C599 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 27.1615f
C600 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.09966f
C601 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA4.EN 1.2771f
C602 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 1.70987f
C603 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.111867f
C604 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.352238f
C605 VPWR a_8822_43288# 0.394205f
C606 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.301485f
C607 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.205884f
C608 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S 0.106927f
C609 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C610 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.17528f
C611 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.154232f
C612 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 27.1625f
C613 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.41635f
C614 VPWR a_9990_5622# 0.470814f
C615 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN 0.144331f
C616 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.449584f
C617 VPWR a_15230_40296# 0.455577f
C618 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.10132f
C619 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.791379f
C620 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_SAR8B_CV_0.D<7> 0.241356f
C621 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_28556# 0.135353f
C622 VPWR a_20270_44168# 0.340085f
C623 VPWR SUNSAR_SAR8B_CV_0.D<1> 5.18522f
C624 VPWR a_15210_32076# 0.436368f
C625 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.297363f
C626 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.449584f
C627 VPWR a_5150_42408# 0.391292f
C628 VPWR a_5130_36828# 0.395767f
C629 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.3401f
C630 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.182408f
C631 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.143554f
C632 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_11322_35068# 0.129098f
C633 VPWR a_13862_40296# 0.457343f
C634 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.34399f
C635 VPWR a_15210_35068# 0.394528f
C636 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.271482f
C637 VPWR a_18902_44168# 0.3405f
C638 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C639 VPWR a_15210_35948# 0.417826f
C640 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C641 VPWR a_13842_32076# 0.436368f
C642 VPWR a_15210_28908# 0.395394f
C643 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.19724f
C644 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C645 VPWR a_16542_2630# 0.448659f
C646 VPWR a_3782_42408# 0.391292f
C647 VPWR a_3762_36828# 0.395857f
C648 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.103734f
C649 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 4.36162f
C650 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.291229f
C651 VPWR a_9990_5974# 0.451043f
C652 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3686# 0.16579f
C653 VPWR a_5150_43288# 0.394205f
C654 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3334# 0.163985f
C655 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.193518f
C656 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_41880# 0.100592f
C657 VPWR a_13842_35068# 0.394528f
C658 VPWR a_13842_35948# 0.417826f
C659 VPWR a_13842_28908# 0.395394f
C660 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6519f
C661 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80606f
C662 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.449584f
C663 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA2.EN 1.2771f
C664 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S 0.152518f
C665 VPWR a_23922_34540# 0.502044f
C666 VPWR a_23922_26796# 0.442318f
C667 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA7.EN 0.438277f
C668 VPWR a_3782_43288# 0.394205f
C669 uo_out[7] TIE_L2 0.100011f
C670 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.238862f
C671 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.301485f
C672 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S 0.104609f
C673 uio_out[0] TIE_L 0.44106f
C674 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.205884f
C675 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.625035f
C676 VPWR SUNSAR_SAR8B_CV_0.D<2> 5.20829f
C677 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.665724f
C678 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C679 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.686731f
C680 VPWR SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.714341f
C681 SUNSAR_CAPT8B_CV_0.XA5.XA2.A a_22790_42408# 0.10248f
C682 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 13.6523f
C683 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.303978f
C684 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.305166f
C685 VPWR a_10190_40296# 0.455675f
C686 SUNSAR_SAR8B_CV_0.XA1.EN a_2610_28556# 0.132757f
C687 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_15230_42760# 0.111734f
C688 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.271482f
C689 uio_oe[0] TIE_L 1.21913f
C690 VPWR a_15230_44168# 0.340085f
C691 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S 0.106927f
C692 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.A 0.744161f
C693 VPWR a_10170_32076# 0.436368f
C694 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.898003f
C695 VPWR SUNSAR_SAR8B_CV_0.XA20.CK_CMP 1.1111f
C696 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S 0.150467f
C697 SUNSAR_SAR8B_CV_0.XA7.XA12.A a_21402_36828# 0.104051f
C698 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.13078f
C699 VPWR a_8822_40296# 0.457343f
C700 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.107823f
C701 VPWR a_10170_35068# 0.394528f
C702 VPWR a_13862_44168# 0.3405f
C703 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S 0.106927f
C704 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C705 VPWR a_10170_35948# 0.417826f
C706 VPWR a_8802_32076# 0.436368f
C707 VPWR a_10170_28908# 0.395394f
C708 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.34383f
C709 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.898003f
C710 VPWR SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.723713f
C711 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_21422_42408# 0.113479f
C712 VPWR a_20250_26796# 0.441753f
C713 ui_in[0] tt_um_TT06_SAR_done_0.DONE 0.198829f
C714 VPWR SUNSAR_CAPT8B_CV_0.XA6.B 0.86364f
C715 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3686# 0.16579f
C716 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.145738f
C717 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_7650_35068# 0.127528f
C718 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C719 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN 0.253395f
C720 VPWR a_8802_35068# 0.394528f
C721 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.143023f
C722 clk TIE_L 0.146712f
C723 VPWR SUNSAR_SAR8B_CV_0.D<3> 5.17056f
C724 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.11536f
C725 VPWR a_8802_35948# 0.417826f
C726 VPWR a_8802_28908# 0.395394f
C727 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.55251f
C728 VPWR a_9990_2630# 0.447504f
C729 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.39041f
C730 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.898003f
C731 VPWR SUNSAR_SAR8B_CV_0.XA7.CEIN 2.28789f
C732 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C733 VPWR a_18882_26796# 0.442908f
C734 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.352238f
C735 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA6.EN 0.503825f
C736 VPWR a_23942_43640# 0.412992f
C737 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C738 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.301485f
C739 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S 0.104609f
C740 uo_out[0] TIE_L 0.280844f
C741 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.205884f
C742 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 0.625175f
C743 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C744 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.A 0.504864f
C745 ua[0] SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.241597f
C746 VPWR a_16542_2982# 0.490338f
C747 SUNSAR_SAR8B_CV_0.XA7.XA11.A a_21402_36300# 0.13402f
C748 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C749 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.898003f
C750 VPWR SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.720096f
C751 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.152052f
C752 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.104122f
C753 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S 0.112098f
C754 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 3.57448f
C755 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 0.305131f
C756 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_21402_35420# 0.160931f
C757 VPWR a_5150_40296# 0.455605f
C758 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.40569f
C759 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.791351f
C760 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_13862_42760# 0.113305f
C761 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.142977f
C762 VPWR a_10190_44168# 0.340085f
C763 uo_out[1] TIE_L 0.50141f
C764 VPWR a_5130_32076# 0.436368f
C765 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.100365f
C766 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.898003f
C767 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C768 VPWR SUNSAR_SAR8B_CV_0.XA6.CEIN 1.0603f
C769 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.280191f
C770 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.339883f
C771 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S 0.155821f
C772 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S 0.112858f
C773 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_20250_35420# 0.133834f
C774 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.143554f
C775 VPWR a_3782_40296# 0.457343f
C776 VPWR a_5130_35068# 0.394528f
C777 VPWR a_8822_44168# 0.3405f
C778 uo_out[2] TIE_L 0.156661f
C779 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C780 VPWR SUNSAR_SAR8B_CV_0.D<4> 5.15123f
C781 VPWR a_5130_35948# 0.417826f
C782 VPWR a_3762_32076# 0.436368f
C783 VPWR a_5130_28908# 0.395394f
C784 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.55251f
C785 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189112f
C786 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C787 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.898003f
C788 VPWR SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.723728f
C789 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.152045f
C790 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_17750_42408# 0.111909f
C791 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 4.24834f
C792 VPWR a_15210_26796# 0.441753f
C793 SUNSAR_SAR8B_CV_0.XA6.XA12.A a_17730_36828# 0.10248f
C794 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S 0.106927f
C795 VPWR a_3762_35068# 0.394528f
C796 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.142956f
C797 uo_out[3] TIE_L 0.185333f
C798 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.137975f
C799 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S 0.106927f
C800 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.A 0.744161f
C801 VPWR a_3762_35948# 0.417826f
C802 VPWR a_3762_28908# 0.395394f
C803 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.898003f
C804 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C805 VPWR SUNSAR_SAR8B_CV_0.XA5.CEIN 2.30385f
C806 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C807 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S 0.150467f
C808 VPWR a_13842_26796# 0.442908f
C809 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA5.EN 0.438277f
C810 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_6282_35068# 0.129098f
C811 VPWR a_23942_40648# 0.489579f
C812 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C813 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.301485f
C814 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.271482f
C815 uo_out[4] TIE_L 0.31941f
C816 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.625035f
C817 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.205884f
C818 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S 0.106927f
C819 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.618979f
C820 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.100365f
C821 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.898003f
C822 VPWR SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.720133f
C823 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.154232f
C824 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_16382_42408# 0.113479f
C825 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.303978f
C826 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 1.77563f
C827 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_18882_35420# 0.133834f
C828 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 3.86364f
C829 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.142977f
C830 VPWR a_5150_44168# 0.340085f
C831 uo_out[5] TIE_L 1.3092f
C832 VPWR SUNSAR_SAR8B_CV_0.D<5> 5.14531f
C833 VPWR SUNSAR_SAR8B_CV_0.XA20.XA12.Y 1.13456f
C834 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.324111f
C835 VPWR a_9990_2982# 0.491909f
C836 VPWR a_23942_42760# 0.388156f
C837 VPWR SUNSAR_SAR8B_CV_0.XA4.CEIN 1.06031f
C838 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.3401f
C839 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C840 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 4.25569f
C841 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.13078f
C842 SUNSAR_SAR8B_CV_0.XA5.XA12.A a_16362_36828# 0.104051f
C843 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S 0.106927f
C844 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_17730_35420# 0.160931f
C845 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 0.635098f
C846 SUNSAR_CAPT8B_CV_0.XA5.B a_22790_41000# 0.11811f
C847 VPWR a_3782_44168# 0.3405f
C848 uo_out[6] TIE_L 0.204625f
C849 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.105016f
C850 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.174995f
C851 VPWR SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.774301f
C852 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S 0.104609f
C853 VPWR a_16542_3334# 0.380282f
C854 SUNSAR_SAR8B_CV_0.XA6.XA11.A a_17730_36300# 0.13253f
C855 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C856 VPWR SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.723762f
C857 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.104122f
C858 VPWR a_10170_26796# 0.441753f
C859 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 0.305131f
C860 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.145738f
C861 VPWR a_20270_40648# 0.492579f
C862 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_10190_42760# 0.111734f
C863 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_41880# 0.100592f
C864 VPWR SUNSAR_SAR8B_CV_0.XA6.DONE 0.246222f
C865 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.142956f
C866 VPWR a_20250_30316# 0.403745f
C867 uo_out[7] TIE_L 0.471918f
C868 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.475004f
C869 VPWR SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.780003f
C870 tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G 0.186749f
C871 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.2165f
C872 VPWR SUNSAR_SAR8B_CV_0.XA3.CEIN 2.30393f
C873 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.300065f
C874 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S 0.155821f
C875 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.352238f
C876 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA4.EN 0.503825f
C877 VPWR a_8802_26796# 0.442908f
C878 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 1.77562f
C879 VPWR a_18902_40648# 0.491225f
C880 VPWR SUNSAR_SAR8B_CV_0.XA5.DONE 0.245452f
C881 VPWR a_18882_30316# 0.403802f
C882 VPWR TIE_L 0.387688f
C883 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.205884f
C884 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 0.625175f
C885 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.419738f
C886 VPWR SUNSAR_SAR8B_CV_0.D<6> 5.17441f
C887 VPWR SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.779986f
C888 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S 0.104609f
C889 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.10225f
C890 SUNSAR_SAR8B_CV_0.XA5.XA11.A a_16362_36300# 0.13402f
C891 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C892 VPWR a_20270_42760# 0.391454f
C893 VPWR SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.720114f
C894 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_12710_42408# 0.111909f
C895 VPWR tt_um_TT06_SAR_done_0.DONE 8.46867f
C896 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S 0.101001f
C897 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_2610_35068# 0.127528f
C898 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C899 VPWR SUNSAR_SAR8B_CV_0.XA4.DONE 0.246222f
C900 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.142977f
C901 VPWR a_23942_44344# 0.342053f
C902 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.11099f
C903 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S 0.106927f
C904 VPWR SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.780003f
C905 VPWR a_18902_42760# 0.391454f
C906 VPWR SUNSAR_SAR8B_CV_0.XA2.CEIN 1.0603f
C907 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C908 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S 0.150467f
C909 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.143554f
C910 VPWR SUNSAR_SAR8B_CV_0.XA3.DONE 0.245452f
C911 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87301f
C912 VPWR a_20250_28204# 0.361706f
C913 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.419738f
C914 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S 0.106927f
C915 VPWR SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.779986f
C916 VPWR SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.728492f
C917 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.26609f
C918 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_11342_42408# 0.113479f
C919 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S 0.112858f
C920 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.386305f
C921 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.215804f
C922 SUNSAR_SAR8B_CV_0.XA4.XA12.A a_12690_36828# 0.10248f
C923 VPWR a_5130_26796# 0.441753f
C924 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S 0.106927f
C925 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.309657f
C926 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_16362_35420# 0.160931f
C927 VPWR a_15230_40648# 0.492579f
C928 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_8822_42760# 0.113305f
C929 VPWR SUNSAR_SAR8B_CV_0.XA2.DONE 0.246222f
C930 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.142956f
C931 VPWR a_15210_30316# 0.404384f
C932 VPWR a_18882_28204# 0.36179f
C933 VPWR SUNSAR_SAR8B_CV_0.D<7> 3.61291f
C934 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.744161f
C935 VPWR SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.780003f
C936 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.86675f
C937 VPWR a_9990_3334# 0.380282f
C938 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.155424f
C939 VPWR SUNSAR_SAR8B_CV_0.XA1.CEIN 2.30575f
C940 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C941 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S 0.112858f
C942 VPWR a_3762_26796# 0.442908f
C943 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA3.EN 0.434116f
C944 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_15210_35420# 0.133834f
C945 VPWR a_13862_40648# 0.491225f
C946 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_42408# 0.100131f
C947 VPWR SUNSAR_SAR8B_CV_0.XA1.DONE 0.245452f
C948 VPWR a_13842_30316# 0.404384f
C949 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.205884f
C950 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.08082f
C951 VPWR SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.779986f
C952 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C953 VPWR a_15230_42760# 0.391454f
C954 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.152052f
C955 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.473354f
C956 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.104122f
C957 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 4.2492f
C958 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 1.77562f
C959 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 4.0111f
C960 VPWR SUNSAR_SAR8B_CV_0.XA0.DONE 0.247527f
C961 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.433299f
C962 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.142977f
C963 VPWR a_23942_41880# 0.398828f
C964 VPWR SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.784656f
C965 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S 0.104609f
C966 VPWR a_13862_42760# 0.391454f
C967 VPWR a_20250_37180# 0.469114f
C968 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.149144f
C969 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145339f
C970 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S 0.155821f
C971 VPWR a_23922_27148# 0.483246f
C972 SUNSAR_SAR8B_CV_0.XA3.XA12.A a_11322_36828# 0.104051f
C973 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S 0.106927f
C974 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.437693f
C975 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C976 VPWR a_23922_35420# 0.416528f
C977 VPWR a_15210_28204# 0.361706f
C978 VPWR a_23922_36300# 0.472384f
C979 VPWR SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 1.56028f
C980 SUNSAR_SAR8B_CV_0.XA4.XA11.A a_12690_36300# 0.13253f
C981 VPWR a_18882_37180# 0.473682f
C982 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_7670_42408# 0.111909f
C983 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.182595f
C984 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.101001f
C985 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_13842_35420# 0.133834f
C986 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C987 VPWR a_10190_40648# 0.492624f
C988 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.2199f
C989 VPWR a_10170_30316# 0.404384f
C990 VPWR a_13842_28204# 0.36179f
C991 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.199516f
C992 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1615f
C993 VPWR SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.183853f
C994 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C995 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S 0.150467f
C996 SUNSAR_CAPT8B_CV_0.XA6.A a_22790_41880# 0.111538f
C997 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 4.27988f
C998 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA2.EN 0.491653f
C999 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 1.77562f
C1000 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_12690_35420# 0.160931f
C1001 VPWR a_8822_40648# 0.491225f
C1002 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.398331f
C1003 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.134182f
C1004 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.98135f
C1005 VPWR a_8802_30316# 0.404384f
C1006 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.20727f
C1007 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.205884f
C1008 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C1009 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.449584f
C1010 VPWR a_20270_41880# 0.395781f
C1011 VPWR a_20250_32956# 0.433941f
C1012 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S 0.104609f
C1013 SUNSAR_SAR8B_CV_0.XA3.XA11.A a_11322_36300# 0.13402f
C1014 VPWR a_10190_42760# 0.391454f
C1015 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_6302_42408# 0.113479f
C1016 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.375196f
C1017 VPWR a_20250_27148# 0.470364f
C1018 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.324105f
C1019 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.305131f
C1020 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.437693f
C1021 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.25689f
C1022 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_5150_42760# 0.111734f
C1023 VPWR a_20250_35420# 0.39661f
C1024 VPWR a_18902_41880# 0.395781f
C1025 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.744161f
C1026 VPWR a_20250_36300# 0.395776f
C1027 VPWR a_18882_32956# 0.436368f
C1028 VPWR SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.183853f
C1029 VPWR a_8822_42760# 0.391454f
C1030 VPWR a_15210_37180# 0.474036f
C1031 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C1032 VPWR a_18882_27148# 0.471462f
C1033 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.138f
C1034 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C1035 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.79343f
C1036 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C1037 VPWR a_18882_35420# 0.39968f
C1038 VPWR a_10170_28204# 0.361706f
C1039 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.178111f
C1040 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.449584f
C1041 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.174995f
C1042 VPWR a_18882_36300# 0.399161f
C1043 VPWR a_16542_4038# 0.379979f
C1044 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.765539f
C1045 TIE_L TIE_L1 0.257793f
C1046 VPWR a_13842_37180# 0.473697f
C1047 SUNSAR_SAR8B_CV_0.XA2.XA12.A a_7650_36828# 0.10248f
C1048 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.158152f
C1049 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S 0.106927f
C1050 VPWR a_5150_40648# 0.492592f
C1051 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233744f
C1052 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C1053 VPWR a_5130_30316# 0.404384f
C1054 VPWR a_8802_28204# 0.36179f
C1055 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.50324f
C1056 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6519f
C1057 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.4271f
C1058 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C1059 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.303428f
C1060 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.383512f
C1061 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA1.EN 0.11341f
C1062 VPWR a_3782_40648# 0.491225f
C1063 VPWR a_3762_30316# 0.404384f
C1064 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C1065 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.205884f
C1066 VPWR a_15230_41880# 0.395781f
C1067 VPWR a_15210_32956# 0.436368f
C1068 VPWR a_5150_42760# 0.391454f
C1069 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.244517f
C1070 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_2630_42408# 0.111909f
C1071 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S 0.112858f
C1072 VPWR a_15210_27148# 0.470364f
C1073 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.220689f
C1074 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.30523f
C1075 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 1.77562f
C1076 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.224309f
C1077 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.527529f
C1078 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_11322_35420# 0.160931f
C1079 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.394834f
C1080 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_3782_42760# 0.113305f
C1081 VPWR a_15210_35420# 0.39968f
C1082 VPWR a_13862_41880# 0.395781f
C1083 VPWR a_15210_36300# 0.398846f
C1084 VPWR a_13842_32956# 0.436368f
C1085 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S 0.104609f
C1086 VPWR a_3782_42760# 0.391454f
C1087 VPWR a_10170_37180# 0.474068f
C1088 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C1089 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_SAR8B_CV_0.D<1> 0.241356f
C1090 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S 0.112858f
C1091 VPWR a_13842_27148# 0.471462f
C1092 SUNSAR_SAR8B_CV_0.XA1.XA12.A a_6282_36828# 0.104051f
C1093 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S 0.106927f
C1094 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_10170_35420# 0.133834f
C1095 VPWR a_13842_35420# 0.39968f
C1096 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.07223f
C1097 VPWR SUNSAR_SAR8B_CV_0.XA20.CPO 6.88568f
C1098 VPWR a_5130_28204# 0.361706f
C1099 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C1100 ui_in[0] SUNSAR_CAPT8B_CV_0.XA5.B 0.172623f
C1101 VPWR a_13842_36300# 0.399161f
C1102 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.762388f
C1103 SUNSAR_SAR8B_CV_0.XA2.XA11.A a_7650_36300# 0.13253f
C1104 VPWR a_8802_37180# 0.473729f
C1105 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.18614f
C1106 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<1> 0.297507f
C1107 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 4.24508f
C1108 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.377598f
C1109 VPWR a_23942_41000# 0.390551f
C1110 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C1111 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 5.19722f
C1112 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.432466f
C1113 VPWR a_23922_30844# 0.425847f
C1114 VPWR a_3762_28204# 0.36179f
C1115 ua[1] ua[0] 3.85017f
C1116 clk SUNSAR_CAPT8B_CV_0.XA5.B 0.210661f
C1117 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.55251f
C1118 VPWR a_9990_4038# 0.379979f
C1119 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.127551f
C1120 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.145048f
C1121 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA20.CPO 0.328435f
C1122 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 1.77562f
C1123 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_42408# 0.100131f
C1124 VPWR a_10190_41880# 0.395781f
C1125 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C1126 VPWR a_10170_32956# 0.436368f
C1127 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S 0.104609f
C1128 SUNSAR_SAR8B_CV_0.XA1.XA11.A a_6282_36300# 0.13402f
C1129 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.693521f
C1130 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.293159f
C1131 VPWR a_10170_27148# 0.470364f
C1132 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_8802_35420# 0.133834f
C1133 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C1134 VPWR a_10170_35420# 0.39968f
C1135 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C1136 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.429492f
C1137 VPWR a_8822_41880# 0.395781f
C1138 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.744161f
C1139 VPWR a_10170_36300# 0.398846f
C1140 VPWR a_8802_32956# 0.436368f
C1141 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31666f
C1142 VPWR a_23942_43112# 0.393308f
C1143 VPWR a_5130_37180# 0.474051f
C1144 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C1145 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.D<2> 0.297715f
C1146 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 4.25322f
C1147 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA6.CEIN 0.432008f
C1148 VPWR a_8802_27148# 0.471462f
C1149 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.527529f
C1150 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_7650_35420# 0.160931f
C1151 VPWR a_20270_41000# 0.388156f
C1152 VPWR a_8802_35420# 0.39968f
C1153 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S 0.137646f
C1154 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C1155 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C1156 ua[2] VGND 0.117454f
C1157 ua[3] VGND 0.117454f
C1158 ua[4] VGND 0.118698f
C1159 ua[5] VGND 0.120088f
C1160 ua[6] VGND 0.120088f
C1161 ua[7] VGND 0.111009f
C1162 ua[0] VGND 9.399512f
C1163 ua[1] VGND 8.540812f
C1164 uio_out[0] VGND 8.52142f
C1165 uio_oe[0] VGND 7.87718f
C1166 ui_in[0] VGND 5.40407f
C1167 clk VGND 6.22723f
C1168 uo_out[0] VGND 2.40292f
C1169 uo_out[1] VGND 1.50319f
C1170 uo_out[2] VGND 1.42895f
C1171 uo_out[3] VGND 1.68048f
C1172 uo_out[4] VGND 1.55276f
C1173 uo_out[5] VGND 1.75883f
C1174 uo_out[6] VGND 3.667369f
C1175 uo_out[7] VGND 4.218073f
C1176 VPWR VGND 0.515222p
C1177 TIE_L1 VGND 1.33691f
C1178 TIE_L2 VGND 1.67804f
C1179 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93609f
C1180 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93609f
C1181 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.5533f
C1182 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.5533f
C1183 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.334839f
C1184 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.334839f
C1185 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.469f
C1186 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.469f
C1187 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43533f
C1188 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43533f
C1189 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67745f
C1190 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67745f
C1191 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.6684f
C1192 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.6684f
C1193 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.574499f
C1194 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.574499f
C1195 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33412f
C1196 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33412f
C1197 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.469f
C1198 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.469f
C1199 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43533f
C1200 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43533f
C1201 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67745f
C1202 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67745f
C1203 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.6684f
C1204 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.6684f
C1205 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.575099f
C1206 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.575099f
C1207 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33412f
C1208 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33412f
C1209 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.469f
C1210 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.469f
C1211 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43533f
C1212 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43533f
C1213 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67745f
C1214 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67745f
C1215 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.6684f
C1216 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.6684f
C1217 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.571799f
C1218 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.571799f
C1219 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33412f
C1220 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33412f
C1221 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.471901f
C1222 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.471901f
C1223 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.439809f
C1224 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44253f
C1225 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.3859f
C1226 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.38266f
C1227 a_15390_2630# VGND 0.542161f $ **FLOATING
C1228 a_13950_2630# VGND 0.427094f $ **FLOATING
C1229 a_12582_2630# VGND 0.426679f $ **FLOATING
C1230 a_11142_2630# VGND 0.543317f $ **FLOATING
C1231 a_15390_2982# VGND 0.491607f $ **FLOATING
C1232 a_13950_2982# VGND 0.352472f $ **FLOATING
C1233 a_12582_2982# VGND 0.352472f $ **FLOATING
C1234 a_11142_2982# VGND 0.490037f $ **FLOATING
C1235 a_15390_3334# VGND 0.374919f $ **FLOATING
C1236 a_13950_3334# VGND 0.352438f $ **FLOATING
C1237 a_12582_3334# VGND 0.352438f $ **FLOATING
C1238 a_11142_3334# VGND 0.374919f $ **FLOATING
C1239 a_13950_3686# VGND 0.352418f $ **FLOATING
C1240 a_12582_3686# VGND 0.352418f $ **FLOATING
C1241 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND 41.5268f
C1242 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.70146f
C1243 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.70146f
C1244 a_15390_4038# VGND 0.397033f $ **FLOATING
C1245 a_13950_4038# VGND 0.354407f $ **FLOATING
C1246 a_12582_4038# VGND 0.354407f $ **FLOATING
C1247 a_11142_4038# VGND 0.397033f $ **FLOATING
C1248 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND 0.103625f
C1249 a_13950_4390# VGND 0.352432f $ **FLOATING
C1250 a_12582_4390# VGND 0.352432f $ **FLOATING
C1251 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND 0.103625f
C1252 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VGND 3.1165f
C1253 a_15390_4566# VGND 0.389036f $ **FLOATING
C1254 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VGND 3.07938f
C1255 a_11142_4566# VGND 0.389036f $ **FLOATING
C1256 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VGND 0.970036f
C1257 a_13950_4742# VGND 0.352456f $ **FLOATING
C1258 a_12582_4742# VGND 0.352456f $ **FLOATING
C1259 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND 0.7964f
C1260 a_15390_4918# VGND 0.470144f $ **FLOATING
C1261 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND 0.7964f
C1262 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VGND 0.970036f
C1263 a_11142_4918# VGND 0.471715f $ **FLOATING
C1264 a_13950_5094# VGND 0.353103f $ **FLOATING
C1265 a_12582_5094# VGND 0.353103f $ **FLOATING
C1266 a_15390_5270# VGND 0.492927f $ **FLOATING
C1267 a_11142_5270# VGND 0.491356f $ **FLOATING
C1268 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND 0.596866f
C1269 a_13950_5446# VGND 0.433341f $ **FLOATING
C1270 a_12582_5446# VGND 0.433756f $ **FLOATING
C1271 a_15390_5622# VGND 0.47219f $ **FLOATING
C1272 a_15390_5974# VGND 0.541341f $ **FLOATING
C1273 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND 0.596866f
C1274 a_11142_5622# VGND 0.47376f $ **FLOATING
C1275 a_11142_5974# VGND 0.540186f $ **FLOATING
C1276 a_22770_26796# VGND 0.529341f $ **FLOATING
C1277 a_21402_26796# VGND 0.531659f $ **FLOATING
C1278 a_17730_26796# VGND 0.530834f $ **FLOATING
C1279 a_16362_26796# VGND 0.531989f $ **FLOATING
C1280 a_12690_26796# VGND 0.530834f $ **FLOATING
C1281 a_11322_26796# VGND 0.531989f $ **FLOATING
C1282 a_7650_26796# VGND 0.530213f $ **FLOATING
C1283 a_6282_26796# VGND 0.530979f $ **FLOATING
C1284 a_2610_26796# VGND 0.531178f $ **FLOATING
C1285 a_22770_27148# VGND 0.499848f $ **FLOATING
C1286 a_21402_27148# VGND 0.467094f $ **FLOATING
C1287 a_17730_27148# VGND 0.471508f $ **FLOATING
C1288 a_16362_27148# VGND 0.467722f $ **FLOATING
C1289 a_12690_27148# VGND 0.471508f $ **FLOATING
C1290 a_11322_27148# VGND 0.467722f $ **FLOATING
C1291 a_7650_27148# VGND 0.470266f $ **FLOATING
C1292 a_6282_27148# VGND 0.465734f $ **FLOATING
C1293 a_2610_27148# VGND 0.47123f $ **FLOATING
C1294 a_21402_27500# VGND 0.385968f $ **FLOATING
C1295 a_17730_27500# VGND 0.387712f $ **FLOATING
C1296 a_16362_27500# VGND 0.386249f $ **FLOATING
C1297 a_12690_27500# VGND 0.387712f $ **FLOATING
C1298 a_11322_27500# VGND 0.386249f $ **FLOATING
C1299 a_7650_27500# VGND 0.38671f $ **FLOATING
C1300 a_6282_27500# VGND 0.384229f $ **FLOATING
C1301 a_2610_27500# VGND 0.387675f $ **FLOATING
C1302 a_21402_27852# VGND 0.370125f $ **FLOATING
C1303 a_17730_27852# VGND 0.370785f $ **FLOATING
C1304 a_16362_27852# VGND 0.368771f $ **FLOATING
C1305 a_12690_27852# VGND 0.370785f $ **FLOATING
C1306 a_11322_27852# VGND 0.368771f $ **FLOATING
C1307 a_7650_27852# VGND 0.369543f $ **FLOATING
C1308 a_6282_27852# VGND 0.366751f $ **FLOATING
C1309 a_2610_27852# VGND 0.370508f $ **FLOATING
C1310 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND 0.506947f
C1311 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND 0.502211f
C1312 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND 0.477244f
C1313 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND 0.502211f
C1314 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND 0.477244f
C1315 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND 0.502211f
C1316 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND 0.477244f
C1317 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND 0.502211f
C1318 a_21402_28204# VGND 0.405715f $ **FLOATING
C1319 a_17730_28204# VGND 0.406284f $ **FLOATING
C1320 a_16362_28204# VGND 0.406284f $ **FLOATING
C1321 a_12690_28204# VGND 0.406284f $ **FLOATING
C1322 a_11322_28204# VGND 0.406284f $ **FLOATING
C1323 a_7650_28204# VGND 0.405133f $ **FLOATING
C1324 a_6282_28204# VGND 0.404355f $ **FLOATING
C1325 a_2610_28204# VGND 0.406098f $ **FLOATING
C1326 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND 0.608956f
C1327 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND 0.741242f
C1328 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND 0.749251f
C1329 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND 0.735502f
C1330 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND 0.749251f
C1331 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND 0.735502f
C1332 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND 0.746591f
C1333 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND 0.73057f
C1334 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND 0.74895f
C1335 a_22770_28556# VGND 0.401649f $ **FLOATING
C1336 a_21402_28556# VGND 0.387558f $ **FLOATING
C1337 a_17730_28556# VGND 0.388127f $ **FLOATING
C1338 a_16362_28556# VGND 0.388127f $ **FLOATING
C1339 a_12690_28556# VGND 0.388127f $ **FLOATING
C1340 a_11322_28556# VGND 0.388127f $ **FLOATING
C1341 a_7650_28556# VGND 0.386976f $ **FLOATING
C1342 a_6282_28556# VGND 0.386198f $ **FLOATING
C1343 a_2610_28556# VGND 0.38794f $ **FLOATING
C1344 a_21402_28908# VGND 0.394283f $ **FLOATING
C1345 a_17730_28908# VGND 0.394852f $ **FLOATING
C1346 a_16362_28908# VGND 0.394852f $ **FLOATING
C1347 a_12690_28908# VGND 0.394852f $ **FLOATING
C1348 a_11322_28908# VGND 0.394852f $ **FLOATING
C1349 a_7650_28908# VGND 0.393701f $ **FLOATING
C1350 a_6282_28908# VGND 0.392923f $ **FLOATING
C1351 a_2610_28908# VGND 0.394666f $ **FLOATING
C1352 a_21402_29612# VGND 0.395457f $ **FLOATING
C1353 a_17730_29612# VGND 0.396116f $ **FLOATING
C1354 a_16362_29612# VGND 0.395588f $ **FLOATING
C1355 a_12690_29612# VGND 0.396116f $ **FLOATING
C1356 a_11322_29612# VGND 0.395588f $ **FLOATING
C1357 a_7650_29612# VGND 0.394965f $ **FLOATING
C1358 a_6282_29612# VGND 0.393746f $ **FLOATING
C1359 a_2610_29612# VGND 0.395923f $ **FLOATING
C1360 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318647f
C1361 a_22770_29964# VGND 0.400512f $ **FLOATING
C1362 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND 0.103281f
C1363 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N VGND 1.27143f
C1364 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND 0.100021f
C1365 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N VGND 1.26503f
C1366 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND 0.100021f
C1367 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N VGND 1.26391f
C1368 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND 0.100021f
C1369 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N VGND 1.26503f
C1370 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND 0.100021f
C1371 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N VGND 1.26391f
C1372 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND 0.100021f
C1373 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N VGND 1.25938f
C1374 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND 0.100021f
C1375 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N VGND 1.25329f
C1376 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND 0.100021f
C1377 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N VGND 1.26407f
C1378 a_21402_30316# VGND 0.401758f $ **FLOATING
C1379 a_17730_30316# VGND 0.401074f $ **FLOATING
C1380 a_16362_30316# VGND 0.401074f $ **FLOATING
C1381 a_12690_30316# VGND 0.401074f $ **FLOATING
C1382 a_11322_30316# VGND 0.401074f $ **FLOATING
C1383 a_7650_30316# VGND 0.399923f $ **FLOATING
C1384 a_6282_30316# VGND 0.399145f $ **FLOATING
C1385 a_2610_30316# VGND 0.400881f $ **FLOATING
C1386 SUNSAR_SAR8B_CV_0.XA20.CPO VGND 18.232008f
C1387 a_22770_30844# VGND 0.421853f $ **FLOATING
C1388 a_21402_31196# VGND 0.4255f $ **FLOATING
C1389 a_17730_31196# VGND 0.426069f $ **FLOATING
C1390 a_16362_31196# VGND 0.426069f $ **FLOATING
C1391 a_12690_31196# VGND 0.426069f $ **FLOATING
C1392 a_11322_31196# VGND 0.426069f $ **FLOATING
C1393 a_7650_31196# VGND 0.424917f $ **FLOATING
C1394 a_6282_31196# VGND 0.42414f $ **FLOATING
C1395 a_2610_31196# VGND 0.425876f $ **FLOATING
C1396 a_22770_31724# VGND 0.423601f $ **FLOATING
C1397 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 3.362181f
C1398 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 3.414612f
C1399 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 3.341801f
C1400 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 3.414612f
C1401 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 3.341801f
C1402 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 9.493475f
C1403 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.903188f
C1404 a_21402_32076# VGND 0.426091f $ **FLOATING
C1405 a_17730_32076# VGND 0.42666f $ **FLOATING
C1406 a_16362_32076# VGND 0.42666f $ **FLOATING
C1407 a_12690_32076# VGND 0.42666f $ **FLOATING
C1408 a_11322_32076# VGND 0.42666f $ **FLOATING
C1409 a_7650_32076# VGND 0.42666f $ **FLOATING
C1410 a_6282_32076# VGND 0.42666f $ **FLOATING
C1411 a_2610_32076# VGND 0.426468f $ **FLOATING
C1412 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND 1.55564f
C1413 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C1414 a_21402_32956# VGND 0.426069f $ **FLOATING
C1415 a_17730_32956# VGND 0.426069f $ **FLOATING
C1416 a_16362_32956# VGND 0.426069f $ **FLOATING
C1417 a_12690_32956# VGND 0.426069f $ **FLOATING
C1418 a_11322_32956# VGND 0.426069f $ **FLOATING
C1419 a_7650_32956# VGND 0.426069f $ **FLOATING
C1420 a_6282_32956# VGND 0.426069f $ **FLOATING
C1421 a_2610_32956# VGND 0.425876f $ **FLOATING
C1422 a_22770_33132# VGND 0.403395f $ **FLOATING
C1423 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 3.39445f
C1424 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.477508f
C1425 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.385042f
C1426 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.477508f
C1427 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.385042f
C1428 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 11.707785f
C1429 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 12.318709f
C1430 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 18.293753f
C1431 a_21402_33836# VGND 0.426756f $ **FLOATING
C1432 a_17730_33836# VGND 0.426756f $ **FLOATING
C1433 a_16362_33836# VGND 0.426756f $ **FLOATING
C1434 a_12690_33836# VGND 0.426756f $ **FLOATING
C1435 a_11322_33836# VGND 0.426756f $ **FLOATING
C1436 a_7650_33836# VGND 0.426756f $ **FLOATING
C1437 a_6282_33836# VGND 0.426756f $ **FLOATING
C1438 a_2610_33836# VGND 0.426472f $ **FLOATING
C1439 SUNSAR_SAR8B_CV_0.SARN VGND 71.1589f
C1440 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND 0.149691f
C1441 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND 0.515385f
C1442 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C1443 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND 0.149691f
C1444 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 10.934954f
C1445 a_22770_34540# VGND 0.39377f $ **FLOATING
C1446 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND 0.102f
C1447 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND 0.149691f
C1448 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 10.467578f
C1449 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND 0.149691f
C1450 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 9.520044f
C1451 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND 0.102f
C1452 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND 0.102f
C1453 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND 0.149691f
C1454 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 10.720038f
C1455 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND 0.149691f
C1456 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 11.337016f
C1457 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND 0.102f
C1458 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND 0.102f
C1459 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND 0.149691f
C1460 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 13.150025f
C1461 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND 0.149691f
C1462 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 16.484587f
C1463 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND 0.102f
C1464 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND 0.102f
C1465 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND 0.102f
C1466 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 11.386106f
C1467 a_21402_34716# VGND 0.39476f $ **FLOATING
C1468 a_17730_34716# VGND 0.39476f $ **FLOATING
C1469 a_16362_34716# VGND 0.39476f $ **FLOATING
C1470 a_12690_34716# VGND 0.39476f $ **FLOATING
C1471 a_11322_34716# VGND 0.39476f $ **FLOATING
C1472 a_7650_34716# VGND 0.39476f $ **FLOATING
C1473 a_6282_34716# VGND 0.39476f $ **FLOATING
C1474 a_2610_34716# VGND 0.394567f $ **FLOATING
C1475 a_22770_34892# VGND 0.394644f $ **FLOATING
C1476 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 2.276f
C1477 SUNSAR_SAR8B_CV_0.XA7.EN VGND 4.51439f
C1478 SUNSAR_SAR8B_CV_0.XA6.EN VGND 5.161865f
C1479 SUNSAR_SAR8B_CV_0.XA5.EN VGND 4.27708f
C1480 SUNSAR_SAR8B_CV_0.XA4.EN VGND 5.202775f
C1481 SUNSAR_SAR8B_CV_0.XA3.EN VGND 4.42572f
C1482 SUNSAR_SAR8B_CV_0.XA2.EN VGND 5.144325f
C1483 SUNSAR_SAR8B_CV_0.XA1.EN VGND 4.39222f
C1484 a_21402_35068# VGND 0.389563f $ **FLOATING
C1485 a_17730_35068# VGND 0.389563f $ **FLOATING
C1486 a_16362_35068# VGND 0.389563f $ **FLOATING
C1487 a_12690_35068# VGND 0.389563f $ **FLOATING
C1488 a_11322_35068# VGND 0.389563f $ **FLOATING
C1489 a_7650_35068# VGND 0.389563f $ **FLOATING
C1490 a_6282_35068# VGND 0.389563f $ **FLOATING
C1491 a_2610_35068# VGND 0.38937f $ **FLOATING
C1492 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C1493 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C1494 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C1495 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C1496 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C1497 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C1498 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557214f
C1499 a_22770_35420# VGND 0.395535f $ **FLOATING
C1500 a_21402_35420# VGND 0.389041f $ **FLOATING
C1501 a_17730_35420# VGND 0.388925f $ **FLOATING
C1502 a_16362_35420# VGND 0.389297f $ **FLOATING
C1503 a_12690_35420# VGND 0.388925f $ **FLOATING
C1504 a_11322_35420# VGND 0.389297f $ **FLOATING
C1505 a_7650_35420# VGND 0.388925f $ **FLOATING
C1506 a_6282_35420# VGND 0.389297f $ **FLOATING
C1507 a_2610_35420# VGND 0.389015f $ **FLOATING
C1508 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND 1.07685f
C1509 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND 0.112889f
C1510 SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND 1.50901f
C1511 SUNSAR_SAR8B_CV_0.XA7.XA9.B VGND 1.53168f
C1512 SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND 1.50964f
C1513 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND 0.112889f
C1514 SUNSAR_SAR8B_CV_0.XA6.XA9.B VGND 1.54335f
C1515 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND 0.112889f
C1516 SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND 1.51005f
C1517 SUNSAR_SAR8B_CV_0.XA5.XA9.B VGND 1.53305f
C1518 SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND 1.50964f
C1519 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND 0.112889f
C1520 SUNSAR_SAR8B_CV_0.XA4.XA9.B VGND 1.54335f
C1521 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND 0.112889f
C1522 SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND 1.51005f
C1523 SUNSAR_SAR8B_CV_0.XA3.XA9.B VGND 1.53305f
C1524 SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND 1.50964f
C1525 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND 0.112889f
C1526 SUNSAR_SAR8B_CV_0.XA2.XA9.B VGND 1.54335f
C1527 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND 0.112889f
C1528 SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND 1.51005f
C1529 SUNSAR_SAR8B_CV_0.XA1.XA9.B VGND 1.53305f
C1530 SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND 1.51935f
C1531 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND 0.112889f
C1532 SUNSAR_SAR8B_CV_0.XA0.XA9.B VGND 1.61753f
C1533 a_22770_35948# VGND 0.414038f $ **FLOATING
C1534 a_21402_35948# VGND 0.390722f $ **FLOATING
C1535 a_17730_35948# VGND 0.391291f $ **FLOATING
C1536 a_16362_35948# VGND 0.391291f $ **FLOATING
C1537 a_12690_35948# VGND 0.391291f $ **FLOATING
C1538 a_11322_35948# VGND 0.391291f $ **FLOATING
C1539 a_7650_35948# VGND 0.391291f $ **FLOATING
C1540 a_6282_35948# VGND 0.391291f $ **FLOATING
C1541 a_2610_35948# VGND 0.391099f $ **FLOATING
C1542 SUNSAR_SAR8B_CV_0.XA20.XA12.Y VGND 0.789814f
C1543 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C1544 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C1545 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C1546 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C1547 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C1548 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C1549 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C1550 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.895311f
C1551 a_22770_36300# VGND 0.472701f $ **FLOATING
C1552 a_21402_36300# VGND 0.393831f $ **FLOATING
C1553 a_17730_36300# VGND 0.394738f $ **FLOATING
C1554 a_16362_36300# VGND 0.3944f $ **FLOATING
C1555 a_12690_36300# VGND 0.394718f $ **FLOATING
C1556 a_11322_36300# VGND 0.3944f $ **FLOATING
C1557 a_7650_36300# VGND 0.394715f $ **FLOATING
C1558 a_6282_36300# VGND 0.3944f $ **FLOATING
C1559 a_2610_36300# VGND 0.394523f $ **FLOATING
C1560 a_22770_36652# VGND 0.542245f $ **FLOATING
C1561 SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND 0.881626f
C1562 SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND 0.884627f
C1563 SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND 0.877071f
C1564 SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND 0.884604f
C1565 SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND 0.877059f
C1566 SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND 0.884603f
C1567 SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND 0.877071f
C1568 SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND 0.892649f
C1569 SUNSAR_SAR8B_CV_0.XB2.TIE_L VGND 33.050705f
C1570 a_21402_36828# VGND 0.414041f $ **FLOATING
C1571 a_17730_36828# VGND 0.413952f $ **FLOATING
C1572 a_16362_36828# VGND 0.413659f $ **FLOATING
C1573 a_12690_36828# VGND 0.413942f $ **FLOATING
C1574 a_11322_36828# VGND 0.413658f $ **FLOATING
C1575 a_7650_36828# VGND 0.413944f $ **FLOATING
C1576 a_6282_36828# VGND 0.413659f $ **FLOATING
C1577 a_2610_36828# VGND 0.413594f $ **FLOATING
C1578 SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND 1.08552f
C1579 SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND 2.06017f
C1580 SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND 1.10839f
C1581 SUNSAR_SAR8B_CV_0.XA7.CEIN VGND 1.45333f
C1582 SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND 1.06778f
C1583 SUNSAR_SAR8B_CV_0.XA6.CEIN VGND 1.71757f
C1584 SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND 1.10834f
C1585 SUNSAR_SAR8B_CV_0.XA5.CEIN VGND 1.52588f
C1586 SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND 1.06777f
C1587 SUNSAR_SAR8B_CV_0.XA4.CEIN VGND 1.71756f
C1588 SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND 1.10835f
C1589 SUNSAR_SAR8B_CV_0.XA3.CEIN VGND 1.52589f
C1590 SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND 1.06778f
C1591 SUNSAR_SAR8B_CV_0.XA2.CEIN VGND 1.71756f
C1592 SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND 1.11927f
C1593 SUNSAR_SAR8B_CV_0.XA1.CEIN VGND 1.53308f
C1594 a_21402_37180# VGND 0.47501f $ **FLOATING
C1595 a_17730_37180# VGND 0.474809f $ **FLOATING
C1596 a_16362_37180# VGND 0.476355f $ **FLOATING
C1597 a_12690_37180# VGND 0.47479f $ **FLOATING
C1598 a_11322_37180# VGND 0.476354f $ **FLOATING
C1599 a_7650_37180# VGND 0.474794f $ **FLOATING
C1600 a_6282_37180# VGND 0.476355f $ **FLOATING
C1601 a_2610_37180# VGND 0.474277f $ **FLOATING
C1602 a_21402_37532# VGND 0.546649f $ **FLOATING
C1603 a_17730_37532# VGND 0.548986f $ **FLOATING
C1604 a_16362_37532# VGND 0.547631f $ **FLOATING
C1605 a_12690_37532# VGND 0.548815f $ **FLOATING
C1606 a_11322_37532# VGND 0.547631f $ **FLOATING
C1607 a_7650_37532# VGND 0.548857f $ **FLOATING
C1608 a_6282_37532# VGND 0.547634f $ **FLOATING
C1609 a_2610_37532# VGND 0.546853f $ **FLOATING
C1610 a_27575_39955# VGND 0.440387f $ **FLOATING
C1611 a_27575_40307# VGND 0.408627f $ **FLOATING
C1612 tt_um_TT06_SAR_done_0.x3.MP1.G VGND 1.07773f
C1613 a_27575_40659# VGND 0.389133f $ **FLOATING
C1614 tt_um_TT06_SAR_done_0.x4.MP0.G VGND 0.822801f
C1615 a_27575_41011# VGND 0.472703f $ **FLOATING
C1616 a_27575_41363# VGND 0.532318f $ **FLOATING
C1617 a_22790_40296# VGND 0.546732f $ **FLOATING
C1618 a_21422_40296# VGND 0.54563f $ **FLOATING
C1619 a_17750_40296# VGND 0.546813f $ **FLOATING
C1620 a_16382_40296# VGND 0.547966f $ **FLOATING
C1621 a_12710_40296# VGND 0.546813f $ **FLOATING
C1622 a_11342_40296# VGND 0.547969f $ **FLOATING
C1623 a_7670_40296# VGND 0.54681f $ **FLOATING
C1624 a_6302_40296# VGND 0.547966f $ **FLOATING
C1625 a_2630_40296# VGND 0.54539f $ **FLOATING
C1626 a_22790_40648# VGND 0.492438f $ **FLOATING
C1627 a_21422_40648# VGND 0.49034f $ **FLOATING
C1628 a_17750_40648# VGND 0.492453f $ **FLOATING
C1629 a_16382_40648# VGND 0.490883f $ **FLOATING
C1630 a_12710_40648# VGND 0.492453f $ **FLOATING
C1631 a_11342_40648# VGND 0.490883f $ **FLOATING
C1632 a_7670_40648# VGND 0.492453f $ **FLOATING
C1633 a_6302_40648# VGND 0.490883f $ **FLOATING
C1634 a_2630_40648# VGND 0.492826f $ **FLOATING
C1635 a_22790_41000# VGND 0.388777f $ **FLOATING
C1636 a_21422_41000# VGND 0.388174f $ **FLOATING
C1637 a_17750_41000# VGND 0.388174f $ **FLOATING
C1638 a_16382_41000# VGND 0.388174f $ **FLOATING
C1639 a_12710_41000# VGND 0.388174f $ **FLOATING
C1640 a_11342_41000# VGND 0.388174f $ **FLOATING
C1641 a_7670_41000# VGND 0.388174f $ **FLOATING
C1642 a_6302_41000# VGND 0.388174f $ **FLOATING
C1643 a_2630_41000# VGND 0.388638f $ **FLOATING
C1644 a_22790_41352# VGND 0.374594f $ **FLOATING
C1645 a_21422_41352# VGND 0.393558f $ **FLOATING
C1646 a_17750_41352# VGND 0.393558f $ **FLOATING
C1647 a_16382_41352# VGND 0.393558f $ **FLOATING
C1648 a_12710_41352# VGND 0.393558f $ **FLOATING
C1649 a_11342_41352# VGND 0.393558f $ **FLOATING
C1650 a_7670_41352# VGND 0.393558f $ **FLOATING
C1651 a_6302_41352# VGND 0.393558f $ **FLOATING
C1652 a_2630_41352# VGND 0.394022f $ **FLOATING
C1653 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND 0.803097f
C1654 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND 0.107737f
C1655 SUNSAR_SAR8B_CV_0.D<1> VGND 15.247869f
C1656 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND 0.107643f
C1657 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND 0.107643f
C1658 SUNSAR_SAR8B_CV_0.D<2> VGND 14.272022f
C1659 SUNSAR_SAR8B_CV_0.D<3> VGND 13.258019f
C1660 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND 0.107643f
C1661 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND 0.107643f
C1662 SUNSAR_SAR8B_CV_0.D<4> VGND 13.431784f
C1663 SUNSAR_SAR8B_CV_0.D<5> VGND 14.641789f
C1664 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND 0.107643f
C1665 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND 0.107643f
C1666 SUNSAR_SAR8B_CV_0.D<6> VGND 13.740876f
C1667 SUNSAR_SAR8B_CV_0.D<7> VGND 17.95158f
C1668 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND 0.107643f
C1669 a_22790_41880# VGND 0.394408f $ **FLOATING
C1670 a_21422_41880# VGND 0.395138f $ **FLOATING
C1671 a_17750_41880# VGND 0.395707f $ **FLOATING
C1672 a_16382_41880# VGND 0.395707f $ **FLOATING
C1673 a_12710_41880# VGND 0.395707f $ **FLOATING
C1674 a_11342_41880# VGND 0.395707f $ **FLOATING
C1675 a_7670_41880# VGND 0.395707f $ **FLOATING
C1676 a_6302_41880# VGND 0.395707f $ **FLOATING
C1677 a_2630_41880# VGND 0.396052f $ **FLOATING
C1678 SUNSAR_CAPT8B_CV_0.XA5.B VGND 1.96193f
C1679 a_22790_42408# VGND 0.410698f $ **FLOATING
C1680 a_21422_42408# VGND 0.389697f $ **FLOATING
C1681 a_17750_42408# VGND 0.390266f $ **FLOATING
C1682 a_16382_42408# VGND 0.390266f $ **FLOATING
C1683 a_12710_42408# VGND 0.390266f $ **FLOATING
C1684 a_11342_42408# VGND 0.390266f $ **FLOATING
C1685 a_7670_42408# VGND 0.390266f $ **FLOATING
C1686 a_6302_42408# VGND 0.390266f $ **FLOATING
C1687 a_2630_42408# VGND 0.390612f $ **FLOATING
C1688 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C1689 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND 1.28758f
C1690 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND 1.27933f
C1691 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND 1.27933f
C1692 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND 1.27933f
C1693 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND 1.27933f
C1694 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND 1.27933f
C1695 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND 1.27933f
C1696 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND 1.29578f
C1697 a_22790_42760# VGND 0.378208f $ **FLOATING
C1698 a_21422_42760# VGND 0.393027f $ **FLOATING
C1699 a_17750_42760# VGND 0.393596f $ **FLOATING
C1700 a_16382_42760# VGND 0.393596f $ **FLOATING
C1701 a_12710_42760# VGND 0.393596f $ **FLOATING
C1702 a_11342_42760# VGND 0.393596f $ **FLOATING
C1703 a_7670_42760# VGND 0.393596f $ **FLOATING
C1704 a_6302_42760# VGND 0.393596f $ **FLOATING
C1705 a_2630_42760# VGND 0.393942f $ **FLOATING
C1706 a_22790_43112# VGND 0.388427f $ **FLOATING
C1707 SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND 1.29446f
C1708 SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND 1.29655f
C1709 SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND 1.29655f
C1710 SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND 1.29655f
C1711 SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND 1.29655f
C1712 SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND 1.29655f
C1713 SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND 1.29655f
C1714 SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND 1.29893f
C1715 SUNSAR_CAPT8B_CV_0.XA6.A VGND 2.38038f
C1716 a_21422_43288# VGND 0.394124f $ **FLOATING
C1717 a_17750_43288# VGND 0.394693f $ **FLOATING
C1718 a_16382_43288# VGND 0.394693f $ **FLOATING
C1719 a_12710_43288# VGND 0.394693f $ **FLOATING
C1720 a_11342_43288# VGND 0.394693f $ **FLOATING
C1721 a_7670_43288# VGND 0.394693f $ **FLOATING
C1722 a_6302_43288# VGND 0.394693f $ **FLOATING
C1723 a_2630_43288# VGND 0.395039f $ **FLOATING
C1724 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND 0.103608f
C1725 SUNSAR_CAPT8B_CV_0.XA6.B VGND 1.65375f
C1726 a_22790_43640# VGND 0.387806f $ **FLOATING
C1727 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND 0.112889f
C1728 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN VGND 1.69058f
C1729 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND 0.112889f
C1730 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN VGND 1.69315f
C1731 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND 0.112889f
C1732 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN VGND 1.69315f
C1733 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND 0.112889f
C1734 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN VGND 1.69315f
C1735 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND 0.112889f
C1736 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN VGND 1.69797f
C1737 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND 0.112889f
C1738 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN VGND 1.69797f
C1739 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND 0.112889f
C1740 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN VGND 1.69797f
C1741 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND 0.112889f
C1742 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN VGND 1.69726f
C1743 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.88269f
C1744 a_21422_43816# VGND 0.390629f $ **FLOATING
C1745 a_17750_43816# VGND 0.391198f $ **FLOATING
C1746 a_16382_43816# VGND 0.391198f $ **FLOATING
C1747 a_12710_43816# VGND 0.391198f $ **FLOATING
C1748 a_11342_43816# VGND 0.391198f $ **FLOATING
C1749 a_7670_43816# VGND 0.391198f $ **FLOATING
C1750 a_6302_43816# VGND 0.391198f $ **FLOATING
C1751 a_2630_43816# VGND 0.391544f $ **FLOATING
C1752 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 32.775158f
C1753 a_22790_43992# VGND 0.384235f $ **FLOATING
C1754 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.23582f
C1755 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.23517f
C1756 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.23517f
C1757 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.23517f
C1758 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26123f
C1759 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C1760 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C1761 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C1762 SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND 0.5774f
C1763 a_21422_44168# VGND 0.425534f $ **FLOATING
C1764 a_17750_44168# VGND 0.425449f $ **FLOATING
C1765 a_16382_44168# VGND 0.425864f $ **FLOATING
C1766 a_12710_44168# VGND 0.425449f $ **FLOATING
C1767 a_11342_44168# VGND 0.425864f $ **FLOATING
C1768 a_7670_44168# VGND 0.425449f $ **FLOATING
C1769 a_6302_44168# VGND 0.425864f $ **FLOATING
C1770 a_2630_44168# VGND 0.426034f $ **FLOATING
C1771 TIE_L VGND 6.36945f
C1772 a_22790_44344# VGND 0.423601f $ **FLOATING
C1773 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n0 VGND 0.134084f
C1774 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n1 VGND 0.383793f
C1775 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n2 VGND 4.98541f
C1776 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n3 VGND 5.21883f
C1777 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n4 VGND 0.488995f
C1778 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n5 VGND 0.488995f
C1779 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n6 VGND 9.802549f
C1780 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n7 VGND 4.78669f
C1781 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n8 VGND 9.27166f
C1782 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n9 VGND 1.12383f
C1783 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n10 VGND 9.60336f
C1784 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n11 VGND 4.8841f
C1785 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n12 VGND 5.51583f
C1786 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n13 VGND 13.1294f
C1787 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n14 VGND 5.68794f
C1788 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n15 VGND 0.189948f
C1789 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB4.A VGND 0.325863f
C1790 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n16 VGND 0.383793f
C1791 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n17 VGND 4.98541f
C1792 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n18 VGND 5.21883f
C1793 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n19 VGND 0.488995f
C1794 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n20 VGND 0.488995f
C1795 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n21 VGND 9.802549f
C1796 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n22 VGND 4.78669f
C1797 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n23 VGND 9.27166f
C1798 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n24 VGND 1.12383f
C1799 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n25 VGND 9.60336f
C1800 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n26 VGND 4.8841f
C1801 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n27 VGND 5.51583f
C1802 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n28 VGND 13.1294f
C1803 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n29 VGND 5.68794f
C1804 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n30 VGND 0.189948f
C1805 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n31 VGND 0.611883f
C1806 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n32 VGND 0.383793f
C1807 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n33 VGND 4.98541f
C1808 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n34 VGND 5.21883f
C1809 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n35 VGND 0.488995f
C1810 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n36 VGND 0.488995f
C1811 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n37 VGND 9.802549f
C1812 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n38 VGND 4.78669f
C1813 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n39 VGND 9.27166f
C1814 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n40 VGND 1.12383f
C1815 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n41 VGND 9.60336f
C1816 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n42 VGND 4.8841f
C1817 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n43 VGND 5.51583f
C1818 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n44 VGND 13.1294f
C1819 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n45 VGND 5.68794f
C1820 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n46 VGND 0.189948f
C1821 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n47 VGND 0.581839f
C1822 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n48 VGND 0.383793f
C1823 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n49 VGND 4.98541f
C1824 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n50 VGND 5.21883f
C1825 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n51 VGND 0.488995f
C1826 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n52 VGND 0.488995f
C1827 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n53 VGND 9.802549f
C1828 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n54 VGND 4.78669f
C1829 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n55 VGND 9.27166f
C1830 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n56 VGND 1.12383f
C1831 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n57 VGND 9.60336f
C1832 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n58 VGND 4.8841f
C1833 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n59 VGND 5.51583f
C1834 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n60 VGND 13.1294f
C1835 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n61 VGND 5.68794f
C1836 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n62 VGND 0.189948f
C1837 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n63 VGND 0.319324f
C1838 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n64 VGND 0.383793f
C1839 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n65 VGND 4.98541f
C1840 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n66 VGND 5.21883f
C1841 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n67 VGND 0.488995f
C1842 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n68 VGND 0.488995f
C1843 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n69 VGND 9.802549f
C1844 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n70 VGND 4.78669f
C1845 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n71 VGND 9.27166f
C1846 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n72 VGND 1.12383f
C1847 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n73 VGND 9.60336f
C1848 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n74 VGND 4.8841f
C1849 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n75 VGND 5.51583f
C1850 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n76 VGND 13.1294f
C1851 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n77 VGND 5.68794f
C1852 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n78 VGND 0.189948f
C1853 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.XCAPB0.A VGND 0.30117f
C1854 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n79 VGND 1.01237f
C1855 SUNSAR_SAR8B_CV_0.XB2.XA4.GNG.n80 VGND 0.329585f
C1856 SUNSAR_SAR8B_CV_0.XA7.ENO.t3 VGND 0.118384f
C1857 SUNSAR_SAR8B_CV_0.XA7.ENO.t2 VGND 0.116907f
C1858 SUNSAR_SAR8B_CV_0.XA7.ENO.n1 VGND 0.252453f
C1859 SUNSAR_SAR8B_CV_0.XA7.ENO.n2 VGND 0.124505f
C1860 SUNSAR_SAR8B_CV_0.XA7.ENO.n3 VGND 0.248709f
C1861 SUNSAR_SAR8B_CV_0.XA7.ENO.t4 VGND 0.118384f
C1862 SUNSAR_SAR8B_CV_0.XA7.ENO.t5 VGND 0.114198f
C1863 SUNSAR_SAR8B_CV_0.XA7.ENO.n5 VGND 1.10167f
C1864 SUNSAR_SAR8B_CV_0.XA7.ENO.n7 VGND 1.62495f
C1865 uo_out[6].n1 VGND 0.112549f
C1866 uo_out[6].n3 VGND 0.217632f
C1867 uo_out[6].n6 VGND 0.720805f
C1868 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n0 VGND 0.102978f
C1869 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n3 VGND 0.102978f
C1870 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n4 VGND 0.102978f
C1871 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n5 VGND 0.102978f
C1872 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n8 VGND 0.31929f
C1873 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_OP.n9 VGND 0.344724f
C1874 SUNSAR_SAR8B_CV_0.XB2.CKN.n1 VGND 0.161451f
C1875 SUNSAR_SAR8B_CV_0.XB2.CKN.n3 VGND 0.117006f
C1876 SUNSAR_SAR8B_CV_0.XB2.CKN.n4 VGND 0.117006f
C1877 SUNSAR_SAR8B_CV_0.XB2.CKN.n7 VGND 0.186157f
C1878 SUNSAR_SAR8B_CV_0.XB2.XA4.MP0.G VGND 0.113391f
C1879 SUNSAR_SAR8B_CV_0.XB2.CKN.n11 VGND 0.241449f
C1880 SUNSAR_SAR8B_CV_0.XB2.CKN.n12 VGND 0.300724f
C1881 uo_out[7].n0 VGND 0.177819f
C1882 uo_out[7].n1 VGND 0.135771f
C1883 uo_out[7].n6 VGND 0.76451f
C1884 SUNSAR_SAR8B_CV_0.D<0>.n2 VGND 0.125441f
C1885 SUNSAR_SAR8B_CV_0.D<0>.n3 VGND 0.106281f
C1886 SUNSAR_SAR8B_CV_0.D<0>.n4 VGND 0.237622f
C1887 SUNSAR_SAR8B_CV_0.D<0>.n6 VGND 0.639161f
C1888 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP0.G VGND 0.121566f
C1889 SUNSAR_SAR8B_CV_0.D<0>.n11 VGND 0.230363f
C1890 SUNSAR_SAR8B_CV_0.D<0>.n12 VGND 1.16213f
C1891 SUNSAR_SAR8B_CV_0.D<0>.n13 VGND 1.45057f
C1892 SUNSAR_SAR8B_CV_0.D<0>.n20 VGND 0.114807f
C1893 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n1 VGND 0.256077f
C1894 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n2 VGND 0.203326f
C1895 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n4 VGND 0.20339f
C1896 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n5 VGND 0.402663f
C1897 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n8 VGND 0.123619f
C1898 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n10 VGND 0.391361f
C1899 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n11 VGND 0.236748f
C1900 SUNSAR_CAPT8B_CV_0.XG12.XA2.MN0.G VGND 0.108664f
C1901 SUNSAR_CAPT8B_CV_0.XG12.XA1.Y.n13 VGND 0.14197f
C1902 ua[0].n2 VGND 1.39243f
C1903 ua[0].n15 VGND 0.1295f
C1904 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n0 VGND 0.1444f
C1905 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n1 VGND 0.130728f
C1906 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n2 VGND 0.130728f
C1907 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n3 VGND 0.1444f
C1908 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n4 VGND 0.1444f
C1909 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n5 VGND 0.1444f
C1910 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n6 VGND 0.130728f
C1911 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n7 VGND 0.130728f
C1912 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_ON.n9 VGND 0.11907f
C1913 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.D VGND 0.100265f
C1914 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n0 VGND 0.425177f
C1915 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n1 VGND 4.75946f
C1916 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n2 VGND 0.105629f
C1917 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n4 VGND 0.146554f
C1918 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n5 VGND 0.203243f
C1919 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n6 VGND 0.105629f
C1920 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n7 VGND 0.145294f
C1921 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n8 VGND 0.209128f
C1922 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n11 VGND 0.216814f
C1923 SUNSAR_SAR8B_CV_0.XDAC2.CP<1>.n12 VGND 0.403927f
C1924 SUNSAR_SAR8B_CV_0.XA5.CP0.n0 VGND 0.110522f
C1925 SUNSAR_SAR8B_CV_0.XA5.CP0.n1 VGND 0.100058f
C1926 SUNSAR_SAR8B_CV_0.XA5.CP0.n2 VGND 0.100058f
C1927 SUNSAR_SAR8B_CV_0.XA5.CP0.n3 VGND 0.110522f
C1928 SUNSAR_SAR8B_CV_0.XA5.CP0.n4 VGND 0.110522f
C1929 SUNSAR_SAR8B_CV_0.XA5.CP0.n5 VGND 0.110522f
C1930 SUNSAR_SAR8B_CV_0.XA5.CP0.n6 VGND 0.100058f
C1931 SUNSAR_SAR8B_CV_0.XA5.CP0.n7 VGND 0.100058f
C1932 SUNSAR_SAR8B_CV_0.XA5.CP0.n9 VGND 0.117745f
C1933 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n1 VGND 0.256077f
C1934 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n2 VGND 0.203326f
C1935 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n4 VGND 0.20339f
C1936 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n5 VGND 0.402663f
C1937 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n8 VGND 0.123619f
C1938 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n10 VGND 0.391361f
C1939 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n11 VGND 0.236748f
C1940 SUNSAR_CAPT8B_CV_0.XI14.XA2.MN0.G VGND 0.108664f
C1941 SUNSAR_CAPT8B_CV_0.XI14.XA1.Y.n13 VGND 0.14197f
C1942 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n1 VGND 0.141664f
C1943 SUNSAR_SAR8B_CV_0.XA20.XA2.MN6.G VGND 0.137288f
C1944 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.t14 VGND 0.103258f
C1945 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n2 VGND 0.141664f
C1946 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n3 VGND 0.141003f
C1947 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n5 VGND 0.15648f
C1948 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n6 VGND 0.141664f
C1949 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n7 VGND 0.141664f
C1950 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n8 VGND 0.15648f
C1951 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n9 VGND 0.15648f
C1952 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n10 VGND 0.15648f
C1953 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n11 VGND 0.141664f
C1954 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n12 VGND 0.126187f
C1955 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n14 VGND 0.821361f
C1956 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n15 VGND 0.250881f
C1957 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n16 VGND 0.132395f
C1958 SUNSAR_SAR8B_CV_0.XA20.XA2.VMR.n18 VGND 0.180043f
C1959 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n0 VGND 0.131525f
C1960 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n2 VGND 0.148791f
C1961 SUNSAR_SAR8B_CV_0.XB1.XA3.MN1.D VGND 0.292689f
C1962 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n3 VGND 0.202878f
C1963 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n4 VGND 3.85261f
C1964 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n5 VGND 0.407483f
C1965 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n6 VGND 0.407483f
C1966 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n7 VGND 9.128111f
C1967 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n8 VGND 13.252201f
C1968 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n9 VGND 0.329004f
C1969 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n10 VGND 13.252201f
C1970 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n11 VGND 0.407483f
C1971 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n12 VGND 0.407483f
C1972 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n13 VGND 5.54943f
C1973 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n14 VGND 4.85685f
C1974 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n15 VGND 9.526259f
C1975 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n16 VGND 4.989491f
C1976 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n17 VGND 4.75996f
C1977 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n18 VGND 9.128111f
C1978 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n19 VGND 1.17804f
C1979 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n20 VGND 9.72281f
C1980 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n21 VGND 4.95706f
C1981 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n22 VGND 5.56704f
C1982 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n23 VGND 0.162841f
C1983 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB4.B VGND 0.322338f
C1984 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n24 VGND 0.329004f
C1985 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n25 VGND 4.95706f
C1986 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n26 VGND 4.989491f
C1987 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n27 VGND 9.526259f
C1988 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n28 VGND 1.17804f
C1989 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n29 VGND 9.72281f
C1990 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n30 VGND 0.407483f
C1991 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n31 VGND 9.128111f
C1992 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n32 VGND 4.75996f
C1993 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n33 VGND 0.407483f
C1994 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n34 VGND 4.85685f
C1995 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n35 VGND 5.54943f
C1996 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n36 VGND 13.252201f
C1997 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n37 VGND 5.56704f
C1998 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n38 VGND 0.162841f
C1999 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n39 VGND 0.605263f
C2000 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n40 VGND 0.329004f
C2001 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n41 VGND 4.95706f
C2002 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n42 VGND 4.989491f
C2003 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n43 VGND 9.526259f
C2004 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n44 VGND 1.17804f
C2005 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n45 VGND 9.72281f
C2006 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n46 VGND 0.407483f
C2007 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n47 VGND 9.128111f
C2008 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n48 VGND 4.75996f
C2009 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n49 VGND 0.407483f
C2010 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n50 VGND 4.85685f
C2011 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n51 VGND 5.54943f
C2012 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n52 VGND 13.252201f
C2013 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n53 VGND 5.56704f
C2014 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n54 VGND 0.162841f
C2015 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n55 VGND 0.575545f
C2016 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n56 VGND 0.329004f
C2017 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n57 VGND 4.95706f
C2018 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n58 VGND 4.989491f
C2019 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n59 VGND 9.526259f
C2020 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n60 VGND 1.17804f
C2021 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n61 VGND 9.72281f
C2022 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n62 VGND 0.407483f
C2023 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n63 VGND 9.128111f
C2024 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n64 VGND 4.75996f
C2025 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n65 VGND 0.407483f
C2026 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n66 VGND 4.85685f
C2027 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n67 VGND 5.54943f
C2028 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n68 VGND 13.252201f
C2029 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n69 VGND 5.56704f
C2030 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n70 VGND 0.162841f
C2031 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n71 VGND 0.605263f
C2032 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB0.B VGND 0.322338f
C2033 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n72 VGND 0.162841f
C2034 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n73 VGND 4.75996f
C2035 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n74 VGND 4.989491f
C2036 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n75 VGND 0.329004f
C2037 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n76 VGND 5.54943f
C2038 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n77 VGND 4.85685f
C2039 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n78 VGND 9.526259f
C2040 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n79 VGND 1.17804f
C2041 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n80 VGND 9.72282f
C2042 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n81 VGND 2.53222f
C2043 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n82 VGND 3.31179f
C2044 SUNSAR_SAR8B_CV_0.XB1.XA3.B.n83 VGND 2.38206f
C2045 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n0 VGND 0.102978f
C2046 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n3 VGND 0.102978f
C2047 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n4 VGND 0.102978f
C2048 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n5 VGND 0.102978f
C2049 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n8 VGND 0.31929f
C2050 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_OP.n9 VGND 0.344724f
C2051 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n1 VGND 0.256077f
C2052 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n2 VGND 0.203326f
C2053 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n4 VGND 0.20339f
C2054 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n5 VGND 0.402663f
C2055 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n8 VGND 0.123619f
C2056 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n10 VGND 0.391361f
C2057 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n11 VGND 0.236748f
C2058 SUNSAR_CAPT8B_CV_0.XC08.XA2.MN0.G VGND 0.108664f
C2059 SUNSAR_CAPT8B_CV_0.XC08.XA1.Y.n13 VGND 0.14197f
C2060 SUNSAR_SAR8B_CV_0.XA5.ENO.n1 VGND 0.164081f
C2061 SUNSAR_SAR8B_CV_0.XA5.ENO.n3 VGND 0.161647f
C2062 SUNSAR_SAR8B_CV_0.XA5.ENO.n5 VGND 0.716027f
C2063 SUNSAR_SAR8B_CV_0.XA5.ENO.n6 VGND 0.122071f
C2064 SUNSAR_SAR8B_CV_0.XA5.ENO.n8 VGND 0.460551f
C2065 SUNSAR_SAR8B_CV_0.XA5.ENO.n9 VGND 0.237982f
C2066 SUNSAR_SAR8B_CV_0.XA5.ENO.n13 VGND 0.265622f
C2067 SUNSAR_SAR8B_CV_0.XA5.ENO.n15 VGND 1.05613f
C2068 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.D VGND 0.103605f
C2069 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n2 VGND 0.102978f
C2070 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n5 VGND 0.102978f
C2071 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n6 VGND 0.102978f
C2072 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n7 VGND 0.102978f
C2073 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n10 VGND 0.185977f
C2074 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_OP.n11 VGND 0.431108f
C2075 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n0 VGND 0.138624f
C2076 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n1 VGND 0.125499f
C2077 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n2 VGND 0.125499f
C2078 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n3 VGND 0.138624f
C2079 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n4 VGND 0.138624f
C2080 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n5 VGND 0.138624f
C2081 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n6 VGND 0.125499f
C2082 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n7 VGND 0.125499f
C2083 SUNSAR_SAR8B_CV_0.XA6.XA1.CHL_ON.n9 VGND 0.114307f
C2084 SUNSAR_SAR8B_CV_0.XA1.ENO.n0 VGND 0.164081f
C2085 SUNSAR_SAR8B_CV_0.XA1.ENO.n5 VGND 0.122071f
C2086 SUNSAR_SAR8B_CV_0.XA1.ENO.n7 VGND 0.460551f
C2087 SUNSAR_SAR8B_CV_0.XA1.ENO.n8 VGND 0.237982f
C2088 SUNSAR_SAR8B_CV_0.XA1.ENO.n12 VGND 0.716027f
C2089 SUNSAR_SAR8B_CV_0.XA1.ENO.n13 VGND 1.05613f
C2090 SUNSAR_SAR8B_CV_0.XA1.ENO.n15 VGND 0.265622f
C2091 SUNSAR_SAR8B_CV_0.XA1.ENO.n17 VGND 0.161647f
C2092 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n2 VGND 0.360526f
C2093 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n4 VGND 0.630025f
C2094 SUNSAR_SAR8B_CV_0.XA20.XA1.CKN.n5 VGND 0.104409f
C2095 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n0 VGND 0.105044f
C2096 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n1 VGND 0.420065f
C2097 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n2 VGND 4.5f
C2098 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n3 VGND 0.232891f
C2099 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n4 VGND 0.232891f
C2100 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n5 VGND 0.100295f
C2101 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n6 VGND 0.274879f
C2102 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n7 VGND 0.200277f
C2103 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n8 VGND 0.100295f
C2104 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n10 VGND 0.180425f
C2105 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n11 VGND 0.100295f
C2106 SUNSAR_SAR8B_CV_0.XDAC2.CP<2>.n13 VGND 0.218314f
C2107 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.D VGND 0.152072f
C2108 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n0 VGND 0.111648f
C2109 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n1 VGND 0.1444f
C2110 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n2 VGND 0.130728f
C2111 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n3 VGND 0.130728f
C2112 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n4 VGND 0.1444f
C2113 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n5 VGND 0.1444f
C2114 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n6 VGND 0.1444f
C2115 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n7 VGND 0.130728f
C2116 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_ON.n8 VGND 0.176497f
C2117 SUNSAR_SAR8B_CV_0.XA4.CN1.n2 VGND 0.111486f
C2118 SUNSAR_SAR8B_CV_0.XA4.CN1.n3 VGND 0.10093f
C2119 SUNSAR_SAR8B_CV_0.XA4.CN1.n4 VGND 0.10093f
C2120 SUNSAR_SAR8B_CV_0.XA4.CN1.n5 VGND 0.111486f
C2121 SUNSAR_SAR8B_CV_0.XA4.CN1.n6 VGND 0.111486f
C2122 SUNSAR_SAR8B_CV_0.XA4.CN1.n7 VGND 0.111486f
C2123 SUNSAR_SAR8B_CV_0.XA4.CN1.n8 VGND 0.10093f
C2124 SUNSAR_SAR8B_CV_0.XA4.CN1.n12 VGND 0.109181f
C2125 SUNSAR_SAR8B_CV_0.D<2>.n2 VGND 0.156423f
C2126 SUNSAR_SAR8B_CV_0.D<2>.n3 VGND 0.132532f
C2127 SUNSAR_SAR8B_CV_0.D<2>.n4 VGND 0.296312f
C2128 SUNSAR_SAR8B_CV_0.D<2>.n6 VGND 0.797026f
C2129 SUNSAR_SAR8B_CV_0.D<2>.n9 VGND 0.110573f
C2130 SUNSAR_SAR8B_CV_0.D<2>.t10 VGND 0.114016f
C2131 SUNSAR_SAR8B_CV_0.D<2>.t11 VGND 0.110199f
C2132 SUNSAR_SAR8B_CV_0.D<2>.n11 VGND 0.284379f
C2133 SUNSAR_SAR8B_CV_0.D<2>.n12 VGND 0.598339f
C2134 SUNSAR_SAR8B_CV_0.D<2>.n14 VGND 0.607933f
C2135 SUNSAR_SAR8B_CV_0.D<2>.n15 VGND 2.07028f
C2136 SUNSAR_SAR8B_CV_0.D<2>.n16 VGND 3.06123f
C2137 SUNSAR_SAR8B_CV_0.D<2>.n17 VGND 3.22646f
C2138 SUNSAR_SAR8B_CV_0.D<2>.n24 VGND 0.143163f
C2139 SUNSAR_SAR8B_CV_0.D<2>.n26 VGND 0.105733f
C2140 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n0 VGND 0.347864f
C2141 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n1 VGND 4.68702f
C2142 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n2 VGND 0.102823f
C2143 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n4 VGND 0.142661f
C2144 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n5 VGND 0.197845f
C2145 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n6 VGND 0.102823f
C2146 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n7 VGND 0.141435f
C2147 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n8 VGND 0.203573f
C2148 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n11 VGND 0.211055f
C2149 SUNSAR_SAR8B_CV_0.XDAC2.CP<3>.n12 VGND 0.393199f
C2150 SUNSAR_SAR8B_CV_0.D<6>.n3 VGND 0.1537f
C2151 SUNSAR_SAR8B_CV_0.D<6>.n4 VGND 0.130224f
C2152 SUNSAR_SAR8B_CV_0.D<6>.n5 VGND 0.291154f
C2153 SUNSAR_SAR8B_CV_0.D<6>.n7 VGND 0.783151f
C2154 SUNSAR_SAR8B_CV_0.D<6>.n11 VGND 0.103892f
C2155 SUNSAR_SAR8B_CV_0.D<6>.n12 VGND 0.140671f
C2156 SUNSAR_SAR8B_CV_0.D<6>.t9 VGND 0.112031f
C2157 SUNSAR_SAR8B_CV_0.D<6>.t10 VGND 0.108281f
C2158 SUNSAR_SAR8B_CV_0.D<6>.n16 VGND 0.28226f
C2159 SUNSAR_SAR8B_CV_0.D<6>.n17 VGND 1.19748f
C2160 SUNSAR_SAR8B_CV_0.D<6>.n18 VGND 2.06862f
C2161 SUNSAR_SAR8B_CV_0.D<6>.n19 VGND 3.07478f
C2162 SUNSAR_SAR8B_CV_0.D<6>.n20 VGND 3.66491f
C2163 SUNSAR_SAR8B_CV_0.D<6>.n24 VGND 0.108648f
C2164 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n0 VGND 0.1444f
C2165 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n1 VGND 0.130728f
C2166 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n2 VGND 0.130728f
C2167 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n3 VGND 0.1444f
C2168 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n4 VGND 0.1444f
C2169 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n5 VGND 0.1444f
C2170 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n6 VGND 0.130728f
C2171 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n7 VGND 0.130728f
C2172 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_ON.n9 VGND 0.11907f
C2173 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.D VGND 0.100265f
C2174 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n1 VGND 0.131284f
C2175 SUNSAR_SAR8B_CV_0.XA20.XA3.MN6.G VGND 0.136136f
C2176 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.t15 VGND 0.102391f
C2177 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n2 VGND 0.140475f
C2178 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n3 VGND 0.155167f
C2179 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n4 VGND 0.140475f
C2180 SUNSAR_SAR8B_CV_0.XA20.XA3.MP4.G VGND 0.246081f
C2181 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n5 VGND 0.155167f
C2182 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n6 VGND 0.140475f
C2183 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n7 VGND 0.140475f
C2184 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n8 VGND 0.155167f
C2185 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n9 VGND 0.155167f
C2186 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n10 VGND 0.155167f
C2187 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n11 VGND 0.140475f
C2188 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n12 VGND 0.140475f
C2189 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n13 VGND 0.448445f
C2190 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n15 VGND 0.220454f
C2191 SUNSAR_SAR8B_CV_0.XA20.XA2.CO.n16 VGND 0.178532f
C2192 SUNSAR_SAR8B_CV_0.XA20.XA2.MP3.D VGND 0.114275f
C2193 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP1.G VGND 0.126429f
C2194 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN1.G VGND 0.417001f
C2195 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN0.G VGND 0.299703f
C2196 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n2 VGND 0.140462f
C2197 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP1.G VGND 0.126429f
C2198 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n4 VGND 0.402711f
C2199 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n6 VGND 0.318237f
C2200 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP1.G VGND 0.126429f
C2201 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN1.G VGND 0.417001f
C2202 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN0.G VGND 0.299703f
C2203 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n8 VGND 0.140462f
C2204 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP1.G VGND 0.126429f
C2205 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n10 VGND 0.402711f
C2206 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n12 VGND 0.318237f
C2207 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP1.G VGND 0.126429f
C2208 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN1.G VGND 0.417001f
C2209 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN0.G VGND 0.299703f
C2210 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n14 VGND 0.140462f
C2211 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP1.G VGND 0.126429f
C2212 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n16 VGND 0.402711f
C2213 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n18 VGND 0.318237f
C2214 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP1.G VGND 0.126429f
C2215 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN1.G VGND 0.417001f
C2216 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN0.G VGND 0.299703f
C2217 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n20 VGND 0.502191f
C2218 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n21 VGND 1.05459f
C2219 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n22 VGND 0.779358f
C2220 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n23 VGND 0.737524f
C2221 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n24 VGND 0.779358f
C2222 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n25 VGND 0.737524f
C2223 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n26 VGND 0.819123f
C2224 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n27 VGND 0.643965f
C2225 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP1.G VGND 0.126429f
C2226 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n28 VGND 0.402711f
C2227 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n29 VGND 0.31799f
C2228 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n34 VGND 0.700488f
C2229 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n35 VGND 0.307664f
C2230 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n38 VGND 0.122293f
C2231 SUNSAR_SAR8B_CV_0.XA0.CMP_ON.n41 VGND 0.122293f
C2232 SUNSAR_SAR8B_CV_0.XA20.XA3a.MP2.D VGND 0.112811f
C2233 SUNSAR_SAR8B_CV_0.XA3.CP0.n0 VGND 0.110522f
C2234 SUNSAR_SAR8B_CV_0.XA3.CP0.n1 VGND 0.100058f
C2235 SUNSAR_SAR8B_CV_0.XA3.CP0.n2 VGND 0.100058f
C2236 SUNSAR_SAR8B_CV_0.XA3.CP0.n3 VGND 0.110522f
C2237 SUNSAR_SAR8B_CV_0.XA3.CP0.n4 VGND 0.110522f
C2238 SUNSAR_SAR8B_CV_0.XA3.CP0.n5 VGND 0.110522f
C2239 SUNSAR_SAR8B_CV_0.XA3.CP0.n6 VGND 0.100058f
C2240 SUNSAR_SAR8B_CV_0.XA3.CP0.n7 VGND 0.100058f
C2241 SUNSAR_SAR8B_CV_0.XA3.CP0.n9 VGND 0.117745f
C2242 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n0 VGND 0.102978f
C2243 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n3 VGND 0.102978f
C2244 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n4 VGND 0.102978f
C2245 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n5 VGND 0.102978f
C2246 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n8 VGND 0.31929f
C2247 SUNSAR_SAR8B_CV_0.XA3.XA1.CHL_OP.n9 VGND 0.344724f
C2248 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n1 VGND 0.225363f
C2249 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n2 VGND 0.372287f
C2250 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n5 VGND 0.131858f
C2251 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n7 VGND 0.389189f
C2252 SUNSAR_CAPT8B_CV_0.XH13.XA2.MN0.G VGND 0.108664f
C2253 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n8 VGND 0.168986f
C2254 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n10 VGND 0.236748f
C2255 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n13 VGND 0.147362f
C2256 SUNSAR_CAPT8B_CV_0.XH13.XA1.Y.n15 VGND 0.259645f
C2257 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n0 VGND 0.383793f
C2258 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n1 VGND 4.98541f
C2259 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB4.A VGND 2.39335f
C2260 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n2 VGND 5.21883f
C2261 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n3 VGND 0.488995f
C2262 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n4 VGND 0.488995f
C2263 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n5 VGND 9.802549f
C2264 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n6 VGND 4.78669f
C2265 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n7 VGND 9.27166f
C2266 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n8 VGND 1.12383f
C2267 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n9 VGND 9.60336f
C2268 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n10 VGND 4.8841f
C2269 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n11 VGND 5.51583f
C2270 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n12 VGND 13.1294f
C2271 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n13 VGND 3.2946f
C2272 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n14 VGND 0.506002f
C2273 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n15 VGND 0.383793f
C2274 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n16 VGND 4.98541f
C2275 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB3.A VGND 2.39335f
C2276 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n17 VGND 5.21883f
C2277 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n18 VGND 0.488995f
C2278 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n19 VGND 0.488995f
C2279 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n20 VGND 9.802549f
C2280 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n21 VGND 4.78669f
C2281 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n22 VGND 9.27166f
C2282 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n23 VGND 1.12383f
C2283 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n24 VGND 9.60336f
C2284 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n25 VGND 4.8841f
C2285 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n26 VGND 5.51583f
C2286 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n27 VGND 13.1294f
C2287 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n28 VGND 3.2946f
C2288 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n29 VGND 0.220704f
C2289 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n30 VGND 0.631704f
C2290 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n31 VGND 0.383793f
C2291 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n32 VGND 4.98541f
C2292 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB2.A VGND 2.39335f
C2293 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n33 VGND 5.21883f
C2294 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n34 VGND 0.488995f
C2295 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n35 VGND 0.488995f
C2296 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n36 VGND 9.802549f
C2297 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n37 VGND 4.78669f
C2298 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n38 VGND 9.27166f
C2299 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n39 VGND 1.12383f
C2300 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n40 VGND 9.60336f
C2301 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n41 VGND 4.8841f
C2302 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n42 VGND 5.51583f
C2303 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n43 VGND 13.1294f
C2304 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n44 VGND 3.2946f
C2305 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n45 VGND 0.220704f
C2306 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n46 VGND 0.591851f
C2307 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n47 VGND 0.383793f
C2308 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n48 VGND 4.98541f
C2309 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB1.A VGND 2.39335f
C2310 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n49 VGND 5.21883f
C2311 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n50 VGND 0.488995f
C2312 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n51 VGND 0.488995f
C2313 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n52 VGND 9.802549f
C2314 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n53 VGND 4.78669f
C2315 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n54 VGND 9.27166f
C2316 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n55 VGND 1.12383f
C2317 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n56 VGND 9.60336f
C2318 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n57 VGND 4.8841f
C2319 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n58 VGND 5.51583f
C2320 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n59 VGND 13.1294f
C2321 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n60 VGND 3.2946f
C2322 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n61 VGND 0.220704f
C2323 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n62 VGND 0.329336f
C2324 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n63 VGND 0.383793f
C2325 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n64 VGND 4.98541f
C2326 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.XCAPB0.A VGND 2.39335f
C2327 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n65 VGND 5.21883f
C2328 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n66 VGND 0.488995f
C2329 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n67 VGND 0.488995f
C2330 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n68 VGND 9.802549f
C2331 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n69 VGND 4.78669f
C2332 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n70 VGND 9.27166f
C2333 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n71 VGND 1.12383f
C2334 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n72 VGND 9.60336f
C2335 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n73 VGND 4.8841f
C2336 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n74 VGND 5.51583f
C2337 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n75 VGND 13.1294f
C2338 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n76 VGND 3.2946f
C2339 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n77 VGND 0.481257f
C2340 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n78 VGND 1.05738f
C2341 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n79 VGND 0.133633f
C2342 SUNSAR_SAR8B_CV_0.XB1.XA4.GNG.n80 VGND 0.291714f
C2343 SUNSAR_SAR8B_CV_0.XA3.ENO.n0 VGND 0.164081f
C2344 SUNSAR_SAR8B_CV_0.XA3.ENO.n5 VGND 0.122071f
C2345 SUNSAR_SAR8B_CV_0.XA3.ENO.n7 VGND 0.460551f
C2346 SUNSAR_SAR8B_CV_0.XA3.ENO.n8 VGND 0.237982f
C2347 SUNSAR_SAR8B_CV_0.XA3.ENO.n12 VGND 0.716027f
C2348 SUNSAR_SAR8B_CV_0.XA3.ENO.n13 VGND 1.05613f
C2349 SUNSAR_SAR8B_CV_0.XA3.ENO.n15 VGND 0.265622f
C2350 SUNSAR_SAR8B_CV_0.XA3.ENO.n17 VGND 0.161647f
C2351 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n1 VGND 0.256077f
C2352 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n2 VGND 0.203326f
C2353 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n4 VGND 0.20339f
C2354 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n5 VGND 0.402663f
C2355 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n8 VGND 0.123619f
C2356 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n10 VGND 0.391361f
C2357 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n11 VGND 0.236748f
C2358 SUNSAR_CAPT8B_CV_0.XE10.XA2.MN0.G VGND 0.108664f
C2359 SUNSAR_CAPT8B_CV_0.XE10.XA1.Y.n13 VGND 0.14197f
C2360 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n1 VGND 0.225363f
C2361 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n2 VGND 0.372287f
C2362 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n5 VGND 0.131858f
C2363 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n7 VGND 0.389189f
C2364 SUNSAR_CAPT8B_CV_0.XB07.XA2.MN0.G VGND 0.108664f
C2365 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n8 VGND 0.168986f
C2366 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n10 VGND 0.236748f
C2367 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n13 VGND 0.147362f
C2368 SUNSAR_CAPT8B_CV_0.XB07.XA1.Y.n15 VGND 0.259645f
C2369 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n5 VGND 0.170541f
C2370 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n6 VGND 3.68898f
C2371 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n13 VGND 0.179516f
C2372 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n18 VGND 0.531431f
C2373 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n19 VGND 3.34373f
C2374 SUNSAR_SAR8B_CV_0.XB1.TIE_L.n20 VGND 2.28514f
C2375 ua[1].n1 VGND 1.35775f
C2376 ua[1].n15 VGND 0.152982f
C2377 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.D VGND 0.103605f
C2378 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n2 VGND 0.102978f
C2379 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n5 VGND 0.102978f
C2380 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n6 VGND 0.102978f
C2381 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n7 VGND 0.102978f
C2382 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n10 VGND 0.185977f
C2383 SUNSAR_SAR8B_CV_0.XA2.XA1.CHL_OP.n11 VGND 0.431108f
C2384 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n1 VGND 0.225363f
C2385 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n2 VGND 0.372287f
C2386 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n5 VGND 0.131858f
C2387 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n7 VGND 0.389189f
C2388 SUNSAR_CAPT8B_CV_0.XD09.XA2.MN0.G VGND 0.108664f
C2389 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n8 VGND 0.168986f
C2390 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n10 VGND 0.236748f
C2391 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n13 VGND 0.147362f
C2392 SUNSAR_CAPT8B_CV_0.XD09.XA1.Y.n15 VGND 0.259645f
C2393 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n1 VGND 0.225363f
C2394 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n2 VGND 0.372287f
C2395 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n5 VGND 0.131858f
C2396 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n7 VGND 0.389189f
C2397 SUNSAR_CAPT8B_CV_0.XF11.XA2.MN0.G VGND 0.108664f
C2398 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n8 VGND 0.168986f
C2399 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n10 VGND 0.236748f
C2400 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n13 VGND 0.147362f
C2401 SUNSAR_CAPT8B_CV_0.XF11.XA1.Y.n15 VGND 0.259645f
C2402 SUNSAR_SAR8B_CV_0.SARP.t0 VGND 0.24003f
C2403 SUNSAR_SAR8B_CV_0.SARP.n0 VGND 0.148714f
C2404 SUNSAR_SAR8B_CV_0.SARP.n1 VGND 0.108353f
C2405 SUNSAR_SAR8B_CV_0.SARP.t4 VGND 0.24003f
C2406 SUNSAR_SAR8B_CV_0.SARP.n3 VGND 0.32617f
C2407 SUNSAR_SAR8B_CV_0.SARP.t5 VGND 0.24003f
C2408 SUNSAR_SAR8B_CV_0.SARP.n4 VGND 0.19119f
C2409 SUNSAR_SAR8B_CV_0.SARP.n5 VGND 0.445407f
C2410 SUNSAR_SAR8B_CV_0.SARP.t7 VGND 0.24003f
C2411 SUNSAR_SAR8B_CV_0.SARP.n6 VGND 0.19119f
C2412 SUNSAR_SAR8B_CV_0.SARP.n7 VGND 0.429071f
C2413 SUNSAR_SAR8B_CV_0.SARP.n8 VGND 0.221314f
C2414 SUNSAR_SAR8B_CV_0.SARP.t6 VGND 0.24003f
C2415 SUNSAR_SAR8B_CV_0.SARP.n9 VGND 0.105299f
C2416 SUNSAR_SAR8B_CV_0.SARP.n11 VGND 0.719468f
C2417 SUNSAR_SAR8B_CV_0.SARP.n12 VGND 2.27763f
C2418 SUNSAR_SAR8B_CV_0.SARP.n13 VGND 2.8494f
C2419 SUNSAR_SAR8B_CV_0.SARP.n14 VGND 2.98449f
C2420 SUNSAR_SAR8B_CV_0.SARP.n15 VGND 2.99867f
C2421 SUNSAR_SAR8B_CV_0.SARP.n16 VGND 2.99867f
C2422 SUNSAR_SAR8B_CV_0.SARP.n17 VGND 2.99867f
C2423 SUNSAR_SAR8B_CV_0.SARP.n18 VGND 2.99867f
C2424 SUNSAR_SAR8B_CV_0.SARP.n19 VGND 2.99867f
C2425 SUNSAR_SAR8B_CV_0.SARP.n20 VGND 2.99867f
C2426 SUNSAR_SAR8B_CV_0.SARP.n21 VGND 2.99867f
C2427 SUNSAR_SAR8B_CV_0.SARP.n22 VGND 2.99867f
C2428 SUNSAR_SAR8B_CV_0.SARP.n23 VGND 2.99867f
C2429 SUNSAR_SAR8B_CV_0.SARP.n24 VGND 2.99867f
C2430 SUNSAR_SAR8B_CV_0.SARP.n25 VGND 2.99867f
C2431 SUNSAR_SAR8B_CV_0.SARP.n26 VGND 2.99867f
C2432 SUNSAR_SAR8B_CV_0.SARP.n27 VGND 2.99867f
C2433 SUNSAR_SAR8B_CV_0.SARP.n28 VGND 2.99867f
C2434 SUNSAR_SAR8B_CV_0.SARP.n29 VGND 2.99867f
C2435 SUNSAR_SAR8B_CV_0.SARP.n30 VGND 2.99867f
C2436 SUNSAR_SAR8B_CV_0.SARP.n31 VGND 2.99867f
C2437 SUNSAR_SAR8B_CV_0.SARP.n32 VGND 2.99867f
C2438 SUNSAR_SAR8B_CV_0.SARP.n33 VGND 2.99867f
C2439 SUNSAR_SAR8B_CV_0.SARP.n34 VGND 2.99867f
C2440 SUNSAR_SAR8B_CV_0.SARP.n35 VGND 2.99867f
C2441 SUNSAR_SAR8B_CV_0.SARP.n36 VGND 2.99867f
C2442 SUNSAR_SAR8B_CV_0.SARP.n37 VGND 2.99867f
C2443 SUNSAR_SAR8B_CV_0.SARP.n38 VGND 2.99867f
C2444 SUNSAR_SAR8B_CV_0.SARP.n39 VGND 2.99867f
C2445 SUNSAR_SAR8B_CV_0.SARP.n40 VGND 2.99867f
C2446 SUNSAR_SAR8B_CV_0.SARP.n41 VGND 2.99867f
C2447 SUNSAR_SAR8B_CV_0.SARP.n42 VGND 2.99867f
C2448 SUNSAR_SAR8B_CV_0.SARP.n43 VGND 2.99867f
C2449 SUNSAR_SAR8B_CV_0.SARP.n44 VGND 3.14902f
C2450 SUNSAR_SAR8B_CV_0.SARP.n45 VGND 2.99867f
C2451 SUNSAR_SAR8B_CV_0.SARP.n46 VGND 2.99867f
C2452 SUNSAR_SAR8B_CV_0.SARP.n47 VGND 2.99867f
C2453 SUNSAR_SAR8B_CV_0.SARP.n48 VGND 2.99867f
C2454 SUNSAR_SAR8B_CV_0.SARP.n49 VGND 2.99867f
C2455 SUNSAR_SAR8B_CV_0.SARP.n50 VGND 2.99867f
C2456 SUNSAR_SAR8B_CV_0.SARP.n51 VGND 2.99867f
C2457 SUNSAR_SAR8B_CV_0.SARP.n52 VGND 2.99867f
C2458 SUNSAR_SAR8B_CV_0.SARP.n53 VGND 2.99867f
C2459 SUNSAR_SAR8B_CV_0.SARP.n54 VGND 2.99867f
C2460 SUNSAR_SAR8B_CV_0.SARP.n55 VGND 2.99867f
C2461 SUNSAR_SAR8B_CV_0.SARP.n56 VGND 2.99867f
C2462 SUNSAR_SAR8B_CV_0.SARP.n57 VGND 2.99867f
C2463 SUNSAR_SAR8B_CV_0.SARP.n58 VGND 2.99867f
C2464 SUNSAR_SAR8B_CV_0.SARP.n59 VGND 2.99867f
C2465 SUNSAR_SAR8B_CV_0.SARP.n60 VGND 2.99867f
C2466 SUNSAR_SAR8B_CV_0.SARP.n61 VGND 2.99867f
C2467 SUNSAR_SAR8B_CV_0.SARP.n62 VGND 2.99867f
C2468 SUNSAR_SAR8B_CV_0.SARP.n63 VGND 2.99867f
C2469 SUNSAR_SAR8B_CV_0.SARP.n64 VGND 2.99867f
C2470 SUNSAR_SAR8B_CV_0.SARP.n65 VGND 2.99867f
C2471 SUNSAR_SAR8B_CV_0.SARP.n66 VGND 2.99867f
C2472 SUNSAR_SAR8B_CV_0.SARP.n67 VGND 2.99867f
C2473 SUNSAR_SAR8B_CV_0.SARP.n68 VGND 2.99867f
C2474 SUNSAR_SAR8B_CV_0.SARP.n69 VGND 2.99867f
C2475 SUNSAR_SAR8B_CV_0.SARP.n70 VGND 2.99867f
C2476 SUNSAR_SAR8B_CV_0.SARP.n71 VGND 2.99867f
C2477 SUNSAR_SAR8B_CV_0.SARP.n72 VGND 2.99867f
C2478 SUNSAR_SAR8B_CV_0.SARP.n73 VGND 2.99867f
C2479 SUNSAR_SAR8B_CV_0.SARP.n74 VGND 2.99867f
C2480 SUNSAR_SAR8B_CV_0.SARP.n75 VGND 2.98449f
C2481 SUNSAR_SAR8B_CV_0.SARP.t17 VGND 0.141596f
C2482 SUNSAR_SAR8B_CV_0.SARP.n77 VGND 0.430551f
C2483 SUNSAR_SAR8B_CV_0.SARP.t15 VGND 0.141596f
C2484 SUNSAR_SAR8B_CV_0.SARP.n78 VGND 0.475581f
C2485 SUNSAR_SAR8B_CV_0.SARP.t16 VGND 0.141596f
C2486 SUNSAR_SAR8B_CV_0.SARP.n79 VGND 0.475581f
C2487 SUNSAR_SAR8B_CV_0.SARP.t10 VGND 0.141596f
C2488 SUNSAR_SAR8B_CV_0.SARP.n80 VGND 0.475581f
C2489 SUNSAR_SAR8B_CV_0.SARP.t9 VGND 0.141596f
C2490 SUNSAR_SAR8B_CV_0.SARP.n81 VGND 0.36479f
C2491 SUNSAR_SAR8B_CV_0.SARP.n82 VGND 0.171873f
C2492 SUNSAR_SAR8B_CV_0.SARP.t12 VGND 0.141596f
C2493 SUNSAR_SAR8B_CV_0.SARP.n83 VGND 0.430551f
C2494 SUNSAR_SAR8B_CV_0.SARP.t8 VGND 0.141596f
C2495 SUNSAR_SAR8B_CV_0.SARP.n84 VGND 0.475581f
C2496 SUNSAR_SAR8B_CV_0.SARP.t11 VGND 0.141596f
C2497 SUNSAR_SAR8B_CV_0.SARP.n85 VGND 0.475581f
C2498 SUNSAR_SAR8B_CV_0.SARP.t14 VGND 0.141596f
C2499 SUNSAR_SAR8B_CV_0.SARP.n86 VGND 0.475581f
C2500 SUNSAR_SAR8B_CV_0.SARP.t13 VGND 0.141596f
C2501 SUNSAR_SAR8B_CV_0.SARP.n87 VGND 0.36479f
C2502 SUNSAR_SAR8B_CV_0.SARP.n88 VGND 0.90714f
C2503 SUNSAR_SAR8B_CV_0.SARP.n89 VGND 8.80934f
C2504 SUNSAR_SAR8B_CV_0.SARP.n90 VGND 3.32668f
C2505 SUNSAR_SAR8B_CV_0.SARP.n91 VGND 4.22073f
C2506 SUNSAR_SAR8B_CV_0.SARP.n92 VGND 1.60941f
C2507 SUNSAR_SAR8B_CV_0.SARP.n93 VGND 1.60941f
C2508 SUNSAR_SAR8B_CV_0.SARP.n94 VGND 1.60941f
C2509 SUNSAR_SAR8B_CV_0.SARP.n95 VGND 1.60941f
C2510 SUNSAR_SAR8B_CV_0.SARP.n96 VGND 1.60941f
C2511 SUNSAR_SAR8B_CV_0.SARP.n97 VGND 1.60941f
C2512 SUNSAR_SAR8B_CV_0.SARP.n98 VGND 1.60941f
C2513 SUNSAR_SAR8B_CV_0.SARP.n99 VGND 1.60941f
C2514 SUNSAR_SAR8B_CV_0.SARP.n100 VGND 1.60941f
C2515 SUNSAR_SAR8B_CV_0.SARP.n101 VGND 1.60941f
C2516 SUNSAR_SAR8B_CV_0.SARP.n102 VGND 1.60941f
C2517 SUNSAR_SAR8B_CV_0.SARP.n103 VGND 1.60941f
C2518 SUNSAR_SAR8B_CV_0.SARP.n104 VGND 1.60941f
C2519 SUNSAR_SAR8B_CV_0.SARP.n105 VGND 1.60941f
C2520 SUNSAR_SAR8B_CV_0.SARP.n106 VGND 1.60941f
C2521 SUNSAR_SAR8B_CV_0.SARP.n107 VGND 1.60941f
C2522 SUNSAR_SAR8B_CV_0.SARP.n108 VGND 1.60941f
C2523 SUNSAR_SAR8B_CV_0.SARP.n109 VGND 1.60941f
C2524 SUNSAR_SAR8B_CV_0.SARP.n110 VGND 1.60941f
C2525 SUNSAR_SAR8B_CV_0.SARP.n111 VGND 1.60941f
C2526 SUNSAR_SAR8B_CV_0.SARP.n112 VGND 1.60941f
C2527 SUNSAR_SAR8B_CV_0.SARP.n113 VGND 1.60941f
C2528 SUNSAR_SAR8B_CV_0.SARP.n114 VGND 1.60941f
C2529 SUNSAR_SAR8B_CV_0.SARP.n115 VGND 1.60941f
C2530 SUNSAR_SAR8B_CV_0.SARP.n116 VGND 1.60941f
C2531 SUNSAR_SAR8B_CV_0.SARP.n117 VGND 1.60941f
C2532 SUNSAR_SAR8B_CV_0.SARP.n118 VGND 1.60941f
C2533 SUNSAR_SAR8B_CV_0.SARP.n119 VGND 1.60941f
C2534 SUNSAR_SAR8B_CV_0.SARP.n120 VGND 1.59523f
C2535 SUNSAR_SAR8B_CV_0.XDAC1.XC0.CTOP VGND 0.191794f
C2536 SUNSAR_SAR8B_CV_0.SARP.n121 VGND 10.8953f
C2537 SUNSAR_SAR8B_CV_0.SARP.n122 VGND 2.8494f
C2538 SUNSAR_SAR8B_CV_0.SARP.n123 VGND 2.8494f
C2539 SUNSAR_SAR8B_CV_0.SARP.n124 VGND 2.98449f
C2540 SUNSAR_SAR8B_CV_0.SARP.n125 VGND 2.99867f
C2541 SUNSAR_SAR8B_CV_0.SARP.n126 VGND 2.99867f
C2542 SUNSAR_SAR8B_CV_0.SARP.n127 VGND 2.99867f
C2543 SUNSAR_SAR8B_CV_0.SARP.n128 VGND 2.99867f
C2544 SUNSAR_SAR8B_CV_0.SARP.n129 VGND 2.99867f
C2545 SUNSAR_SAR8B_CV_0.SARP.n130 VGND 2.99867f
C2546 SUNSAR_SAR8B_CV_0.SARP.n131 VGND 2.99867f
C2547 SUNSAR_SAR8B_CV_0.SARP.n132 VGND 2.99867f
C2548 SUNSAR_SAR8B_CV_0.SARP.n133 VGND 2.99867f
C2549 SUNSAR_SAR8B_CV_0.SARP.n134 VGND 2.99867f
C2550 SUNSAR_SAR8B_CV_0.SARP.n135 VGND 2.99867f
C2551 SUNSAR_SAR8B_CV_0.SARP.n136 VGND 2.99867f
C2552 SUNSAR_SAR8B_CV_0.SARP.n137 VGND 2.99867f
C2553 SUNSAR_SAR8B_CV_0.SARP.n138 VGND 2.99867f
C2554 SUNSAR_SAR8B_CV_0.SARP.n139 VGND 2.99867f
C2555 SUNSAR_SAR8B_CV_0.SARP.n140 VGND 2.99867f
C2556 SUNSAR_SAR8B_CV_0.SARP.n141 VGND 2.99867f
C2557 SUNSAR_SAR8B_CV_0.SARP.n142 VGND 2.99867f
C2558 SUNSAR_SAR8B_CV_0.SARP.n143 VGND 2.99867f
C2559 SUNSAR_SAR8B_CV_0.SARP.n144 VGND 2.99867f
C2560 SUNSAR_SAR8B_CV_0.SARP.n145 VGND 2.99867f
C2561 SUNSAR_SAR8B_CV_0.SARP.n146 VGND 2.99867f
C2562 SUNSAR_SAR8B_CV_0.SARP.n147 VGND 2.99867f
C2563 SUNSAR_SAR8B_CV_0.SARP.n148 VGND 2.99867f
C2564 SUNSAR_SAR8B_CV_0.SARP.n149 VGND 2.99867f
C2565 SUNSAR_SAR8B_CV_0.SARP.n150 VGND 2.99867f
C2566 SUNSAR_SAR8B_CV_0.SARP.n151 VGND 2.99867f
C2567 SUNSAR_SAR8B_CV_0.SARP.n152 VGND 2.99867f
C2568 SUNSAR_SAR8B_CV_0.SARP.n153 VGND 2.99867f
C2569 SUNSAR_SAR8B_CV_0.SARP.n154 VGND 2.99867f
C2570 SUNSAR_SAR8B_CV_0.SARP.n155 VGND 2.99867f
C2571 SUNSAR_SAR8B_CV_0.SARP.n156 VGND 3.32668f
C2572 SUNSAR_SAR8B_CV_0.SARP.n157 VGND 4.22073f
C2573 SUNSAR_SAR8B_CV_0.SARP.n158 VGND 1.60941f
C2574 SUNSAR_SAR8B_CV_0.SARP.n159 VGND 1.60941f
C2575 SUNSAR_SAR8B_CV_0.SARP.n160 VGND 1.60941f
C2576 SUNSAR_SAR8B_CV_0.SARP.n161 VGND 1.60941f
C2577 SUNSAR_SAR8B_CV_0.SARP.n162 VGND 1.60941f
C2578 SUNSAR_SAR8B_CV_0.SARP.n163 VGND 1.60941f
C2579 SUNSAR_SAR8B_CV_0.SARP.n164 VGND 1.60941f
C2580 SUNSAR_SAR8B_CV_0.SARP.n165 VGND 1.60941f
C2581 SUNSAR_SAR8B_CV_0.SARP.n166 VGND 1.60941f
C2582 SUNSAR_SAR8B_CV_0.SARP.n167 VGND 1.60941f
C2583 SUNSAR_SAR8B_CV_0.SARP.n168 VGND 1.60941f
C2584 SUNSAR_SAR8B_CV_0.SARP.n169 VGND 1.60941f
C2585 SUNSAR_SAR8B_CV_0.SARP.n170 VGND 1.60941f
C2586 SUNSAR_SAR8B_CV_0.SARP.n171 VGND 1.60941f
C2587 SUNSAR_SAR8B_CV_0.SARP.n172 VGND 1.60941f
C2588 SUNSAR_SAR8B_CV_0.SARP.n173 VGND 1.60941f
C2589 SUNSAR_SAR8B_CV_0.SARP.n174 VGND 1.60941f
C2590 SUNSAR_SAR8B_CV_0.SARP.n175 VGND 1.60941f
C2591 SUNSAR_SAR8B_CV_0.SARP.n176 VGND 1.60941f
C2592 SUNSAR_SAR8B_CV_0.SARP.n177 VGND 1.60941f
C2593 SUNSAR_SAR8B_CV_0.SARP.n178 VGND 1.60941f
C2594 SUNSAR_SAR8B_CV_0.SARP.n179 VGND 1.60941f
C2595 SUNSAR_SAR8B_CV_0.SARP.n180 VGND 1.60941f
C2596 SUNSAR_SAR8B_CV_0.SARP.n181 VGND 1.60941f
C2597 SUNSAR_SAR8B_CV_0.SARP.n182 VGND 1.60941f
C2598 SUNSAR_SAR8B_CV_0.SARP.n183 VGND 1.60941f
C2599 SUNSAR_SAR8B_CV_0.SARP.n184 VGND 1.60941f
C2600 SUNSAR_SAR8B_CV_0.SARP.n185 VGND 1.60941f
C2601 SUNSAR_SAR8B_CV_0.SARP.n186 VGND 1.59523f
C2602 SUNSAR_SAR8B_CV_0.SARP.n187 VGND 3.72121f
C2603 SUNSAR_SAR8B_CV_0.SARP.n188 VGND 2.347f
C2604 SUNSAR_SAR8B_CV_0.SARP.t2 VGND 0.26643f
C2605 SUNSAR_SAR8B_CV_0.XB1.M1.S VGND 0.394563f
C2606 SUNSAR_SAR8B_CV_0.SARP.t1 VGND 0.26643f
C2607 SUNSAR_SAR8B_CV_0.XB1.M2.S VGND 0.254849f
C2608 SUNSAR_SAR8B_CV_0.SARP.n192 VGND 0.350613f
C2609 SUNSAR_SAR8B_CV_0.SARP.t3 VGND 0.26643f
C2610 SUNSAR_SAR8B_CV_0.XB1.M3.S VGND 0.254849f
C2611 SUNSAR_SAR8B_CV_0.SARP.n193 VGND 0.350613f
C2612 SUNSAR_SAR8B_CV_0.XB1.M4.S VGND 0.195585f
C2613 SUNSAR_SAR8B_CV_0.XB1.XA3.MP2.G VGND 0.174578f
C2614 SUNSAR_SAR8B_CV_0.XB1.CKN.n1 VGND 0.117006f
C2615 SUNSAR_SAR8B_CV_0.XB1.CKN.n2 VGND 0.117006f
C2616 SUNSAR_SAR8B_CV_0.XB1.CKN.n3 VGND 0.113905f
C2617 SUNSAR_SAR8B_CV_0.XB1.CKN.n5 VGND 0.191959f
C2618 SUNSAR_SAR8B_CV_0.XB1.XA4.MP0.G VGND 0.113391f
C2619 SUNSAR_SAR8B_CV_0.XB1.CKN.n7 VGND 0.323035f
C2620 SUNSAR_SAR8B_CV_0.XB1.CKN.n8 VGND 0.287424f
C2621 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n2 VGND 3.03099f
C2622 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n3 VGND 0.273946f
C2623 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n4 VGND 1.78848f
C2624 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n5 VGND 4.19212f
C2625 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW.n6 VGND 0.123571f
C2626 SUNSAR_SAR8B_CV_0.XA7.CP0.n0 VGND 0.114773f
C2627 SUNSAR_SAR8B_CV_0.XA7.CP0.n1 VGND 0.103906f
C2628 SUNSAR_SAR8B_CV_0.XA7.CP0.n2 VGND 0.103906f
C2629 SUNSAR_SAR8B_CV_0.XA7.CP0.n3 VGND 0.114773f
C2630 SUNSAR_SAR8B_CV_0.XA7.CP0.n4 VGND 0.114773f
C2631 SUNSAR_SAR8B_CV_0.XA7.CP0.n5 VGND 0.114773f
C2632 SUNSAR_SAR8B_CV_0.XA7.CP0.n6 VGND 0.103906f
C2633 SUNSAR_SAR8B_CV_0.XA7.CP0.n7 VGND 0.103906f
C2634 SUNSAR_SAR8B_CV_0.XA7.CP0.n9 VGND 0.122274f
C2635 SUNSAR_SAR8B_CV_0.XA7.CP0.n16 VGND 0.100223f
C2636 tt_um_TT06_SAR_done_0.DONE VGND 0.412317f
C2637 SUNSAR_SAR8B_CV_0.DONE.n4 VGND 0.114408f
C2638 SUNSAR_SAR8B_CV_0.DONE.n5 VGND 0.42406f
C2639 SUNSAR_SAR8B_CV_0.DONE.n6 VGND 0.114408f
C2640 SUNSAR_SAR8B_CV_0.DONE.n7 VGND 0.453177f
C2641 SUNSAR_SAR8B_CV_0.DONE.n8 VGND 0.114408f
C2642 SUNSAR_SAR8B_CV_0.DONE.n9 VGND 0.453177f
C2643 SUNSAR_SAR8B_CV_0.DONE.n10 VGND 0.114408f
C2644 SUNSAR_SAR8B_CV_0.DONE.n11 VGND 0.453177f
C2645 SUNSAR_SAR8B_CV_0.DONE.n12 VGND 0.114408f
C2646 SUNSAR_SAR8B_CV_0.DONE.n13 VGND 0.453177f
C2647 SUNSAR_SAR8B_CV_0.DONE.n14 VGND 0.114408f
C2648 SUNSAR_SAR8B_CV_0.DONE.n15 VGND 0.453177f
C2649 SUNSAR_SAR8B_CV_0.DONE.n16 VGND 0.114408f
C2650 SUNSAR_SAR8B_CV_0.DONE.n17 VGND 0.453177f
C2651 SUNSAR_SAR8B_CV_0.DONE.n18 VGND 0.114408f
C2652 SUNSAR_SAR8B_CV_0.DONE.n19 VGND 0.419309f
C2653 SUNSAR_SAR8B_CV_0.DONE.n20 VGND 0.473087f
C2654 SUNSAR_SAR8B_CV_0.DONE.n21 VGND 0.78828f
C2655 SUNSAR_SAR8B_CV_0.XA5.CN1.n0 VGND 0.111486f
C2656 SUNSAR_SAR8B_CV_0.XA5.CN1.n1 VGND 0.10093f
C2657 SUNSAR_SAR8B_CV_0.XA5.CN1.n2 VGND 0.10093f
C2658 SUNSAR_SAR8B_CV_0.XA5.CN1.n3 VGND 0.111486f
C2659 SUNSAR_SAR8B_CV_0.XA5.CN1.n4 VGND 0.111486f
C2660 SUNSAR_SAR8B_CV_0.XA5.CN1.n5 VGND 0.111486f
C2661 SUNSAR_SAR8B_CV_0.XA5.CN1.n6 VGND 0.10093f
C2662 SUNSAR_SAR8B_CV_0.XA5.CN1.n10 VGND 0.118772f
C2663 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.D VGND 0.152072f
C2664 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n0 VGND 0.111648f
C2665 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n1 VGND 0.1444f
C2666 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n2 VGND 0.130728f
C2667 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n3 VGND 0.130728f
C2668 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n4 VGND 0.1444f
C2669 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n5 VGND 0.1444f
C2670 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n6 VGND 0.1444f
C2671 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n7 VGND 0.130728f
C2672 SUNSAR_SAR8B_CV_0.XA5.XA1.CHL_ON.n8 VGND 0.176497f
C2673 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n1 VGND 0.361801f
C2674 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n2 VGND 3.94329f
C2675 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n3 VGND 0.17066f
C2676 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n4 VGND 0.17066f
C2677 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n6 VGND 0.201429f
C2678 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n7 VGND 0.146762f
C2679 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n10 VGND 0.132214f
C2680 SUNSAR_SAR8B_CV_0.XDAC2.CP<0>.n13 VGND 0.159979f
C2681 SUNSAR_SAR8B_CV_0.XA6.CP0.n3 VGND 0.110522f
C2682 SUNSAR_SAR8B_CV_0.XA6.CP0.n4 VGND 0.100058f
C2683 SUNSAR_SAR8B_CV_0.XA6.CP0.n5 VGND 0.100058f
C2684 SUNSAR_SAR8B_CV_0.XA6.CP0.n6 VGND 0.110522f
C2685 SUNSAR_SAR8B_CV_0.XA6.CP0.n7 VGND 0.110522f
C2686 SUNSAR_SAR8B_CV_0.XA6.CP0.n8 VGND 0.110522f
C2687 SUNSAR_SAR8B_CV_0.XA6.CP0.n9 VGND 0.100058f
C2688 SUNSAR_SAR8B_CV_0.XA6.CP0.n10 VGND 0.186761f
C2689 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n0 VGND 0.102978f
C2690 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n3 VGND 0.102978f
C2691 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n4 VGND 0.102978f
C2692 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n5 VGND 0.102978f
C2693 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n8 VGND 0.31929f
C2694 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_OP.n9 VGND 0.344724f
C2695 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n0 VGND 0.11502f
C2696 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n1 VGND 0.381182f
C2697 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n2 VGND 5.29322f
C2698 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n3 VGND 0.25501f
C2699 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n4 VGND 0.25501f
C2700 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n5 VGND 0.109821f
C2701 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n6 VGND 0.300986f
C2702 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n7 VGND 0.219299f
C2703 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n8 VGND 0.109821f
C2704 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n10 VGND 0.197561f
C2705 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n11 VGND 0.109821f
C2706 SUNSAR_SAR8B_CV_0.XDAC2.CP<4>.n13 VGND 0.239049f
C2707 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n3 VGND 0.201952f
C2708 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n4 VGND 4.13388f
C2709 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n6 VGND 0.185267f
C2710 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n7 VGND 0.134148f
C2711 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n10 VGND 0.237968f
C2712 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n11 VGND 0.215436f
C2713 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t13 VGND 0.150375f
C2714 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t15 VGND 0.150375f
C2715 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n12 VGND 0.215436f
C2716 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n13 VGND 0.237968f
C2717 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t8 VGND 0.150375f
C2718 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t9 VGND 0.150375f
C2719 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n14 VGND 0.237968f
C2720 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t14 VGND 0.150375f
C2721 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t12 VGND 0.150375f
C2722 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n15 VGND 0.237968f
C2723 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n16 VGND 0.215436f
C2724 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t10 VGND 0.150375f
C2725 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.t11 VGND 0.150375f
C2726 SUNSAR_SAR8B_CV_0.XDAC1.CP<4>.n17 VGND 0.402118f
C2727 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n1 VGND 0.133651f
C2728 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n2 VGND 0.246608f
C2729 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n3 VGND 0.133651f
C2730 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n4 VGND 0.323828f
C2731 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n5 VGND 0.133651f
C2732 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n6 VGND 0.323828f
C2733 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n7 VGND 0.133651f
C2734 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n8 VGND 0.323828f
C2735 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n9 VGND 0.133651f
C2736 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n10 VGND 0.323828f
C2737 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n11 VGND 0.133651f
C2738 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n12 VGND 4.57855f
C2739 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n13 VGND 0.147328f
C2740 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n14 VGND 0.147328f
C2741 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n16 VGND 0.17389f
C2742 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n17 VGND 0.126697f
C2743 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n20 VGND 0.114138f
C2744 SUNSAR_SAR8B_CV_0.XDAC2.CP<8>.n23 VGND 0.138107f
C2745 SUNSAR_SAR8B_CV_0.D<1>.n4 VGND 0.130137f
C2746 SUNSAR_SAR8B_CV_0.D<1>.n5 VGND 0.115919f
C2747 SUNSAR_SAR8B_CV_0.D<1>.n6 VGND 0.463516f
C2748 SUNSAR_SAR8B_CV_0.D<1>.n7 VGND 0.487274f
C2749 SUNSAR_SAR8B_CV_0.D<1>.n8 VGND 0.100562f
C2750 SUNSAR_SAR8B_CV_0.D<1>.n10 VGND 0.23659f
C2751 SUNSAR_SAR8B_CV_0.D<1>.n12 VGND 0.461328f
C2752 SUNSAR_SAR8B_CV_0.D<1>.n13 VGND 0.555262f
C2753 SUNSAR_SAR8B_CV_0.D<1>.n14 VGND 1.75501f
C2754 SUNSAR_SAR8B_CV_0.D<1>.n15 VGND 2.59997f
C2755 SUNSAR_SAR8B_CV_0.D<1>.n16 VGND 2.73083f
C2756 SUNSAR_SAR8B_CV_0.D<1>.n24 VGND 0.119106f
C2757 SUNSAR_SAR8B_CV_0.XA6.CN1.n2 VGND 0.111486f
C2758 SUNSAR_SAR8B_CV_0.XA6.CN1.n3 VGND 0.10093f
C2759 SUNSAR_SAR8B_CV_0.XA6.CN1.n4 VGND 0.10093f
C2760 SUNSAR_SAR8B_CV_0.XA6.CN1.n5 VGND 0.111486f
C2761 SUNSAR_SAR8B_CV_0.XA6.CN1.n6 VGND 0.111486f
C2762 SUNSAR_SAR8B_CV_0.XA6.CN1.n7 VGND 0.111486f
C2763 SUNSAR_SAR8B_CV_0.XA6.CN1.n8 VGND 0.10093f
C2764 SUNSAR_SAR8B_CV_0.XA6.CN1.n12 VGND 0.109181f
C2765 SUNSAR_SAR8B_CV_0.XA7.CN1.n0 VGND 0.111486f
C2766 SUNSAR_SAR8B_CV_0.XA7.CN1.n1 VGND 0.10093f
C2767 SUNSAR_SAR8B_CV_0.XA7.CN1.n2 VGND 0.10093f
C2768 SUNSAR_SAR8B_CV_0.XA7.CN1.n3 VGND 0.111486f
C2769 SUNSAR_SAR8B_CV_0.XA7.CN1.n4 VGND 0.111486f
C2770 SUNSAR_SAR8B_CV_0.XA7.CN1.n5 VGND 0.111486f
C2771 SUNSAR_SAR8B_CV_0.XA7.CN1.n6 VGND 0.10093f
C2772 SUNSAR_SAR8B_CV_0.XA7.CN1.n10 VGND 0.118772f
C2773 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.D VGND 0.152072f
C2774 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n0 VGND 0.111648f
C2775 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n1 VGND 0.1444f
C2776 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n2 VGND 0.130728f
C2777 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n3 VGND 0.130728f
C2778 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n4 VGND 0.1444f
C2779 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n5 VGND 0.1444f
C2780 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n6 VGND 0.1444f
C2781 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n7 VGND 0.130728f
C2782 SUNSAR_SAR8B_CV_0.XA7.XA1.CHL_ON.n8 VGND 0.176497f
C2783 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n0 VGND 0.1444f
C2784 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n1 VGND 0.130728f
C2785 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n2 VGND 0.130728f
C2786 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n3 VGND 0.1444f
C2787 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n4 VGND 0.1444f
C2788 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n5 VGND 0.1444f
C2789 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n6 VGND 0.130728f
C2790 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n7 VGND 0.130728f
C2791 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_ON.n9 VGND 0.11907f
C2792 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.D VGND 0.100265f
C2793 SUNSAR_SAR8B_CV_0.EN.t0 VGND 0.111998f
C2794 SUNSAR_SAR8B_CV_0.EN.t1 VGND 0.127751f
C2795 SUNSAR_CAPT8B_CV_0.XA5a.MP0.D VGND 0.223258f
C2796 SUNSAR_SAR8B_CV_0.EN.n1 VGND 0.133422f
C2797 SUNSAR_SAR8B_CV_0.EN.n3 VGND 0.157584f
C2798 SUNSAR_SAR8B_CV_0.EN.n5 VGND 0.452906f
C2799 SUNSAR_SAR8B_CV_0.EN.n6 VGND 0.176982f
C2800 SUNSAR_SAR8B_CV_0.EN.n7 VGND 0.706547f
C2801 SUNSAR_SAR8B_CV_0.EN.n8 VGND 0.18242f
C2802 SUNSAR_SAR8B_CV_0.EN.n10 VGND 0.15763f
C2803 SUNSAR_SAR8B_CV_0.EN.n11 VGND 0.249566f
C2804 SUNSAR_SAR8B_CV_0.EN.n12 VGND 0.479383f
C2805 SUNSAR_SAR8B_CV_0.EN.n13 VGND 0.586856f
C2806 SUNSAR_SAR8B_CV_0.EN.n14 VGND 0.200896f
C2807 SUNSAR_SAR8B_CV_0.EN.n15 VGND 0.221907f
C2808 SUNSAR_SAR8B_CV_0.EN.n16 VGND 0.198172f
C2809 SUNSAR_SAR8B_CV_0.EN.n17 VGND 0.649437f
C2810 SUNSAR_SAR8B_CV_0.EN.n18 VGND 0.173522f
C2811 SUNSAR_SAR8B_CV_0.EN.n19 VGND 0.200896f
C2812 SUNSAR_SAR8B_CV_0.EN.n20 VGND 0.221907f
C2813 SUNSAR_SAR8B_CV_0.EN.n21 VGND 0.158095f
C2814 SUNSAR_SAR8B_CV_0.EN.n25 VGND 0.168089f
C2815 SUNSAR_SAR8B_CV_0.EN.n26 VGND 0.168089f
C2816 SUNSAR_SAR8B_CV_0.EN.n27 VGND 0.200896f
C2817 SUNSAR_SAR8B_CV_0.EN.n28 VGND 0.221907f
C2818 SUNSAR_SAR8B_CV_0.EN.n29 VGND 0.178353f
C2819 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP0.G VGND 0.62328f
C2820 SUNSAR_SAR8B_CV_0.EN.n30 VGND 0.200896f
C2821 SUNSAR_SAR8B_CV_0.EN.n31 VGND 0.221907f
C2822 SUNSAR_SAR8B_CV_0.EN.n32 VGND 0.200896f
C2823 SUNSAR_SAR8B_CV_0.EN.n33 VGND 0.591764f
C2824 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.G VGND 0.161327f
C2825 SUNSAR_SAR8B_CV_0.EN.n37 VGND 0.81243f
C2826 SUNSAR_SAR8B_CV_0.EN.n38 VGND 0.81243f
C2827 SUNSAR_SAR8B_CV_0.EN.n39 VGND 0.586856f
C2828 SUNSAR_SAR8B_CV_0.EN.n40 VGND 0.200896f
C2829 SUNSAR_SAR8B_CV_0.EN.n41 VGND 0.221907f
C2830 SUNSAR_SAR8B_CV_0.EN.n42 VGND 0.198172f
C2831 SUNSAR_SAR8B_CV_0.EN.n43 VGND 0.649437f
C2832 SUNSAR_SAR8B_CV_0.EN.n44 VGND 0.173522f
C2833 SUNSAR_SAR8B_CV_0.EN.n45 VGND 0.200896f
C2834 SUNSAR_SAR8B_CV_0.EN.n46 VGND 0.221907f
C2835 SUNSAR_SAR8B_CV_0.EN.n47 VGND 0.158095f
C2836 SUNSAR_SAR8B_CV_0.EN.n51 VGND 0.168089f
C2837 SUNSAR_SAR8B_CV_0.EN.n52 VGND 0.168089f
C2838 SUNSAR_SAR8B_CV_0.EN.n53 VGND 0.200896f
C2839 SUNSAR_SAR8B_CV_0.EN.n54 VGND 0.221907f
C2840 SUNSAR_SAR8B_CV_0.EN.n55 VGND 0.178353f
C2841 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP0.G VGND 0.62328f
C2842 SUNSAR_SAR8B_CV_0.EN.n56 VGND 0.200896f
C2843 SUNSAR_SAR8B_CV_0.EN.n57 VGND 0.221907f
C2844 SUNSAR_SAR8B_CV_0.EN.n58 VGND 0.200896f
C2845 SUNSAR_SAR8B_CV_0.EN.n59 VGND 0.591764f
C2846 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.G VGND 0.161327f
C2847 SUNSAR_SAR8B_CV_0.EN.n63 VGND 0.81243f
C2848 SUNSAR_SAR8B_CV_0.EN.n64 VGND 0.81243f
C2849 SUNSAR_SAR8B_CV_0.EN.n65 VGND 0.586856f
C2850 SUNSAR_SAR8B_CV_0.EN.n66 VGND 0.200896f
C2851 SUNSAR_SAR8B_CV_0.EN.n67 VGND 0.221907f
C2852 SUNSAR_SAR8B_CV_0.EN.n68 VGND 0.198172f
C2853 SUNSAR_SAR8B_CV_0.EN.n69 VGND 0.649437f
C2854 SUNSAR_SAR8B_CV_0.EN.n70 VGND 0.173522f
C2855 SUNSAR_SAR8B_CV_0.EN.n71 VGND 0.200896f
C2856 SUNSAR_SAR8B_CV_0.EN.n72 VGND 0.221907f
C2857 SUNSAR_SAR8B_CV_0.EN.n73 VGND 0.158095f
C2858 SUNSAR_SAR8B_CV_0.EN.n77 VGND 0.168089f
C2859 SUNSAR_SAR8B_CV_0.EN.n78 VGND 0.168089f
C2860 SUNSAR_SAR8B_CV_0.EN.n79 VGND 0.200896f
C2861 SUNSAR_SAR8B_CV_0.EN.n80 VGND 0.221907f
C2862 SUNSAR_SAR8B_CV_0.EN.n81 VGND 0.178353f
C2863 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP0.G VGND 0.62328f
C2864 SUNSAR_SAR8B_CV_0.EN.n82 VGND 0.200896f
C2865 SUNSAR_SAR8B_CV_0.EN.n83 VGND 0.221907f
C2866 SUNSAR_SAR8B_CV_0.EN.n84 VGND 0.200896f
C2867 SUNSAR_SAR8B_CV_0.EN.n85 VGND 0.591764f
C2868 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.G VGND 0.161327f
C2869 SUNSAR_SAR8B_CV_0.EN.n89 VGND 0.81243f
C2870 SUNSAR_SAR8B_CV_0.EN.n90 VGND 0.81243f
C2871 SUNSAR_SAR8B_CV_0.EN.n91 VGND 0.586856f
C2872 SUNSAR_SAR8B_CV_0.EN.n92 VGND 0.200896f
C2873 SUNSAR_SAR8B_CV_0.EN.n93 VGND 0.221907f
C2874 SUNSAR_SAR8B_CV_0.EN.n94 VGND 0.198172f
C2875 SUNSAR_SAR8B_CV_0.EN.n95 VGND 0.649437f
C2876 SUNSAR_SAR8B_CV_0.EN.n96 VGND 0.173522f
C2877 SUNSAR_SAR8B_CV_0.EN.n97 VGND 0.200896f
C2878 SUNSAR_SAR8B_CV_0.EN.n98 VGND 0.221907f
C2879 SUNSAR_SAR8B_CV_0.EN.n99 VGND 0.158095f
C2880 SUNSAR_SAR8B_CV_0.EN.n103 VGND 0.168089f
C2881 SUNSAR_SAR8B_CV_0.EN.n104 VGND 0.168089f
C2882 SUNSAR_SAR8B_CV_0.EN.n105 VGND 0.200896f
C2883 SUNSAR_SAR8B_CV_0.EN.n106 VGND 0.221907f
C2884 SUNSAR_SAR8B_CV_0.EN.n107 VGND 0.178353f
C2885 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP0.G VGND 0.62328f
C2886 SUNSAR_SAR8B_CV_0.EN.n108 VGND 0.200896f
C2887 SUNSAR_SAR8B_CV_0.EN.n109 VGND 0.221907f
C2888 SUNSAR_SAR8B_CV_0.EN.n110 VGND 0.200896f
C2889 SUNSAR_SAR8B_CV_0.EN.n111 VGND 0.591764f
C2890 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.G VGND 0.161327f
C2891 SUNSAR_SAR8B_CV_0.EN.n115 VGND 4.37092f
C2892 SUNSAR_CAPT8B_CV_0.EN VGND 4.01063f
C2893 SUNSAR_SAR8B_CV_0.EN.n116 VGND 0.247383f
C2894 SUNSAR_SAR8B_CV_0.D<5>.n4 VGND 0.142448f
C2895 SUNSAR_SAR8B_CV_0.D<5>.n5 VGND 0.126885f
C2896 SUNSAR_SAR8B_CV_0.D<5>.n6 VGND 0.507365f
C2897 SUNSAR_SAR8B_CV_0.D<5>.n7 VGND 0.533371f
C2898 SUNSAR_SAR8B_CV_0.D<5>.n8 VGND 0.110075f
C2899 SUNSAR_SAR8B_CV_0.D<5>.t9 VGND 0.103829f
C2900 SUNSAR_SAR8B_CV_0.D<5>.t11 VGND 0.100354f
C2901 SUNSAR_SAR8B_CV_0.D<5>.n10 VGND 0.253308f
C2902 SUNSAR_SAR8B_CV_0.D<5>.n12 VGND 0.503439f
C2903 SUNSAR_SAR8B_CV_0.D<5>.n14 VGND 0.578149f
C2904 SUNSAR_SAR8B_CV_0.D<5>.n15 VGND 1.93127f
C2905 SUNSAR_SAR8B_CV_0.D<5>.n16 VGND 0.535745f
C2906 SUNSAR_SAR8B_CV_0.D<5>.n17 VGND 0.693727f
C2907 SUNSAR_SAR8B_CV_0.D<5>.n18 VGND 0.610407f
C2908 SUNSAR_SAR8B_CV_0.D<5>.n19 VGND 1.9592f
C2909 SUNSAR_SAR8B_CV_0.D<5>.n20 VGND 2.37359f
C2910 SUNSAR_SAR8B_CV_0.D<5>.n28 VGND 0.130373f
C2911 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n2 VGND 0.135375f
C2912 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n3 VGND 0.122557f
C2913 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n4 VGND 0.122557f
C2914 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n5 VGND 0.135375f
C2915 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n6 VGND 0.135375f
C2916 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n7 VGND 0.135375f
C2917 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n8 VGND 0.122557f
C2918 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n11 VGND 0.164672f
C2919 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n12 VGND 0.357211f
C2920 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n13 VGND 0.164672f
C2921 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n14 VGND 0.493133f
C2922 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n15 VGND 0.164672f
C2923 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n16 VGND 0.421448f
C2924 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n17 VGND 0.164672f
C2925 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n18 VGND 2.30721f
C2926 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n19 VGND 3.0983f
C2927 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n21 VGND 0.132576f
C2928 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n24 VGND 0.114886f
C2929 SUNSAR_SAR8B_CV_0.XDAC2.CP<5>.n27 VGND 0.114886f
C2930 SUNSAR_SAR8B_CV_0.D<7>.n13 VGND 0.193847f
C2931 SUNSAR_SAR8B_CV_0.D<7>.n15 VGND 0.276504f
C2932 SUNSAR_SAR8B_CV_0.D<7>.n19 VGND 0.105783f
C2933 SUNSAR_SAR8B_CV_0.D<7>.n21 VGND 0.105783f
C2934 SUNSAR_SAR8B_CV_0.D<7>.n23 VGND 0.105783f
C2935 SUNSAR_SAR8B_CV_0.D<7>.n25 VGND 0.105783f
C2936 SUNSAR_SAR8B_CV_0.D<7>.n27 VGND 0.847145f
C2937 SUNSAR_SAR8B_CV_0.D<7>.n28 VGND 1.11546f
C2938 SUNSAR_SAR8B_CV_0.D<7>.n29 VGND 0.813962f
C2939 SUNSAR_SAR8B_CV_0.D<7>.n30 VGND 0.633723f
C2940 SUNSAR_SAR8B_CV_0.D<4>.n3 VGND 0.145913f
C2941 SUNSAR_SAR8B_CV_0.D<4>.n4 VGND 0.123627f
C2942 SUNSAR_SAR8B_CV_0.D<4>.n5 VGND 0.276403f
C2943 SUNSAR_SAR8B_CV_0.D<4>.n7 VGND 0.743476f
C2944 SUNSAR_SAR8B_CV_0.D<4>.n12 VGND 0.133545f
C2945 SUNSAR_SAR8B_CV_0.D<4>.t10 VGND 0.106355f
C2946 SUNSAR_SAR8B_CV_0.D<4>.t11 VGND 0.102795f
C2947 SUNSAR_SAR8B_CV_0.D<4>.n16 VGND 0.265272f
C2948 SUNSAR_SAR8B_CV_0.D<4>.n18 VGND 0.517599f
C2949 SUNSAR_SAR8B_CV_0.D<4>.n19 VGND 0.621382f
C2950 SUNSAR_SAR8B_CV_0.D<4>.n20 VGND 1.96001f
C2951 SUNSAR_SAR8B_CV_0.D<4>.n21 VGND 2.40683f
C2952 SUNSAR_SAR8B_CV_0.D<4>.n22 VGND 2.65925f
C2953 SUNSAR_SAR8B_CV_0.D<4>.n26 VGND 0.103144f
C2954 SUNSAR_SAR8B_CV_0.XA3.CN1.n4 VGND 0.111486f
C2955 SUNSAR_SAR8B_CV_0.XA3.CN1.n5 VGND 0.10093f
C2956 SUNSAR_SAR8B_CV_0.XA3.CN1.n6 VGND 0.10093f
C2957 SUNSAR_SAR8B_CV_0.XA3.CN1.n7 VGND 0.111486f
C2958 SUNSAR_SAR8B_CV_0.XA3.CN1.n8 VGND 0.111486f
C2959 SUNSAR_SAR8B_CV_0.XA3.CN1.n9 VGND 0.111486f
C2960 SUNSAR_SAR8B_CV_0.XA3.CN1.n10 VGND 0.10093f
C2961 SUNSAR_SAR8B_CV_0.XA3.CN1.n14 VGND 0.118772f
C2962 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n3 VGND 0.140662f
C2963 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n4 VGND 0.344208f
C2964 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n5 VGND 0.422857f
C2965 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n6 VGND 0.422857f
C2966 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n7 VGND 0.422857f
C2967 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n8 VGND 0.422857f
C2968 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n9 VGND 4.16724f
C2969 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n11 VGND 0.129041f
C2970 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n15 VGND 0.165748f
C2971 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n16 VGND 0.150054f
C2972 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t13 VGND 0.104738f
C2973 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t10 VGND 0.104738f
C2974 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n17 VGND 0.150054f
C2975 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n18 VGND 0.165748f
C2976 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t12 VGND 0.104738f
C2977 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t11 VGND 0.104738f
C2978 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n19 VGND 0.165748f
C2979 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t15 VGND 0.104738f
C2980 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t8 VGND 0.104738f
C2981 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n20 VGND 0.165748f
C2982 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n21 VGND 0.150054f
C2983 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t9 VGND 0.104738f
C2984 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.t14 VGND 0.104738f
C2985 SUNSAR_SAR8B_CV_0.XDAC1.CP<8>.n22 VGND 0.280081f
C2986 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.D VGND 0.103605f
C2987 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n2 VGND 0.102978f
C2988 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n5 VGND 0.102978f
C2989 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n6 VGND 0.102978f
C2990 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n7 VGND 0.102978f
C2991 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n10 VGND 0.185977f
C2992 SUNSAR_SAR8B_CV_0.XA0.XA1.CHL_OP.n11 VGND 0.431108f
C2993 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n4 VGND 0.363706f
C2994 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n5 VGND 0.312642f
C2995 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n44 VGND 0.196567f
C2996 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n45 VGND 0.532249f
C2997 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n46 VGND 0.381443f
C2998 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n47 VGND 0.381443f
C2999 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n48 VGND 0.381443f
C3000 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n49 VGND 0.381443f
C3001 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n50 VGND 0.381443f
C3002 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n51 VGND 1.20204f
C3003 SUNSAR_CAPT8B_CV_0.CK_SAMPLE VGND 0.140438f
C3004 SUNSAR_SAR8B_CV_0.CK_SAMPLE.n52 VGND 0.787423f
C3005 SUNSAR_SAR8B_CV_0.D<3>.n4 VGND 0.159682f
C3006 SUNSAR_SAR8B_CV_0.D<3>.n5 VGND 0.142236f
C3007 SUNSAR_SAR8B_CV_0.D<3>.n6 VGND 0.568748f
C3008 SUNSAR_SAR8B_CV_0.D<3>.n7 VGND 0.5979f
C3009 SUNSAR_SAR8B_CV_0.D<3>.n8 VGND 0.123392f
C3010 SUNSAR_SAR8B_CV_0.D<3>.t9 VGND 0.116391f
C3011 SUNSAR_SAR8B_CV_0.D<3>.t11 VGND 0.112495f
C3012 SUNSAR_SAR8B_CV_0.D<3>.n10 VGND 0.290304f
C3013 SUNSAR_SAR8B_CV_0.D<3>.n12 VGND 0.566063f
C3014 SUNSAR_SAR8B_CV_0.D<3>.n13 VGND 0.684236f
C3015 SUNSAR_SAR8B_CV_0.D<3>.n14 VGND 2.1527f
C3016 SUNSAR_SAR8B_CV_0.D<3>.n15 VGND 2.48294f
C3017 SUNSAR_SAR8B_CV_0.D<3>.n16 VGND 2.65688f
C3018 SUNSAR_SAR8B_CV_0.D<3>.n24 VGND 0.146146f
C3019 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n4 VGND 0.113645f
C3020 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n5 VGND 0.101228f
C3021 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n6 VGND 0.404773f
C3022 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n7 VGND 0.425521f
C3023 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n9 VGND 0.22637f
C3024 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n10 VGND 0.285936f
C3025 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n11 VGND 0.285936f
C3026 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n12 VGND 0.285936f
C3027 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n13 VGND 0.285936f
C3028 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n14 VGND 1.83195f
C3029 SUNSAR_SAR8B_CV_0.XDAC1.CP<9>.n18 VGND 0.105641f
C3030 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n0 VGND 0.181013f
C3031 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n1 VGND 0.163874f
C3032 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t12 VGND 0.114384f
C3033 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t9 VGND 0.114384f
C3034 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n2 VGND 0.163874f
C3035 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n3 VGND 0.181013f
C3036 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t11 VGND 0.114384f
C3037 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t13 VGND 0.114384f
C3038 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n4 VGND 0.181013f
C3039 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t15 VGND 0.114384f
C3040 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t10 VGND 0.114384f
C3041 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n5 VGND 0.181013f
C3042 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n6 VGND 0.163874f
C3043 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t8 VGND 0.114384f
C3044 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.t14 VGND 0.114384f
C3045 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n7 VGND 0.145729f
C3046 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n8 VGND 0.171979f
C3047 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n9 VGND 4.05039f
C3048 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n10 VGND 5.3182f
C3049 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n13 VGND 0.192843f
C3050 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n15 VGND 0.110769f
C3051 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n16 VGND 0.153617f
C3052 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n18 VGND 0.153617f
C3053 SUNSAR_SAR8B_CV_0.XDAC2.CP<7>.n20 VGND 0.110769f
C3054 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.D VGND 0.152072f
C3055 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n0 VGND 0.111648f
C3056 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n1 VGND 0.1444f
C3057 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n2 VGND 0.130728f
C3058 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n3 VGND 0.130728f
C3059 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n4 VGND 0.1444f
C3060 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n5 VGND 0.1444f
C3061 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n6 VGND 0.1444f
C3062 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n7 VGND 0.130728f
C3063 SUNSAR_SAR8B_CV_0.XA1.XA1.CHL_ON.n8 VGND 0.176497f
C3064 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n5 VGND 0.114683f
C3065 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n7 VGND 0.10592f
C3066 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n9 VGND 0.161605f
C3067 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n10 VGND 0.321333f
C3068 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n14 VGND 0.178039f
C3069 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n15 VGND 0.295079f
C3070 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n19 VGND 0.161605f
C3071 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n20 VGND 0.321333f
C3072 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n24 VGND 0.178039f
C3073 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n25 VGND 0.295079f
C3074 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n29 VGND 0.161605f
C3075 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n30 VGND 0.321333f
C3076 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n34 VGND 0.178039f
C3077 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n35 VGND 0.295079f
C3078 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n39 VGND 0.161605f
C3079 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n40 VGND 0.321333f
C3080 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n44 VGND 0.656088f
C3081 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n45 VGND 0.626911f
C3082 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n46 VGND 0.626911f
C3083 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n47 VGND 0.626911f
C3084 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n48 VGND 0.626911f
C3085 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n49 VGND 0.658494f
C3086 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n53 VGND 0.178039f
C3087 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n54 VGND 0.295079f
C3088 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n56 VGND 0.411545f
C3089 SUNSAR_SAR8B_CV_0.XA0.CMP_OP.n57 VGND 0.245301f
C3090 SUNSAR_SAR8B_CV_0.XA20.XA1.MN6.G VGND 0.156149f
C3091 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n0 VGND 0.134803f
C3092 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n2 VGND 0.124342f
C3093 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n3 VGND 0.11383f
C3094 SUNSAR_SAR8B_CV_0.XA20.XA2.MN0.G VGND 0.119554f
C3095 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n4 VGND 0.399365f
C3096 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n5 VGND 0.134803f
C3097 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n7 VGND 0.124342f
C3098 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n8 VGND 0.11383f
C3099 SUNSAR_SAR8B_CV_0.XA20.XA3.MN0.G VGND 0.119554f
C3100 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n9 VGND 0.628447f
C3101 SUNSAR_SAR8B_CV_0.XA20.XA4.MN6.G VGND 0.290869f
C3102 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n10 VGND 0.15997f
C3103 SUNSAR_SAR8B_CV_0.XA20.XA1.CK.n11 VGND 0.102716f
C3104 SUNSAR_SAR8B_CV_0.XA20.XA9.MP0.D VGND 0.129257f
C3105 SUNSAR_SAR8B_CV_0.XA4.CP0.n3 VGND 0.110522f
C3106 SUNSAR_SAR8B_CV_0.XA4.CP0.n4 VGND 0.100058f
C3107 SUNSAR_SAR8B_CV_0.XA4.CP0.n5 VGND 0.100058f
C3108 SUNSAR_SAR8B_CV_0.XA4.CP0.n6 VGND 0.110522f
C3109 SUNSAR_SAR8B_CV_0.XA4.CP0.n7 VGND 0.110522f
C3110 SUNSAR_SAR8B_CV_0.XA4.CP0.n8 VGND 0.110522f
C3111 SUNSAR_SAR8B_CV_0.XA4.CP0.n9 VGND 0.100058f
C3112 SUNSAR_SAR8B_CV_0.XA4.CP0.n10 VGND 0.186761f
C3113 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.D VGND 0.103605f
C3114 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n2 VGND 0.102978f
C3115 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n5 VGND 0.102978f
C3116 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n6 VGND 0.102978f
C3117 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n7 VGND 0.102978f
C3118 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n10 VGND 0.185977f
C3119 SUNSAR_SAR8B_CV_0.XA4.XA1.CHL_OP.n11 VGND 0.431108f
C3120 VPWR.n0 VGND 0.458144f
C3121 VPWR.n26 VGND 0.282765f
C3122 VPWR.n27 VGND 0.360086f
C3123 VPWR.n221 VGND 0.284937f
C3124 VPWR.n222 VGND 0.340104f
C3125 VPWR.n253 VGND 0.284937f
C3126 VPWR.t71 VGND 5.37559f
C3127 VPWR.n309 VGND 0.239591f
C3128 VPWR.n344 VGND 0.129734f
C3129 VPWR.n368 VGND 0.281679f
C3130 VPWR.n392 VGND 0.281679f
C3131 VPWR.n433 VGND 0.239591f
C3132 VPWR.t102 VGND 5.37559f
C3133 VPWR.t9 VGND 5.37559f
C3134 VPWR.n598 VGND 5.60932f
C3135 VPWR.n609 VGND 0.240656f
C3136 VPWR.n635 VGND 0.144785f
C3137 VPWR.n645 VGND 0.361389f
C3138 VPWR.n646 VGND 0.361389f
C3139 VPWR.n647 VGND 0.106426f
C3140 VPWR.n679 VGND 0.283851f
C3141 VPWR.n722 VGND 0.283851f
C3142 VPWR.n763 VGND 0.239591f
C3143 VPWR.t17 VGND 5.37559f
C3144 VPWR.t94 VGND 5.37559f
C3145 VPWR.n928 VGND 5.60932f
C3146 VPWR.n939 VGND 0.240656f
C3147 VPWR.n965 VGND 0.142861f
C3148 VPWR.n966 VGND 0.360086f
C3149 VPWR.n967 VGND 0.360086f
C3150 VPWR.n968 VGND 0.106426f
C3151 VPWR.n991 VGND 0.112186f
C3152 VPWR.n995 VGND 0.112186f
C3153 VPWR.t45 VGND 0.245571f
C3154 VPWR.n1002 VGND 0.112186f
C3155 VPWR.n1003 VGND 0.112186f
C3156 VPWR.n1010 VGND 0.213259f
C3157 VPWR.n1032 VGND 0.112186f
C3158 VPWR.n1033 VGND 0.112186f
C3159 VPWR.n1034 VGND 0.112186f
C3160 VPWR.n1041 VGND 0.112186f
C3161 VPWR.n1043 VGND 0.112186f
C3162 VPWR.n1044 VGND 0.112186f
C3163 VPWR.n1053 VGND 0.112186f
C3164 VPWR.n1054 VGND 0.112186f
C3165 VPWR.n1060 VGND 0.112186f
C3166 VPWR.n1061 VGND 0.112186f
C3167 VPWR.t179 VGND 0.245571f
C3168 VPWR.n1068 VGND 2.92997f
C3169 VPWR.n1081 VGND 0.112186f
C3170 VPWR.n1085 VGND 0.112186f
C3171 VPWR.t137 VGND 0.245571f
C3172 VPWR.n1098 VGND 0.112186f
C3173 VPWR.n1099 VGND 0.112186f
C3174 VPWR.n1108 VGND 0.197833f
C3175 VPWR.n1134 VGND 0.112186f
C3176 VPWR.n1135 VGND 0.112186f
C3177 VPWR.n1136 VGND 0.112186f
C3178 VPWR.n1143 VGND 0.112186f
C3179 VPWR.n1145 VGND 0.112186f
C3180 VPWR.n1146 VGND 0.112186f
C3181 VPWR.n1155 VGND 0.112186f
C3182 VPWR.n1156 VGND 0.112186f
C3183 VPWR.n1162 VGND 0.112186f
C3184 VPWR.n1163 VGND 0.112186f
C3185 VPWR.t141 VGND 0.245571f
C3186 VPWR.n1172 VGND 0.885485f
C3187 VPWR.n1173 VGND 2.05652f
C3188 VPWR.n1174 VGND 0.290888p
C3189 VPWR.t21 VGND 5.37559f
C3190 VPWR.n1230 VGND 0.239591f
C3191 VPWR.n1273 VGND 0.282765f
C3192 VPWR.n1274 VGND 0.360086f
C3193 VPWR.n1275 VGND 0.143825f
C3194 VPWR.n1300 VGND 0.240656f
C3195 VPWR.t6 VGND 5.37559f
C3196 VPWR.n1430 VGND 5.60932f
C3197 VPWR.n1445 VGND 0.106426f
C3198 VPWR.n1451 VGND 1.09535f
C3199 VPWR.t98 VGND 0.245571f
C3200 VPWR.n1457 VGND 0.112186f
C3201 VPWR.n1465 VGND 0.112186f
C3202 VPWR.n1472 VGND 0.112186f
C3203 VPWR.n1480 VGND 0.112186f
C3204 VPWR.n1487 VGND 0.112186f
C3205 VPWR.t186 VGND 0.245571f
C3206 VPWR.n1615 VGND 0.112186f
C3207 VPWR.n1616 VGND 0.112186f
C3208 VPWR.n1631 VGND 0.112186f
C3209 VPWR.n1632 VGND 0.112186f
C3210 VPWR.n1647 VGND 0.112186f
C3211 VPWR.n1648 VGND 0.112186f
C3212 VPWR.n1656 VGND 0.112186f
C3213 VPWR.n1670 VGND 0.112186f
C3214 VPWR.n1686 VGND 0.112186f
C3215 VPWR.n1702 VGND 0.112186f
C3216 VPWR.n1703 VGND 0.112186f
C3217 VPWR.n1704 VGND 0.112186f
C3218 VPWR.n1710 VGND 0.112186f
C3219 VPWR.n1711 VGND 0.112186f
C3220 VPWR.n1718 VGND 0.112186f
C3221 VPWR.n1719 VGND 0.112186f
C3222 VPWR.n1720 VGND 0.112186f
C3223 VPWR.n1733 VGND 0.252405f
C3224 VPWR.n1736 VGND 1.39961f
C3225 VPWR.n1765 VGND 0.240656f
C3226 VPWR.t27 VGND 5.37559f
C3227 VPWR.n1895 VGND 5.60932f
C3228 VPWR.n1910 VGND 0.106426f
C3229 VPWR.n1911 VGND 0.361389f
C3230 VPWR.t86 VGND 0.245571f
C3231 VPWR.n1922 VGND 0.112186f
C3232 VPWR.t500 VGND 0.245571f
C3233 VPWR.n1927 VGND 0.112186f
C3234 VPWR.n1928 VGND 0.112186f
C3235 VPWR.n1934 VGND 0.112186f
C3236 VPWR.n1935 VGND 0.112186f
C3237 VPWR.n1936 VGND 0.112186f
C3238 VPWR.t604 VGND 14.895999f
C3239 VPWR.t602 VGND 7.64907f
C3240 VPWR.n1962 VGND 7.41988f
C3241 VPWR.t607 VGND 7.64907f
C3242 VPWR.n1963 VGND 7.34563f
C3243 VPWR.t608 VGND 7.64907f
C3244 VPWR.n1964 VGND 7.34563f
C3245 VPWR.t606 VGND 7.64907f
C3246 VPWR.n1965 VGND 7.34563f
C3247 VPWR.t603 VGND 7.64907f
C3248 VPWR.n1966 VGND 7.34563f
C3249 VPWR.t605 VGND 7.64907f
C3250 VPWR.n1967 VGND 7.34563f
C3251 VPWR.t610 VGND 7.64907f
C3252 VPWR.n1968 VGND 7.34563f
C3253 VPWR.t609 VGND 7.64907f
C3254 VPWR.n1969 VGND 7.535f
C3255 VPWR.n1970 VGND 1.34856f
C3256 VPWR.n1971 VGND 1.53265f
C3257 VPWR.n2017 VGND 0.112186f
C3258 VPWR.t289 VGND 0.245571f
C3259 VPWR.n2022 VGND 0.112186f
C3260 VPWR.n2023 VGND 0.112186f
C3261 VPWR.n2030 VGND 0.112186f
C3262 VPWR.n2032 VGND 0.112186f
C3263 VPWR.n2033 VGND 0.112186f
C3264 VPWR.n2040 VGND 0.112186f
C3265 VPWR.n2041 VGND 0.112186f
C3266 VPWR.n2042 VGND 0.112186f
C3267 VPWR.n2043 VGND 0.112186f
C3268 VPWR.n2050 VGND 0.112186f
C3269 VPWR.n2052 VGND 0.112186f
C3270 VPWR.n2059 VGND 0.112186f
C3271 VPWR.n2060 VGND 0.112186f
C3272 VPWR.n2061 VGND 0.112186f
C3273 VPWR.n2062 VGND 0.112186f
C3274 VPWR.n2068 VGND 0.112186f
C3275 VPWR.n2069 VGND 0.112186f
C3276 VPWR.t30 VGND 0.245571f
C3277 VPWR.n2078 VGND 0.236366f
C3278 VPWR.t60 VGND 2.02122f
C3279 VPWR.t196 VGND 2.02122f
C3280 VPWR.n2134 VGND 2.1091f
C3281 VPWR.n2143 VGND 0.227214f
C3282 VPWR.n2144 VGND 0.229402f
C3283 VPWR.t75 VGND 2.02122f
C3284 VPWR.t106 VGND 2.02122f
C3285 VPWR.n2200 VGND 2.1091f
C3286 VPWR.n2209 VGND 0.227214f
C3287 VPWR.n2210 VGND 0.231229f
C3288 VPWR.t145 VGND 2.02122f
C3289 VPWR.t153 VGND 2.02122f
C3290 VPWR.n2266 VGND 2.1091f
C3291 VPWR.n2275 VGND 0.227214f
C3292 VPWR.n2276 VGND 0.229402f
C3293 VPWR.t56 VGND 2.02122f
C3294 VPWR.t165 VGND 2.02122f
C3295 VPWR.n2332 VGND 2.1091f
C3296 VPWR.n2341 VGND 0.141164f
C3297 VPWR.n2343 VGND 0.12684f
C3298 VPWR.n2345 VGND 6.18132f
C3299 VPWR.n2346 VGND 0.167477p
C3300 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n0 VGND 0.310531f
C3301 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n1 VGND 6.31117f
C3302 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n2 VGND 0.12659f
C3303 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n3 VGND 0.111901f
C3304 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n4 VGND 0.175637f
C3305 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n5 VGND 0.243577f
C3306 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n6 VGND 0.12659f
C3307 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n7 VGND 0.174127f
C3308 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n8 VGND 0.250629f
C3309 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n9 VGND 0.111901f
C3310 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n11 VGND 0.25984f
C3311 SUNSAR_SAR8B_CV_0.XDAC2.CP<6>.n12 VGND 0.484086f
C3312 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n0 VGND 0.23337f
C3313 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n1 VGND 0.211274f
C3314 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t9 VGND 0.147469f
C3315 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t11 VGND 0.147469f
C3316 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n2 VGND 0.211274f
C3317 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n3 VGND 0.23337f
C3318 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t15 VGND 0.147469f
C3319 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t14 VGND 0.147469f
C3320 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n4 VGND 0.23337f
C3321 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t13 VGND 0.147469f
C3322 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t12 VGND 0.147469f
C3323 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n5 VGND 0.23337f
C3324 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n6 VGND 0.211274f
C3325 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t10 VGND 0.147469f
C3326 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.t8 VGND 0.147469f
C3327 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n7 VGND 0.211274f
C3328 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n9 VGND 0.248621f
C3329 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n10 VGND 4.5573f
C3330 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n12 VGND 0.110687f
C3331 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n13 VGND 0.203784f
C3332 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n14 VGND 0.109459f
C3333 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n15 VGND 0.102929f
C3334 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n16 VGND 0.19805f
C3335 SUNSAR_SAR8B_CV_0.XDAC1.CP<6>.n18 VGND 0.142809f
.ends

