* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[1] uio_oe[2]
*+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[1] uio_out[2] uio_out[3]
*+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7] uio_oe[0] uo_out[6]
*+ ui_in[0] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3] uio_out[0]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA0.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=243.9396 ps=1.2855k w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=247.698 ps=1.29678k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R5 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VPWR tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X51 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X52 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X56 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.36 w=1.08 l=0.18
X58 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X62 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X63 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X65 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X66 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X72 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X74 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X76 VGND SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X77 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X78 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X79 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X87 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X88 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X90 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X95 VGND SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X96 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X97 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X98 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X99 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X100 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X101 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X106 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X107 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X108 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R8 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X114 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CNO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X115 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X116 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X118 VGND SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X119 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R9 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X120 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X121 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X122 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X124 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X125 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R11 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X130 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X131 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X132 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X134 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X135 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X136 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X137 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CNO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X140 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R12 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X144 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X146 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X147 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X148 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X149 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X150 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R13 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X155 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X158 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R14 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X160 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X163 VGND SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X166 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X167 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 VPWR SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R15 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X169 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X174 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X175 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X176 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X177 VGND SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R16 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X178 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X181 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X182 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 VPWR SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X185 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X186 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X188 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X193 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X194 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X195 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X198 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X199 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R17 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X201 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X205 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X206 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X207 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X208 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X209 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X210 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X211 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R18 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X212 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X213 VGND SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X214 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X215 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X216 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X217 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R19 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X220 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X221 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X222 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X223 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X224 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X225 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X226 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X227 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X228 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X229 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X230 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X232 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X233 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X235 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X236 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X237 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X239 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X246 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X253 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X255 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X263 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X266 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X268 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 VPWR SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X270 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X275 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X276 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X278 uio_oe[0] tt_um_TT06_SAR_done_0.x4.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R22 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X280 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X282 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X284 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R23 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X286 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X292 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R24 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X294 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X300 uio_out[0] tt_um_TT06_SAR_done_0.x3.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X307 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X308 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X309 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X310 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X311 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X312 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X313 VPWR SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X314 VGND SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA6.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X316 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X318 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R25 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R26 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X321 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X322 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X324 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
D0 VGND ui_in[0] sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X325 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X328 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R27 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X333 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X337 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X338 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X339 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X341 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X342 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X344 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X346 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X347 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X348 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X349 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X351 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X352 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X353 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X355 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X359 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X360 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X363 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X364 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X365 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X366 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X368 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X369 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X370 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X371 VGND SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X372 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R29 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X373 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X374 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X375 VPWR SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X376 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R30 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X377 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X378 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X379 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X381 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X382 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X384 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X385 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X386 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X387 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X389 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X390 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X391 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X393 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R31 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X394 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X395 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X400 VPWR SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R32 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X402 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X404 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X407 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA4.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X410 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R34 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X413 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X414 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X416 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X417 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X418 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X419 SUNSAR_SAR8B_CV_0.XA20.XA11.Y tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X420 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X421 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X422 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X423 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R35 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X424 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X425 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X426 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X427 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X428 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X429 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X430 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X431 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X432 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X433 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X434 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X435 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X436 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X437 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R36 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X440 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X441 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X442 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X443 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R37 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X447 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X449 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X450 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X452 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X453 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X454 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X455 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X457 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X458 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X459 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X462 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X463 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R38 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X464 VPWR SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X465 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X468 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X470 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X471 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X472 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X473 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X474 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 VGND SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X477 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X478 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X479 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X480 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X481 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X482 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X486 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 VGND SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R41 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X489 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X491 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X492 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X493 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X494 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
D1 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X496 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X498 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X499 VPWR SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X500 VGND SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R42 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X501 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X502 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X503 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X505 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X506 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X508 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R43 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X510 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X511 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X512 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X513 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X514 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X515 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R44 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X516 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X517 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X519 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X520 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X521 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X522 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X524 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X525 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X526 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X527 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X528 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X530 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X532 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X533 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X536 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X537 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X540 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X541 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X544 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X545 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X548 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X553 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X554 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X557 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X558 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X560 VGND SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X561 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X562 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X563 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X564 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X565 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 VPWR SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X567 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X568 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X570 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X571 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X572 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X573 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X574 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R46 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X575 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_CAPT8B_CV_0.XA7.MP0.G SUNSAR_CAPT8B_CV_0.XA7.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X578 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X579 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X580 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X581 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X582 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X583 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S SUNSAR_CAPT8B_CV_0.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X584 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X587 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X588 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X589 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X590 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X591 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X592 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X593 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X594 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X595 VGND SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X596 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X598 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X601 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X602 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R48 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X603 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X604 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X605 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X606 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X609 VGND SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X610 VGND SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X613 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X614 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X616 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X618 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X619 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X621 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X624 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X626 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X631 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X637 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X640 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R49 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X642 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X644 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X645 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X647 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X648 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X649 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X650 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X652 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X653 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R51 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X654 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X656 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X657 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X658 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X661 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X663 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X664 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X665 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X666 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R53 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X667 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X668 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X669 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X670 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X674 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X675 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X676 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 VGND SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X680 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X681 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X682 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X683 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X684 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X685 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X686 VPWR SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X687 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X688 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X690 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R54 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X691 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X693 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X694 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X695 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R55 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X696 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X697 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X699 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X700 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X701 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X704 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X705 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X706 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X707 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X709 VGND tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X710 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X713 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X714 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X715 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X716 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X717 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X718 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X719 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X720 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X721 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X722 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R57 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X726 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X727 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X728 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X729 VGND SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X730 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R58 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X731 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X732 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 VPWR SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X734 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X735 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X738 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X740 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X741 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R59 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
R60 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X742 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X745 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X746 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X747 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X749 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R61 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X751 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R62 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X752 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X753 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X754 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X755 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X759 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X760 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X762 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X763 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X765 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X766 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X767 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X768 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 VGND SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CNO VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R64 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X770 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X771 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X773 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X774 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 VPWR SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X777 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X778 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X779 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X780 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X782 VGND SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CNO VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R65 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X783 VGND SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X786 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X787 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X788 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R67 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X790 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X791 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X792 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X793 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X798 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X800 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X802 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X809 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X810 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X813 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X814 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X816 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X817 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X818 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X819 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X821 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X822 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X823 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X824 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X825 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X828 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X829 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X830 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X831 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X832 VPWR SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X833 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X834 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X835 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X836 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X837 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X838 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X839 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R68 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X842 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X843 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X844 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X845 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X846 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X847 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X848 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X849 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X850 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X851 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X852 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X853 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X854 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X855 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X856 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X858 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X859 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X862 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X864 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X867 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X868 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VGND SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X872 VPWR SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X873 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X874 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X875 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X876 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X878 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X879 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X883 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X884 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X886 VGND SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X887 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X890 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X892 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R70 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X893 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X894 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X895 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X896 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X897 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X899 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X901 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R71 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X902 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X903 VGND SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X905 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R72 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X906 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X909 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X910 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R73 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X911 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X912 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X913 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X914 tt_um_TT06_SAR_done_0.x4.MP0.G tt_um_TT06_SAR_done_0.x4.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X915 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X917 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R74 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X918 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X920 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X923 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X924 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X925 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X926 VPWR SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X927 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X928 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X929 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R75 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X930 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X931 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X932 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X933 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X934 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X935 uio_out[0] tt_um_TT06_SAR_done_0.x3.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X936 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X937 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X939 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X940 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X941 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X942 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X943 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R76 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X944 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X945 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X946 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X947 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R77 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X948 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X949 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X950 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X951 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X953 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X954 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X955 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X957 VPWR SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X959 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X961 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X962 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R78 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X963 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X964 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X965 VGND SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA2.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X967 VGND SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 TIE_L SUNSAR_CAPT8B_CV_0.XA7.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X970 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X971 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X972 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X974 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R79 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X975 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X976 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X978 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X980 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X982 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X984 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X985 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X986 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X987 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X988 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X993 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R80 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X994 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X995 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X997 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X999 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
D2 VGND clk sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X1000 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1001 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1002 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1004 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1005 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R81 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1008 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1013 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R82 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X1014 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R83 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1016 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1018 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1019 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1020 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1021 VGND SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1022 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 VPWR SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1025 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1033 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1034 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1035 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1036 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1037 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1038 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1039 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1040 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1041 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1042 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1043 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1044 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1045 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1046 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1047 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1048 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1049 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1050 VGND tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1051 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1052 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1053 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1054 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.098057f
C1 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.010609f
C2 SUNSAR_SAR8B_CV_0.D<4> a_10170_34716# 0.070775f
C3 SUNSAR_CAPT8B_CV_0.XD09.QN TIE_L1 0.012277f
C4 a_8802_30316# VPWR 0.404384f
C5 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_2630_41352# 0.080002f
C6 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_21422_41880# 0.031087f
C7 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_11322_35068# 0.129098f
C8 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.019709f
C9 a_2610_35420# SUNSAR_SAR8B_CV_0.XA0.DONE 0.030547f
C10 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.143554f
C11 a_15210_27500# VPWR 0.382397f
C12 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.34399f
C13 a_3782_44168# SUNSAR_CAPT8B_CV_0.XB07.QN 0.066018f
C14 SUNSAR_SAR8B_CV_0.XA3.XA2.A a_10170_30316# 0.127528f
C15 a_20270_41880# VPWR 0.395781f
C16 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S 0.011178f
C17 SUNSAR_SAR8B_CV_0.D<2> a_15230_41352# 0.06659f
C18 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.097975f
C19 a_20250_32956# VPWR 0.433941f
C20 a_17730_27852# a_17730_27500# 0.010937f
C21 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.2165f
C22 SUNSAR_SAR8B_CV_0.EN a_18882_29612# 0.143959f
C23 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.062692f
C24 a_11142_3334# a_11142_2982# 0.010937f
C25 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B a_16542_2982# 0.011407f
C26 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VPWR 1.06875f
C27 a_17730_32076# SUNSAR_SAR8B_CV_0.XA6.CN1 0.06949f
C28 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C29 a_10190_42760# VPWR 0.391454f
C30 SUNSAR_SAR8B_CV_0.EN tt_um_TT06_SAR_done_0.DONE 0.131506f
C31 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S 0.067572f
C32 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S 0.055627f
C33 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.744161f
C34 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N a_7650_28908# 0.060353f
C35 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.021955f
C36 SUNSAR_SAR8B_CV_0.SARP a_13950_5094# 0.047906f
C37 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.201839f
C38 a_2610_36300# SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.068275f
C39 SUNSAR_SAR8B_CV_0.EN a_3762_30316# 0.077363f
C40 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 5.71192f
C41 SUNSAR_CAPT8B_CV_0.XI14.XA7.C uio_oe[0] 0.010428f
C42 SUNSAR_SAR8B_CV_0.SARP VPWR 0.155428f
C43 a_5150_43288# uo_out[6] 0.071088f
C44 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.093524f
C45 a_17730_35068# SUNSAR_SAR8B_CV_0.XA7.EN 0.067588f
C46 SUNSAR_SAR8B_CV_0.EN a_10170_27500# 0.073293f
C47 a_9990_4566# VPWR 0.413433f
C48 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18126_2928# 0.024512f
C49 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.723061f
C50 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA20.CPO 0.058451f
C51 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.103734f
C52 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_20270_41880# 0.071088f
C53 VPWR uio_oe[0] 1.67769f
C54 uo_out[3] uo_out[2] 0.109993f
C55 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.318734f
C56 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S 0.050207f
C57 a_18902_41000# tt_um_TT06_SAR_done_0.DONE 0.066018f
C58 a_8822_41000# a_8822_40648# 0.010937f
C59 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1615f
C60 a_20250_35420# VPWR 0.39661f
C61 a_3762_36828# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.066018f
C62 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.02121f
C63 a_13862_44168# uo_out[3] 0.041694f
C64 a_20250_27148# a_20250_26796# 0.010937f
C65 a_20270_44168# VPWR 0.340085f
C66 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S 0.010488f
C67 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_41880# 0.100592f
C68 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S 0.021211f
C69 SUNSAR_SAR8B_CV_0.XA3.XA9.B a_11322_35068# 0.011912f
C70 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_10170_35068# 0.089492f
C71 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA1.EN 0.051732f
C72 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.176792f
C73 a_13842_27500# VPWR 0.382189f
C74 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.028261f
C75 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.024085f
C76 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.193521f
C77 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.209683f
C78 TIE_L SUNSAR_CAPT8B_CV_0.XC08.QN 0.013096f
C79 a_2630_44168# SUNSAR_CAPT8B_CV_0.XB07.QN 0.071093f
C80 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.011514f
C81 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_3762_29612# 0.023777f
C82 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.204048f
C83 a_18902_41880# VPWR 0.395781f
C84 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S 0.150467f
C85 a_20250_36300# VPWR 0.395776f
C86 a_18882_37532# a_18882_37180# 0.010937f
C87 a_18882_32956# VPWR 0.436368f
C88 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_5150_42408# 0.076129f
C89 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_6302_42408# 0.098561f
C90 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.12241f
C91 a_11322_35948# SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.071154f
C92 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA20.CNO 0.065777f
C93 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S 0.073313f
C94 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B a_9990_2630# 0.015402f
C95 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR 0.137646f
C96 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_22770_34540# 0.103065f
C97 a_23922_34892# a_23922_34540# 0.010937f
C98 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.133602f
C99 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_16362_31196# 0.010411f
C100 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.012782f
C101 a_8822_42760# VPWR 0.391454f
C102 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_16382_43288# 0.028213f
C103 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S 0.030221f
C104 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.649845f
C105 ui_in[4] ui_in[3] 0.023797f
C106 a_15210_37180# VPWR 0.474036f
C107 SUNSAR_SAR8B_CV_0.XA20.CPO a_21402_28556# 0.014699f
C108 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_3762_27500# 0.033843f
C109 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_13842_27852# 0.028807f
C110 a_2610_28204# a_2610_27852# 0.010937f
C111 SUNSAR_SAR8B_CV_0.EN a_2610_30316# 0.078848f
C112 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80604f
C113 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S uo_out[0] 0.01183f
C114 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S 0.089305f
C115 a_6282_35068# a_6282_34716# 0.010937f
C116 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA2.EN 1.2771f
C117 SUNSAR_SAR8B_CV_0.EN a_8802_27500# 0.071722f
C118 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VPWR 0.452478f
C119 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18054_2928# 0.024512f
C120 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.031784f
C121 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.046398f
C122 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3a.A 1.43919f
C123 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.028032f
C124 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.08285f
C125 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S 0.010423f
C126 SUNSAR_CAPT8B_CV_0.XA5.XA2.A a_23942_42408# 0.091063f
C127 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.055045f
C128 VPWR clk 0.644902f
C129 a_8822_43816# SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.069905f
C130 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 0.093019f
C131 a_28727_41011# VPWR 0.468616f
C132 a_17750_41000# tt_um_TT06_SAR_done_0.DONE 0.070731f
C133 a_18882_35420# VPWR 0.39968f
C134 a_11322_28556# SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.066018f
C135 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.010771f
C136 a_2610_36828# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.072629f
C137 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA7.EN 0.439535f
C138 a_12710_44168# uo_out[3] 0.041178f
C139 a_18902_44168# VPWR 0.3405f
C140 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.023976f
C141 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_SAR8B_CV_0.D<4> 0.393055f
C142 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S 0.021266f
C143 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.DONE 0.034185f
C144 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.238862f
C145 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_16382_42760# 0.091344f
C146 SUNSAR_SAR8B_CV_0.XA2.XA2.A a_8802_30316# 0.129098f
C147 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S 0.013533f
C148 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_2610_29612# 0.040867f
C149 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.019336f
C150 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.284482f
C151 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.040976f
C152 SUNSAR_SAR8B_CV_0.SARN a_13950_3334# 0.037937f
C153 a_18882_36300# VPWR 0.399161f
C154 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S 0.050207f
C155 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.075315f
C156 a_16362_27852# a_16362_27500# 0.010937f
C157 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_42408# 0.031125f
C158 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.199693f
C159 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.432466f
C160 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.626084f
C161 a_10170_35948# SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.067588f
C162 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.205884f
C163 a_9990_3334# a_9990_2982# 0.010937f
C164 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VPWR 1.05322f
C165 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C166 a_16362_32076# SUNSAR_SAR8B_CV_0.XA5.CN1 0.06792f
C167 SUNSAR_CAPT8B_CV_0.XA5.B a_22790_41880# 0.017896f
C168 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_15230_43288# 0.082288f
C169 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_16382_43288# 0.067482f
C170 a_23942_43640# SUNSAR_CAPT8B_CV_0.XA6.B 0.066018f
C171 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S 0.044855f
C172 a_13842_37180# VPWR 0.473697f
C173 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.666402f
C174 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA20.CPO 1.15994f
C175 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C176 a_23922_36652# a_23922_36300# 0.010937f
C177 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S uo_out[0] 0.023976f
C178 a_20250_29612# VPWR 0.398044f
C179 a_3782_43288# uo_out[7] 0.073429f
C180 a_13950_5094# a_13950_4742# 0.010937f
C181 a_5150_43288# VPWR 0.394205f
C182 a_16362_35068# SUNSAR_SAR8B_CV_0.XA6.EN 0.066018f
C183 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_3728# 0.172147f
C184 a_23922_33132# SUNSAR_SAR8B_CV_0.XA20.XA3a.A 0.066404f
C185 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.723071f
C186 SUNSAR_CAPT8B_CV_0.XA5.XA2.A a_22790_42408# 0.10248f
C187 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S 0.089305f
C188 VPWR ui_in[0] 2.01351f
C189 uo_out[4] uo_out[3] 0.854997f
C190 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.010898f
C191 a_16382_41000# tt_um_TT06_SAR_done_0.DONE 0.06916f
C192 a_7670_41000# a_7670_40648# 0.010937f
C193 a_10170_28556# SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.071498f
C194 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.303978f
C195 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.098057f
C196 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 6.86675f
C197 a_18882_27148# a_18882_26796# 0.010937f
C198 a_5130_30316# VPWR 0.404384f
C199 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_SAR8B_CV_0.D<4> 0.241356f
C200 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_15230_42760# 0.111734f
C201 TIE_L SUNSAR_CAPT8B_CV_0.XA7.MP0.G 0.029321f
C202 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.011514f
C203 SUNSAR_SAR8B_CV_0.XA2.XA2.A a_7650_30316# 0.089492f
C204 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_28204# 0.016912f
C205 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.064969f
C206 a_17730_37532# a_17730_37180# 0.010937f
C207 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S 0.022425f
C208 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_SAR8B_CV_0.EN 0.176398f
C209 SUNSAR_SAR8B_CV_0.EN a_15210_29612# 0.143959f
C210 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR 0.138148f
C211 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.093415f
C212 a_22770_34892# a_22770_34540# 0.010937f
C213 a_15210_32076# SUNSAR_SAR8B_CV_0.XA5.CN1 0.067588f
C214 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S 0.012065f
C215 ui_in[5] ui_in[4] 0.023797f
C216 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_43288# 0.031221f
C217 a_22790_43640# SUNSAR_CAPT8B_CV_0.XA6.B 0.081836f
C218 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR 0.097407f
C219 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.079557f
C220 SUNSAR_SAR8B_CV_0.D<3> a_13842_33836# 0.011974f
C221 SUNSAR_CAPT8B_CV_0.XI14.XA7.C uo_out[0] 0.245678f
C222 a_18882_29612# VPWR 0.397362f
C223 a_2630_43288# uo_out[7] 0.066268f
C224 a_3782_43288# VPWR 0.394205f
C225 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C226 a_15210_35068# SUNSAR_SAR8B_CV_0.XA6.EN 0.071277f
C227 a_5130_35068# a_5130_34716# 0.010937f
C228 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24678_3728# 0.0666f
C229 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.014291f
C230 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.449584f
C231 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CN1 0.050197f
C232 a_22770_33132# SUNSAR_SAR8B_CV_0.XA20.XA3a.A 0.067588f
C233 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA20.CPO 0.058427f
C234 VPWR uo_out[0] 1.02382f
C235 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S 0.055045f
C236 a_7670_43816# SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.073123f
C237 SUNSAR_SAR8B_CV_0.XA7.EN a_21402_27148# 0.082474f
C238 tt_um_TT06_SAR_done_0.DONE VPWR 8.70939f
C239 a_15230_41000# tt_um_TT06_SAR_done_0.DONE 0.067588f
C240 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.054448f
C241 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.13078f
C242 SUNSAR_SAR8B_CV_0.D<5> a_8802_34716# 0.069204f
C243 SUNSAR_SAR8B_CV_0.XA7.XA12.A a_21402_36828# 0.104051f
C244 a_11342_44168# uo_out[4] 0.040986f
C245 TIE_L uio_out[0] 0.44106f
C246 a_3762_30316# VPWR 0.404384f
C247 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_8802_35068# 0.091063f
C248 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_13862_42408# 0.015723f
C249 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S 0.036491f
C250 SUNSAR_SAR8B_CV_0.XA20.XA11.Y a_22770_35420# 0.034262f
C251 a_10170_27500# VPWR 0.382397f
C252 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.845515f
C253 a_23942_44344# SUNSAR_CAPT8B_CV_0.XA7.MP0.G 0.096614f
C254 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.126354f
C255 a_15230_41880# VPWR 0.395781f
C256 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.SARP 0.122781f
C257 SUNSAR_SAR8B_CV_0.D<3> a_13862_41352# 0.06816f
C258 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S 0.050648f
C259 a_15210_32956# VPWR 0.436368f
C260 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.86675f
C261 a_15210_27852# a_15210_27500# 0.010937f
C262 SUNSAR_SAR8B_CV_0.EN a_13842_29612# 0.143959f
C263 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_16382_42760# 0.031591f
C264 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S 0.073313f
C265 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA20.CNO 0.066242f
C266 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VPWR 1.06875f
C267 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.033352f
C268 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C269 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C270 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.SARP 0.147435f
C271 a_5150_42760# VPWR 0.391454f
C272 SUNSAR_CAPT8B_CV_0.XI14.XA6.A uo_out[0] 0.014139f
C273 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N a_6282_28908# 0.060353f
C274 SUNSAR_SAR8B_CV_0.XA20.CPO a_17730_28556# 0.014592f
C275 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR 0.112858f
C276 a_22770_36652# a_22770_36300# 0.010937f
C277 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 5.80495f
C278 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN uo_out[0] 0.305166f
C279 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.22339f
C280 a_12582_5094# a_12582_4742# 0.010937f
C281 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S 0.055045f
C282 SUNSAR_SAR8B_CV_0.EN a_5130_27500# 0.073293f
C283 a_13950_5446# ua[0] 0.02841f
C284 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR 0.519052f
C285 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18126_3888# 0.024512f
C286 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.723061f
C287 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_21422_42408# 0.113479f
C288 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S 0.089305f
C289 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_18902_41880# 0.072658f
C290 TIE_L1 uio_oe[0] 0.738069f
C291 uo_out[5] uo_out[4] 1.16093f
C292 uo_out[6] uo_out[3] 0.028786f
C293 VPWR uo_out[1] 1.02322f
C294 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S 0.076714f
C295 SUNSAR_SAR8B_CV_0.XA7.EN a_20250_27148# 0.01235f
C296 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S 0.050207f
C297 a_23942_41000# VPWR 0.390915f
C298 a_13862_41000# tt_um_TT06_SAR_done_0.DONE 0.066018f
C299 a_6302_41000# a_6302_40648# 0.010937f
C300 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6519f
C301 a_15210_35420# VPWR 0.39968f
C302 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.012048f
C303 SUNSAR_SAR8B_CV_0.XA7.XA12.A a_20250_36828# 0.089492f
C304 a_10190_44168# uo_out[4] 0.035338f
C305 a_17730_27148# a_17730_26796# 0.010937f
C306 TIE_L uio_oe[0] 1.21913f
C307 a_15230_44168# VPWR 0.340085f
C308 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_7650_35068# 0.127528f
C309 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.145738f
C310 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_18902_41880# 0.099022f
C311 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.437693f
C312 a_8802_27500# VPWR 0.382189f
C313 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.016209f
C314 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN 0.253395f
C315 a_23942_43112# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.066018f
C316 a_22790_44344# SUNSAR_CAPT8B_CV_0.XA7.MP0.G 0.067588f
C317 a_13862_41880# VPWR 0.395781f
C318 SUNSAR_SAR8B_CV_0.XA1.XA2.A a_6282_30316# 0.091063f
C319 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S 0.011494f
C320 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_23922_29964# 0.035145f
C321 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_28204# 0.017441f
C322 SUNSAR_SAR8B_CV_0.D<3> a_12710_41352# 0.077864f
C323 SUNSAR_SAR8B_CV_0.XA20.CPO a_21402_27852# 0.073814f
C324 a_15210_36300# VPWR 0.398846f
C325 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S 0.050207f
C326 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.030459f
C327 a_16362_37532# a_16362_37180# 0.010937f
C328 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.074964f
C329 a_13842_32956# VPWR 0.436368f
C330 SUNSAR_CAPT8B_CV_0.XA6.B a_22790_43112# 0.012045f
C331 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.062692f
C332 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_42760# 0.031082f
C333 a_23922_28556# VPWR 0.499441f
C334 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.11536f
C335 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S 0.028026f
C336 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.03027f
C337 a_13842_32076# SUNSAR_SAR8B_CV_0.XA4.CN1 0.066018f
C338 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_12690_31196# 0.010411f
C339 a_3782_42760# VPWR 0.391454f
C340 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S 0.012065f
C341 ui_in[6] ui_in[5] 0.023797f
C342 a_10170_37180# VPWR 0.474068f
C343 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N a_5130_28908# 0.023475f
C344 SUNSAR_SAR8B_CV_0.XA20.CPO a_16362_28556# 0.014652f
C345 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_15390_2630# 0.011753f
C346 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR 0.112858f
C347 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S 0.050207f
C348 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S 0.078539f
C349 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.118152f
C350 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.38977f
C351 SUNSAR_CAPT8B_CV_0.XH13.XA7.C uio_oe[0] 0.010428f
C352 a_11142_4918# SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.098163f
C353 a_13842_35068# SUNSAR_SAR8B_CV_0.XA5.EN 0.069707f
C354 a_3762_35068# a_3762_34716# 0.010937f
C355 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S 0.089305f
C356 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S 0.026506f
C357 SUNSAR_SAR8B_CV_0.EN a_3762_27500# 0.071936f
C358 a_16542_4918# VPWR 0.470354f
C359 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18054_3888# 0.024512f
C360 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.014291f
C361 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.449584f
C362 SUNSAR_SAR8B_CV_0.XA7.CP0 a_21402_32956# 0.102695f
C363 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_20270_42408# 0.08955f
C364 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.055045f
C365 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_17750_41880# 0.066018f
C366 VPWR uo_out[2] 1.02322f
C367 m4_11102_44892# uio_oe[0] 0.024961f
C368 uo_out[6] uo_out[4] 0.843602f
C369 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.093019f
C370 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_27148# 0.010025f
C371 a_12710_41000# tt_um_TT06_SAR_done_0.DONE 0.070731f
C372 a_13842_35420# VPWR 0.39968f
C373 a_8802_28556# SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.069927f
C374 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.352238f
C375 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA6.EN 0.503326f
C376 SUNSAR_SAR8B_CV_0.XA20.CPO VPWR 6.88568f
C377 TIE_L clk 0.146712f
C378 a_23942_44344# uio_oe[0] 0.011419f
C379 a_13862_44168# VPWR 0.3405f
C380 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.DONE 0.076485f
C381 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.023976f
C382 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_41880# 0.031087f
C383 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> a_15210_33836# 0.101833f
C384 a_22790_43112# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.071778f
C385 a_23942_43112# SUNSAR_SAR8B_CV_0.EN 0.033775f
C386 SUNSAR_CAPT8B_CV_0.XA5.B clk 0.210661f
C387 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_4038# 0.067824f
C388 SUNSAR_SAR8B_CV_0.XA1.XA2.A a_5130_30316# 0.127528f
C389 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_22770_29964# 0.023357f
C390 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S 0.011062f
C391 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S 0.010193f
C392 SUNSAR_SAR8B_CV_0.XA20.CPO a_20250_27852# 0.066394f
C393 SUNSAR_SAR8B_CV_0.SARN a_13950_3686# 0.049571f
C394 a_13842_36300# VPWR 0.399161f
C395 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.098006f
C396 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.066778f
C397 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S 0.028011f
C398 a_13842_27852# a_13842_27500# 0.010937f
C399 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.205884f
C400 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.077649f
C401 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.432466f
C402 a_8802_35948# SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.066018f
C403 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 0.626356f
C404 SUNSAR_SAR8B_CV_0.D<0> a_20250_32076# 0.020752f
C405 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_3782_42408# 0.031125f
C406 a_22770_28556# VPWR 0.024886f
C407 a_13950_3686# a_13950_3334# 0.010937f
C408 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.014291f
C409 a_12690_32076# SUNSAR_SAR8B_CV_0.XA4.CN1 0.06949f
C410 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.016112f
C411 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S 0.044855f
C412 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP 0.123668f
C413 a_8802_37180# VPWR 0.473729f
C414 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.023017f
C415 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR 4.23254f
C416 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S 0.064105f
C417 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_10170_27852# 0.028807f
C418 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.073351f
C419 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.170578f
C420 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C421 SUNSAR_SAR8B_CV_0.XA7.XA11.A a_21402_36300# 0.13402f
C422 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S 0.016769f
C423 SUNSAR_CAPT8B_CV_0.XA6.B VPWR 0.868246f
C424 a_15210_29612# VPWR 0.397362f
C425 a_11142_4918# SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H 0.015779f
C426 a_9990_4918# SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.067588f
C427 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S uo_out[1] 0.023976f
C428 a_12690_35068# SUNSAR_SAR8B_CV_0.XA5.EN 0.067588f
C429 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.093524f
C430 SUNSAR_SAR8B_CV_0.EN a_2610_27500# 0.079159f
C431 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_21422_41000# 0.115667f
C432 a_12582_5446# ua[1] 0.02841f
C433 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_4688# 0.172147f
C434 SUNSAR_SAR8B_CV_0.XA7.CP0 a_20250_32956# 0.069193f
C435 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.738983f
C436 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.152052f
C437 VPWR uo_out[3] 1.25759f
C438 m4_10366_44892# uio_oe[0] 0.025321f
C439 uo_out[6] uo_out[5] 0.327382f
C440 uo_out[7] uo_out[4] 0.121648f
C441 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.318734f
C442 a_11342_41000# tt_um_TT06_SAR_done_0.DONE 0.06916f
C443 a_5150_41000# a_5150_40648# 0.010937f
C444 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.027995f
C445 a_7650_28556# SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.067588f
C446 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.EN 0.070469f
C447 SUNSAR_SAR8B_CV_0.XA7.CEIN a_21402_36828# 0.073788f
C448 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.033093f
C449 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.054448f
C450 a_22790_44344# uio_oe[0] 0.012146f
C451 a_8822_44168# uo_out[5] 0.036045f
C452 a_23922_30844# VPWR 0.425847f
C453 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 27.1615f
C454 a_16362_27148# a_16362_26796# 0.010937f
C455 SUNSAR_SAR8B_CV_0.XA2.XA9.B a_7650_35068# 0.011912f
C456 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_21402_35420# 0.160931f
C457 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S 0.010488f
C458 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_17750_41880# 0.072448f
C459 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.437693f
C460 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.803935f
C461 a_22790_43112# SUNSAR_SAR8B_CV_0.EN 0.030411f
C462 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] 0.17256f
C463 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_4038# 0.068911f
C464 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.034738f
C465 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S 0.011542f
C466 SUNSAR_SAR8B_CV_0.XA20.CPO a_18882_27852# 0.067964f
C467 a_15210_37532# a_15210_37180# 0.010937f
C468 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S 0.028011f
C469 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.070318f
C470 SUNSAR_SAR8B_CV_0.EN a_10170_29612# 0.143959f
C471 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.12241f
C472 a_7650_35948# SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.072725f
C473 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA20.CNO 0.065836f
C474 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_3782_42408# 0.074559f
C475 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_42408# 0.100131f
C476 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B a_9990_2982# 0.011407f
C477 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S a_16542_3334# 0.023111f
C478 SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR 9.97874f
C479 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_11322_31196# 0.010411f
C480 ui_in[7] ui_in[6] 0.023797f
C481 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_13862_43288# 0.031221f
C482 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S 0.030221f
C483 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.649845f
C484 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S 0.030434f
C485 SUNSAR_SAR8B_CV_0.SARP a_13950_5446# 0.010143f
C486 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR 0.097407f
C487 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.SARN 0.038745f
C488 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.073351f
C489 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.166192f
C490 SUNSAR_SAR8B_CV_0.XA7.XA11.A a_20250_36300# 0.089492f
C491 a_23942_43640# VPWR 0.412992f
C492 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S uo_out[1] 0.01183f
C493 a_13842_29612# VPWR 0.397362f
C494 a_9990_4918# SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H 0.030771f
C495 a_16542_5270# a_16542_4918# 0.010937f
C496 a_2610_35068# a_2610_34716# 0.010937f
C497 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_20270_41000# 0.156079f
C498 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR 0.519052f
C499 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24678_4688# 0.0666f
C500 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 0.026917f
C501 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.011022f
C502 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA20.CNO 0.064502f
C503 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.339883f
C504 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.280191f
C505 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_18902_42408# 0.09112f
C506 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.055045f
C507 VPWR uo_out[4] 1.03021f
C508 m4_9630_44892# uio_oe[0] 0.025289f
C509 uo_out[7] uo_out[5] 1.57818f
C510 a_6302_43816# SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.071553f
C511 SUNSAR_SAR8B_CV_0.XA6.EN a_17730_27148# 0.071936f
C512 a_20270_41000# VPWR 0.388204f
C513 a_10190_41000# tt_um_TT06_SAR_done_0.DONE 0.067588f
C514 SUNSAR_SAR8B_CV_0.XA6.XA12.A a_18882_36828# 0.091063f
C515 SUNSAR_SAR8B_CV_0.XA7.CEIN a_20250_36828# 0.07472f
C516 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.010609f
C517 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.098057f
C518 a_22790_44344# clk 0.010581f
C519 TIE_L uo_out[0] 0.280844f
C520 a_7670_44168# uo_out[5] 0.04067f
C521 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.143554f
C522 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S 0.036491f
C523 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_20250_35420# 0.133834f
C524 SUNSAR_SAR8B_CV_0.XA7.XA9.B a_21402_35420# 0.017683f
C525 a_5130_27500# VPWR 0.382397f
C526 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S 0.028026f
C527 a_10190_41880# VPWR 0.395781f
C528 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.017094f
C529 SUNSAR_SAR8B_CV_0.XA0.XA2.A a_3762_30316# 0.129098f
C530 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.204048f
C531 SUNSAR_CAPT8B_CV_0.XA5.B tt_um_TT06_SAR_done_0.DONE 0.01988f
C532 SUNSAR_SAR8B_CV_0.XA20.CPO a_17730_27852# 0.072221f
C533 a_10170_32956# VPWR 0.436368f
C534 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 27.1615f
C535 a_12690_27852# a_12690_27500# 0.010937f
C536 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.062692f
C537 SUNSAR_SAR8B_CV_0.EN a_8802_29612# 0.143959f
C538 a_20250_28556# VPWR 0.406628f
C539 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S a_15390_3334# 0.036577f
C540 a_12582_3686# a_12582_3334# 0.010937f
C541 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.014291f
C542 a_11322_32076# SUNSAR_SAR8B_CV_0.XA3.CN1 0.06792f
C543 SUNSAR_SAR8B_CV_0.EN VPWR 41.914997f
C544 SUNSAR_CAPT8B_CV_0.XH13.XA6.A uo_out[1] 0.014139f
C545 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_43288# 0.069053f
C546 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_13862_43288# 0.080718f
C547 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S 0.055627f
C548 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.744161f
C549 SUNSAR_SAR8B_CV_0.XA20.CPO a_12690_28556# 0.014592f
C550 a_23942_40648# a_23942_40296# 0.010937f
C551 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_11142_2630# 0.011753f
C552 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S 0.050207f
C553 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.52234f
C554 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189272f
C555 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.166272f
C556 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C557 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN uo_out[1] 0.305131f
C558 a_11322_35068# SUNSAR_SAR8B_CV_0.XA4.EN 0.066018f
C559 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S 0.055045f
C560 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C561 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_2768# 0.049023f
C562 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VPWR 0.452478f
C563 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18126_4848# 0.024512f
C564 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.152045f
C565 SUNSAR_SAR8B_CV_0.XA6.CP0 a_18882_32956# 0.070763f
C566 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.738992f
C567 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_17750_42408# 0.111909f
C568 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S 0.089305f
C569 m4_8894_44892# uio_oe[0] 0.025289f
C570 VPWR uo_out[5] 1.02721f
C571 uo_out[7] uo_out[6] 2.38922f
C572 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S 0.076714f
C573 a_18902_41000# VPWR 0.388305f
C574 a_8822_41000# tt_um_TT06_SAR_done_0.DONE 0.066018f
C575 a_3782_41000# a_3782_40648# 0.010937f
C576 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.55251f
C577 a_10170_35420# VPWR 0.39968f
C578 SUNSAR_SAR8B_CV_0.XA6.XA12.A a_17730_36828# 0.10248f
C579 SUNSAR_SAR8B_CV_0.XA7.CEIN a_18882_36828# 0.015625f
C580 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.02121f
C581 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.111867f
C582 TIE_L uo_out[1] 0.50141f
C583 a_10190_44168# VPWR 0.340085f
C584 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR 2.45124f
C585 a_15210_27148# a_15210_26796# 0.010937f
C586 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_SAR8B_CV_0.D<5> 0.241356f
C587 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.014291f
C588 a_3762_27500# VPWR 0.382189f
C589 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.SARN 0.052813f
C590 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.331207f
C591 a_8822_41880# VPWR 0.395781f
C592 SUNSAR_SAR8B_CV_0.XA0.XA2.A a_2610_30316# 0.089492f
C593 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.276252f
C594 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.010345f
C595 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_28204# 0.016912f
C596 SUNSAR_SAR8B_CV_0.D<4> a_11342_41352# 0.079434f
C597 SUNSAR_CAPT8B_CV_0.XA5.B a_23942_41000# 0.091365f
C598 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S 0.050207f
C599 SUNSAR_SAR8B_CV_0.XA20.CPO a_16362_27852# 0.073806f
C600 a_10170_36300# VPWR 0.398846f
C601 a_13842_37532# a_13842_37180# 0.010937f
C602 a_8802_32956# VPWR 0.436368f
C603 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S 0.073313f
C604 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.138246f
C605 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_13862_42760# 0.031082f
C606 a_18882_28556# VPWR 0.406628f
C607 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.026794f
C608 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.CNO 0.159359f
C609 a_10170_32076# SUNSAR_SAR8B_CV_0.XA3.CN1 0.067588f
C610 a_23942_43112# VPWR 0.393308f
C611 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO 0.464697f
C612 uio_in[0] ui_in[7] 0.023797f
C613 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_12710_43288# 0.028213f
C614 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S 0.026885f
C615 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S 0.024386f
C616 a_5130_37180# VPWR 0.474051f
C617 SUNSAR_SAR8B_CV_0.XA20.CPO a_11322_28556# 0.014652f
C618 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S 0.064105f
C619 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_8802_27852# 0.028807f
C620 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR 4.24041f
C621 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.166192f
C622 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.021942f
C623 SUNSAR_SAR8B_CV_0.D<4> a_10170_33836# 0.011975f
C624 SUNSAR_CAPT8B_CV_0.XH13.XA7.C uo_out[1] 0.245678f
C625 a_15390_5270# a_15390_4918# 0.010937f
C626 a_10170_35068# SUNSAR_SAR8B_CV_0.XA4.EN 0.071277f
C627 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24678_2768# 0.024512f
C628 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18054_4848# 0.024512f
C629 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 0.026917f
C630 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.011022f
C631 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.028032f
C632 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA20.CPO 0.064038f
C633 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C634 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_16382_41880# 0.067588f
C635 m4_8158_44892# uio_oe[0] 0.025289f
C636 VPWR uo_out[6] 1.34623f
C637 SUNSAR_SAR8B_CV_0.XA5.EN a_16362_27148# 0.082474f
C638 a_5150_43816# SUNSAR_CAPT8B_CV_0.XC08.XA7.CN 0.071475f
C639 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S 0.055045f
C640 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S 0.050207f
C641 a_7670_41000# tt_um_TT06_SAR_done_0.DONE 0.070731f
C642 a_8802_35420# VPWR 0.39968f
C643 a_6282_28556# SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.066018f
C644 SUNSAR_SAR8B_CV_0.D<6> a_5130_34716# 0.070775f
C645 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA5.EN 0.439535f
C646 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.010771f
C647 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S 0.011641f
C648 a_6302_44168# uo_out[6] 0.044469f
C649 SUNSAR_CAPT8B_CV_0.XB07.QN TIE_L2 0.012775f
C650 a_8822_44168# VPWR 0.3405f
C651 TIE_L uo_out[2] 0.156661f
C652 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR 2.44986f
C653 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.DONE 0.034185f
C654 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S 0.021266f
C655 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_SAR8B_CV_0.D<5> 0.393076f
C656 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_6282_35068# 0.129098f
C657 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_10190_42408# 0.015723f
C658 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.020079f
C659 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> a_13842_33836# 0.103403f
C660 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.030618f
C661 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S 0.011494f
C662 SUNSAR_SAR8B_CV_0.D<4> a_10190_41352# 0.06659f
C663 SUNSAR_CAPT8B_CV_0.XA5.B a_22790_41000# 0.11811f
C664 SUNSAR_SAR8B_CV_0.XA20.CPO a_15210_27852# 0.066394f
C665 a_8802_36300# VPWR 0.399161f
C666 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.011847f
C667 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S 0.028011f
C668 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.030446f
C669 a_11322_27852# a_11322_27500# 0.010937f
C670 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S a_21402_27500# 0.036993f
C671 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.205884f
C672 SUNSAR_SAR8B_CV_0.D<1> a_18882_32076# 0.020342f
C673 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA20.CNO 0.058767f
C674 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.080525f
C675 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.626084f
C676 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_42760# 0.031591f
C677 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.TIE_L 6.83332f
C678 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.441867f
C679 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.026917f
C680 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 a_23922_31724# 0.023357f
C681 SUNSAR_SAR8B_CV_0.XA20.XA3.CO a_23922_30844# 0.077046f
C682 a_3762_37180# VPWR 0.473713f
C683 a_22790_40648# a_22790_40296# 0.010937f
C684 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.021955f
C685 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_16542_2982# 0.068023f
C686 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.078539f
C687 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.166272f
C688 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.SARN 0.034649f
C689 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S VPWR 0.106927f
C690 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.010347f
C691 a_10170_29612# VPWR 0.397362f
C692 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA9.Y 1.59176f
C693 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18126_2928# 0.0666f
C694 a_9990_4918# VPWR 0.468783f
C695 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_5648# 0.172147f
C696 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 0.012272f
C697 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA20.CNO 0.066024f
C698 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.154232f
C699 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.74103f
C700 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_16382_42408# 0.113479f
C701 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_15230_41880# 0.071088f
C702 a_23942_42760# a_23942_42408# 0.010937f
C703 m4_7422_44892# uio_oe[0] 0.02529f
C704 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.318734f
C705 VPWR uo_out[7] 1.27659f
C706 TIE_L SUNSAR_CAPT8B_CV_0.XA6.B 0.019831f
C707 SUNSAR_SAR8B_CV_0.XA5.EN a_15210_27148# 0.01235f
C708 a_6302_41000# tt_um_TT06_SAR_done_0.DONE 0.06916f
C709 a_2630_41000# a_2630_40648# 0.010937f
C710 a_5130_28556# SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.071498f
C711 SUNSAR_SAR8B_CV_0.XA6.CEIN a_18882_36828# 0.066018f
C712 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.303978f
C713 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.098057f
C714 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.182408f
C715 TIE_L uo_out[3] 0.185333f
C716 a_5150_44168# uo_out[6] 0.035338f
C717 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR 2.45309f
C718 a_13842_27148# a_13842_26796# 0.010937f
C719 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6519f
C720 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_16382_41880# 0.070877f
C721 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S 0.021211f
C722 SUNSAR_SAR8B_CV_0.XA1.XA9.B a_6282_35068# 0.011912f
C723 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_5130_35068# 0.089492f
C724 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_18882_35420# 0.133834f
C725 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B 0.254583f
C726 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.014291f
C727 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.CNO 0.108751f
C728 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 4.31242f
C729 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.035675f
C730 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.CKN 0.101993f
C731 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_28204# 0.017441f
C732 SUNSAR_SAR8B_CV_0.XA20.CPO a_13842_27852# 0.067964f
C733 a_12690_37532# a_12690_37180# 0.010937f
C734 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.106828f
C735 SUNSAR_SAR8B_CV_0.EN a_5130_29612# 0.143959f
C736 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S 0.044855f
C737 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.12241f
C738 a_6282_35948# SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.071154f
C739 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S 0.016737f
C740 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 a_22770_31724# 0.035229f
C741 a_8802_32076# SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.066018f
C742 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_7650_31196# 0.010411f
C743 SUNSAR_SAR8B_CV_0.XA20.XA3.CO a_22770_30844# 0.068231f
C744 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.324243f
C745 uio_in[1] uio_in[0] 0.023797f
C746 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.072852f
C747 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S 0.036094f
C748 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.011346f
C749 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_15390_2982# 0.078536f
C750 SUNSAR_SAR8B_CV_0.XA20.CK_CMP a_23922_35948# 0.067588f
C751 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.166192f
C752 SUNSAR_SAR8B_CV_0.XA6.XA11.A a_18882_36300# 0.091063f
C753 SUNSAR_CAPT8B_CV_0.XI14.XA7.C VPWR 2.97223f
C754 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S uo_out[2] 0.01183f
C755 a_8802_29612# VPWR 0.397362f
C756 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C757 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_23922_34892# 0.069155f
C758 a_8802_35068# SUNSAR_SAR8B_CV_0.XA3.EN 0.069707f
C759 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18054_2928# 0.105547f
C760 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.40569f
C761 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24678_5648# 0.0666f
C762 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S 0.010423f
C763 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.3401f
C764 SUNSAR_SAR8B_CV_0.XA5.CP0 a_16362_32956# 0.102695f
C765 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_15230_42408# 0.08955f
C766 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.B 0.016319f
C767 m4_6686_44892# uio_oe[0] 0.032443f
C768 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.093019f
C769 a_28727_41363# uio_oe[0] 0.027581f
C770 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.010751f
C771 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.018785f
C772 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_27148# 0.010025f
C773 a_15230_41000# VPWR 0.388204f
C774 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S 0.030434f
C775 a_5150_41000# tt_um_TT06_SAR_done_0.DONE 0.067588f
C776 SUNSAR_SAR8B_CV_0.XA5.XA12.A a_16362_36828# 0.104051f
C777 SUNSAR_SAR8B_CV_0.XA6.CEIN a_17730_36828# 0.070731f
C778 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.054448f
C779 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.13078f
C780 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.291229f
C781 TIE_L uo_out[4] 0.31941f
C782 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR 2.45309f
C783 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_17730_35420# 0.160931f
C784 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_16382_41880# 0.031087f
C785 a_20250_27852# VPWR 0.358413f
C786 a_5150_41880# VPWR 0.395781f
C787 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.SARP 0.054558f
C788 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.204048f
C789 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S 0.013533f
C790 SUNSAR_SAR8B_CV_0.XA20.CPO a_12690_27852# 0.072221f
C791 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.070269f
C792 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_21402_34716# 0.072552f
C793 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.097975f
C794 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6519f
C795 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S 0.030221f
C796 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.649845f
C797 a_10170_27852# a_10170_27500# 0.010937f
C798 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.432466f
C799 a_5130_32956# VPWR 0.436368f
C800 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S 0.073313f
C801 SUNSAR_SAR8B_CV_0.EN a_3762_29612# 0.143959f
C802 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.104691f
C803 a_5130_35948# SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.067588f
C804 a_15210_28556# VPWR 0.406628f
C805 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.175342f
C806 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.441867f
C807 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.026917f
C808 a_7650_32076# SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.06949f
C809 SUNSAR_CAPT8B_CV_0.XG12.XA6.A uo_out[2] 0.014222f
C810 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C811 SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR 1.63909f
C812 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.63636f
C813 SUNSAR_SAR8B_CV_0.XA20.CPO a_7650_28556# 0.014592f
C814 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S 0.030434f
C815 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N a_21402_29612# 0.031412f
C816 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.106002f
C817 a_21422_40648# a_21422_40296# 0.010937f
C818 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR 0.112858f
C819 SUNSAR_SAR8B_CV_0.XA20.CK_CMP a_22770_35948# 0.070536f
C820 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.206912f
C821 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.201839f
C822 SUNSAR_SAR8B_CV_0.XA6.XA11.A a_17730_36300# 0.13253f
C823 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S 0.016767f
C824 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN VPWR 1.77591f
C825 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S uo_out[2] 0.023976f
C826 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_22770_34892# 0.089422f
C827 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S 0.026506f
C828 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S 0.055045f
C829 a_7650_35068# SUNSAR_SAR8B_CV_0.XA3.EN 0.067588f
C830 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_3728# 0.049023f
C831 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18126_5808# 0.024512f
C832 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CN1 0.050135f
C833 SUNSAR_SAR8B_CV_0.XA5.CP0 a_15210_32956# 0.069193f
C834 a_22790_42760# a_22790_42408# 0.010937f
C835 TIE_L2 uio_oe[0] 0.014206f
C836 TIE_L1 uo_out[5] 0.275786f
C837 a_27575_41363# uio_oe[0] 0.01232f
C838 a_13862_41000# VPWR 0.388305f
C839 a_28727_41363# a_28727_41011# 0.010937f
C840 a_3782_41000# tt_um_TT06_SAR_done_0.DONE 0.066018f
C841 a_5130_35420# VPWR 0.39968f
C842 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.55251f
C843 SUNSAR_SAR8B_CV_0.XA5.XA12.A a_15210_36828# 0.089492f
C844 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.012048f
C845 TIE_L uo_out[5] 1.3092f
C846 a_3782_44168# uo_out[7] 0.040727f
C847 a_5150_44168# VPWR 0.340085f
C848 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR 2.45309f
C849 a_12690_27148# a_12690_26796# 0.010937f
C850 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_41880# 0.100592f
C851 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.145738f
C852 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C853 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.026917f
C854 a_18882_27852# VPWR 0.358599f
C855 a_3782_41880# VPWR 0.395781f
C856 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_4390# 0.156896f
C857 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.SARP 0.062266f
C858 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S 0.077008f
C859 SUNSAR_SAR8B_CV_0.XA20.CPO a_11322_27852# 0.073806f
C860 a_5130_36300# VPWR 0.398846f
C861 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S 0.050207f
C862 a_11322_37532# a_11322_37180# 0.010937f
C863 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S 0.055627f
C864 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.744161f
C865 a_3762_32956# VPWR 0.436368f
C866 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.06595f
C867 SUNSAR_SAR8B_CV_0.EN a_2610_29612# 0.076552f
C868 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.062692f
C869 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA20.CNO 0.056212f
C870 a_13842_28556# VPWR 0.406628f
C871 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S a_11142_3334# 0.036577f
C872 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.473914f
C873 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.070343f
C874 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S 0.012065f
C875 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_6282_31196# 0.010411f
C876 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C877 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S VPWR 0.097536f
C878 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S 0.050207f
C879 uio_in[2] uio_in[1] 0.023797f
C880 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S 0.026885f
C881 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_11342_43288# 0.028213f
C882 SUNSAR_SAR8B_CV_0.XA20.CPO a_6282_28556# 0.014652f
C883 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N a_3762_28908# 0.023475f
C884 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.073013f
C885 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S 0.030434f
C886 a_20250_37532# VPWR 0.454489f
C887 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.028567f
C888 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S 0.050207f
C889 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.078539f
C890 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR 0.112858f
C891 SUNSAR_SAR8B_CV_0.D<5> a_8802_33836# 0.011974f
C892 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.SARN 0.034649f
C893 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S VPWR 0.106927f
C894 SUNSAR_CAPT8B_CV_0.XG12.XA7.C uo_out[2] 0.246146f
C895 a_11142_5270# a_11142_4918# 0.010937f
C896 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_18902_41000# 0.15757f
C897 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S 0.055045f
C898 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24678_3728# 0.024512f
C899 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C900 a_16542_5270# VPWR 0.489055f
C901 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18054_5808# 0.024512f
C902 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S 0.010423f
C903 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.028032f
C904 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_13862_42408# 0.09112f
C905 TIE_L1 uo_out[6] 0.036047f
C906 a_3782_43816# SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.069905f
C907 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S 0.055045f
C908 SUNSAR_SAR8B_CV_0.XA20.CPO a_22770_29964# 0.01114f
C909 SUNSAR_SAR8B_CV_0.XA4.EN a_12690_27148# 0.071936f
C910 a_2630_41000# tt_um_TT06_SAR_done_0.DONE 0.070731f
C911 a_3762_35420# VPWR 0.39968f
C912 a_3762_28556# SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.069927f
C913 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA4.EN 0.50443f
C914 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.CP0 0.056326f
C915 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.352238f
C916 a_3782_44168# VPWR 0.3405f
C917 TIE_L uo_out[6] 0.204625f
C918 a_2630_44168# uo_out[7] 0.041756f
C919 SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR 2.45309f
C920 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_8822_42408# 0.015723f
C921 SUNSAR_SAR8B_CV_0.XA6.XA9.B a_17730_35420# 0.017683f
C922 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_3762_35068# 0.091063f
C923 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.DONE 0.076485f
C924 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S 0.028026f
C925 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.118161f
C926 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.011542f
C927 a_21402_31196# SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.066018f
C928 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.SARP 0.257526f
C929 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_4390# 0.156514f
C930 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.30776f
C931 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S 0.013533f
C932 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<1> 0.010193f
C933 SUNSAR_SAR8B_CV_0.D<5> a_8822_41352# 0.06816f
C934 SUNSAR_SAR8B_CV_0.XA20.CPO a_10170_27852# 0.066394f
C935 a_3762_36300# VPWR 0.399161f
C936 SUNSAR_SAR8B_CV_0.SARN a_13950_4038# 0.014345f
C937 a_8802_27852# a_8802_27500# 0.010937f
C938 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S 0.026885f
C939 SUNSAR_SAR8B_CV_0.D<7> a_3762_31196# 0.070763f
C940 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.205884f
C941 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 0.626356f
C942 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S a_9990_3334# 0.023111f
C943 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_2630# 0.067363f
C944 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.098257f
C945 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.021241f
C946 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S VPWR 0.097536f
C947 a_6282_32076# SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.06792f
C948 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CN1 0.466783f
C949 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C950 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.019092f
C951 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_SAR8B_CV_0.D<0> 0.010401f
C952 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S 0.055627f
C953 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.A 0.744161f
C954 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_11342_43288# 0.067482f
C955 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_10190_43288# 0.082288f
C956 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N a_2610_28908# 0.060353f
C957 a_18882_37532# VPWR 0.458364f
C958 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.075015f
C959 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.013868f
C960 a_20270_40648# a_20270_40296# 0.010937f
C961 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_11142_2982# 0.080106f
C962 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S 0.064105f
C963 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_5130_27852# 0.028807f
C964 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C965 SUNSAR_SAR8B_CV_0.XA5.XA11.A a_16362_36300# 0.13402f
C966 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.10065f
C967 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN uo_out[2] 0.305131f
C968 a_5130_29612# VPWR 0.397362f
C969 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_17750_41000# 0.114097f
C970 a_6282_35068# SUNSAR_SAR8B_CV_0.XA2.EN 0.066018f
C971 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA7.EN 0.291697f
C972 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18126_3888# 0.0666f
C973 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_6608# 0.172147f
C974 SUNSAR_SAR8B_CV_0.XA7.EN a_21402_30316# 0.06916f
C975 SUNSAR_SAR8B_CV_0.XA4.CP0 a_13842_32956# 0.070763f
C976 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_12710_42408# 0.111909f
C977 a_21422_42760# a_21422_42408# 0.010937f
C978 TIE_L1 uo_out[7] 0.206895f
C979 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S 0.076714f
C980 a_23942_41352# clk 0.067588f
C981 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.015869f
C982 a_27575_41363# a_27575_41011# 0.010937f
C983 a_2610_28556# SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.067588f
C984 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.CP0 0.033345f
C985 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.CP0 0.056173f
C986 SUNSAR_SAR8B_CV_0.XA5.CEIN a_16362_36828# 0.0733f
C987 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.EN 0.070866f
C988 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.054448f
C989 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.033093f
C990 SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR 2.45309f
C991 TIE_L uo_out[7] 0.471918f
C992 a_11322_27148# a_11322_26796# 0.010937f
C993 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.55251f
C994 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S 0.021211f
C995 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_2610_35068# 0.127528f
C996 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C997 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.026917f
C998 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.13041f
C999 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_28204# 0.016912f
C1000 a_20250_31196# SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.067827f
C1001 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR 0.118162f
C1002 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.128204f
C1003 SUNSAR_SAR8B_CV_0.D<5> a_7670_41352# 0.077864f
C1004 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.011542f
C1005 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.031163f
C1006 SUNSAR_SAR8B_CV_0.XA20.CPO a_8802_27852# 0.067964f
C1007 SUNSAR_SAR8B_CV_0.SARN a_12582_4038# 0.032882f
C1008 a_10170_37532# a_10170_37180# 0.010937f
C1009 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_17730_34716# 0.070402f
C1010 SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR 4.93712f
C1011 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 0.010379f
C1012 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.11099f
C1013 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.098494f
C1014 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.098737f
C1015 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.030127f
C1016 SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR 1.63909f
C1017 a_5130_32076# SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.067588f
C1018 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S 0.012065f
C1019 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C1020 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S 0.050207f
C1021 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_43288# 0.031221f
C1022 uio_in[3] uio_in[2] 0.023797f
C1023 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA6.A 0.649845f
C1024 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S 0.030221f
C1025 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.073013f
C1026 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.183415f
C1027 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.016812f
C1028 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_9990_2982# 0.066453f
C1029 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR 3.09702f
C1030 SUNSAR_SAR8B_CV_0.XA5.XA11.A a_15210_36300# 0.089492f
C1031 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN VPWR 1.7759f
C1032 a_9990_5270# a_9990_4918# 0.010937f
C1033 a_3762_29612# VPWR 0.397362f
C1034 a_5130_35068# SUNSAR_SAR8B_CV_0.XA2.EN 0.071277f
C1035 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18054_3888# 0.105547f
C1036 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24678_6608# 0.0666f
C1037 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.074772f
C1038 SUNSAR_SAR8B_CV_0.XA4.CP0 a_12690_32956# 0.101124f
C1039 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.093019f
C1040 TIE_L1 VPWR 0.114647f
C1041 TIE_L SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.045419f
C1042 a_2630_43816# SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.073123f
C1043 a_10190_41000# VPWR 0.388224f
C1044 a_22790_41352# clk 0.073203f
C1045 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S 0.050207f
C1046 SUNSAR_SAR8B_CV_0.XA3.EN a_11322_27148# 0.082474f
C1047 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR 0.106794f
C1048 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.098057f
C1049 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.CP0 0.056326f
C1050 SUNSAR_SAR8B_CV_0.XA4.XA12.A a_13842_36828# 0.091063f
C1051 SUNSAR_SAR8B_CV_0.XA5.CEIN a_15210_36828# 0.07472f
C1052 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.010609f
C1053 TIE_L VPWR 0.387688f
C1054 SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR 2.45309f
C1055 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XA5.B 0.03255f
C1056 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S 0.021266f
C1057 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_SAR8B_CV_0.D<6> 0.39306f
C1058 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.020208f
C1059 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.143554f
C1060 a_15210_27852# VPWR 0.358413f
C1061 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.118161f
C1062 SUNSAR_CAPT8B_CV_0.XA5.B VPWR 1.20915f
C1063 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.CKN 0.101993f
C1064 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S 0.076247f
C1065 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87498f
C1066 SUNSAR_SAR8B_CV_0.XA20.CPO a_7650_27852# 0.072221f
C1067 a_23922_36652# VPWR 0.449853f
C1068 SUNSAR_SAR8B_CV_0.XA20.CNO a_21402_27500# 0.067588f
C1069 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_16362_34716# 0.068905f
C1070 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S a_17730_27500# 0.036993f
C1071 a_7650_27852# a_7650_27500# 0.010937f
C1072 a_23922_33132# VPWR 0.415713f
C1073 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.55549f
C1074 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.432466f
C1075 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_11342_42760# 0.031591f
C1076 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA20.CNO 0.180455f
C1077 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.062692f
C1078 a_3762_35948# SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.066018f
C1079 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.066004f
C1080 SUNSAR_SAR8B_CV_0.D<2> a_15210_32076# 0.020342f
C1081 a_10170_28556# VPWR 0.406628f
C1082 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.093469f
C1083 a_13950_2630# ua[0] 0.020368f
C1084 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.098257f
C1085 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.021241f
C1086 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C1087 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CN1 0.466783f
C1088 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.01601f
C1089 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.233892f
C1090 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S 0.044855f
C1091 SUNSAR_SAR8B_CV_0.XA20.CPO a_2610_28556# 0.014592f
C1092 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S 0.030434f
C1093 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.021304f
C1094 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CEIN 0.07415f
C1095 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.01121f
C1096 a_18902_40648# a_18902_40296# 0.010937f
C1097 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_16542_3334# 0.066018f
C1098 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S 0.050207f
C1099 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.SARN 0.034649f
C1100 SUNSAR_CAPT8B_CV_0.XH13.XA7.C VPWR 2.97208f
C1101 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S uo_out[3] 0.024336f
C1102 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_SAR8B_CV_0.D<3> 0.018133f
C1103 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1104 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.093524f
C1105 a_9990_5270# VPWR 0.490626f
C1106 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_4688# 0.049023f
C1107 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18126_6768# 0.024512f
C1108 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.26609f
C1109 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CN1 0.050197f
C1110 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_11342_42408# 0.113479f
C1111 a_20270_42760# a_20270_42408# 0.010937f
C1112 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.318734f
C1113 a_8822_41000# VPWR 0.388305f
C1114 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.386305f
C1115 SUNSAR_SAR8B_CV_0.XA3.EN a_10170_27148# 0.01235f
C1116 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VPWR 0.658328f
C1117 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 54.2165f
C1118 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.222689f
C1119 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.02121f
C1120 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.CP0 0.056173f
C1121 SUNSAR_SAR8B_CV_0.XA4.XA12.A a_12690_36828# 0.10248f
C1122 SUNSAR_SAR8B_CV_0.XA5.CEIN a_13842_36828# 0.015625f
C1123 a_23942_44344# VPWR 0.342053f
C1124 a_10170_27148# a_10170_26796# 0.010937f
C1125 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_13862_41880# 0.099022f
C1126 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_SAR8B_CV_0.D<6> 0.241356f
C1127 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_16362_35420# 0.160931f
C1128 SUNSAR_SAR8B_CV_0.XA0.XA9.B a_2610_35068# 0.011912f
C1129 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 0.021241f
C1130 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.098257f
C1131 a_13842_27852# VPWR 0.358599f
C1132 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.SARN 0.048717f
C1133 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> a_3762_32956# 0.017384f
C1134 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.129613f
C1135 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_28204# 0.017441f
C1136 a_18882_31196# SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.066256f
C1137 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.363295f
C1138 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S 0.011494f
C1139 SUNSAR_SAR8B_CV_0.XA20.CPO a_6282_27852# 0.073806f
C1140 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S 0.050207f
C1141 SUNSAR_SAR8B_CV_0.XA20.CNO a_20250_27500# 0.066018f
C1142 a_8802_37532# a_8802_37180# 0.010937f
C1143 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.030459f
C1144 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.12241f
C1145 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_42760# 0.031082f
C1146 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S 0.073313f
C1147 a_2610_35948# SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.072725f
C1148 a_8802_28556# VPWR 0.406628f
C1149 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_3334# 0.120042f
C1150 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S 0.028396f
C1151 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C1152 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_2610_31196# 0.010411f
C1153 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA20.CPO 0.057359f
C1154 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S 0.050207f
C1155 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S 0.036094f
C1156 uio_in[4] uio_in[3] 0.023797f
C1157 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.073013f
C1158 SUNSAR_SAR8B_CV_0.XA20.CPO a_21402_28908# 0.08706f
C1159 a_15210_37532# VPWR 0.459576f
C1160 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.093457f
C1161 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_15390_3334# 0.072629f
C1162 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S 0.064105f
C1163 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_3762_27852# 0.028807f
C1164 a_20250_34716# VPWR 0.396749f
C1165 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.155604f
C1166 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S 0.028452f
C1167 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S uo_out[3] 0.01219f
C1168 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR 0.337652f
C1169 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S 0.089305f
C1170 a_3762_35068# SUNSAR_SAR8B_CV_0.XA1.EN 0.069707f
C1171 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR 0.808658f
C1172 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24678_4688# 0.024512f
C1173 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_18054_6768# 0.024512f
C1174 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA20.CNO 0.064528f
C1175 SUNSAR_SAR8B_CV_0.XA3.CP0 a_11322_32956# 0.102695f
C1176 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_10190_42408# 0.08955f
C1177 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S 0.010488f
C1178 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.142061f
C1179 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.018832f
C1180 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_27148# 0.010025f
C1181 a_23942_41352# a_23942_41000# 0.010937f
C1182 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.036144f
C1183 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA3.EN 0.435786f
C1184 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.CP0 0.056326f
C1185 a_20250_31196# VPWR 0.437f
C1186 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_41880# 0.031087f
C1187 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S 0.030434f
C1188 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S 0.036491f
C1189 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.301485f
C1190 SUNSAR_SAR8B_CV_0.XA5.XA9.B a_16362_35420# 0.017683f
C1191 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_15210_35420# 0.133834f
C1192 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.DONE 0.034185f
C1193 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.066203f
C1194 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.118226f
C1195 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S 0.011542f
C1196 a_17730_31196# SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.067588f
C1197 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S VPWR 0.106927f
C1198 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.031841f
C1199 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.151273f
C1200 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S 0.010193f
C1201 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 1.62434f
C1202 SUNSAR_SAR8B_CV_0.XA20.CPO a_5130_27852# 0.066394f
C1203 SUNSAR_SAR8B_CV_0.XA7.XA11.A VPWR 0.718455f
C1204 SUNSAR_SAR8B_CV_0.XA20.CNO a_18882_27500# 0.067588f
C1205 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.098006f
C1206 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S a_16362_27500# 0.036993f
C1207 a_6282_27852# a_6282_27500# 0.010937f
C1208 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR 2.68142f
C1209 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S 0.026885f
C1210 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.08649f
C1211 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S 0.027192f
C1212 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.205884f
C1213 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_2630# 0.068977f
C1214 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_3334# 0.113134f
C1215 a_13950_4038# a_13950_3686# 0.010937f
C1216 a_12582_2630# ua[1] 0.020558f
C1217 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.419738f
C1218 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.058243f
C1219 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C1220 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CN1 0.466783f
C1221 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA20.CPO 0.058001f
C1222 SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR 1.63909f
C1223 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_SAR8B_CV_0.D<1> 0.010401f
C1224 ua[1] ua[2] 0.01847f
C1225 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A 0.057364f
C1226 a_13842_37532# VPWR 0.458421f
C1227 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.178114f
C1228 a_17750_40648# a_17750_40296# 0.010937f
C1229 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.030806f
C1230 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.078539f
C1231 a_18882_34716# VPWR 0.399819f
C1232 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C1233 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S VPWR 0.106927f
C1234 a_13950_5446# a_13950_5094# 0.010937f
C1235 a_23922_29964# VPWR 0.429137f
C1236 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN uo_out[3] 0.309657f
C1237 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_16382_41000# 0.115667f
C1238 a_2610_35068# SUNSAR_SAR8B_CV_0.XA1.EN 0.067588f
C1239 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18126_4848# 0.0666f
C1240 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.473354f
C1241 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.076376f
C1242 SUNSAR_SAR8B_CV_0.XA6.EN a_17730_30316# 0.070731f
C1243 SUNSAR_SAR8B_CV_0.XA3.CP0 a_10170_32956# 0.069193f
C1244 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.152052f
C1245 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.023976f
C1246 a_18902_42760# a_18902_42408# 0.010937f
C1247 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S 0.076714f
C1248 a_23942_43992# SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.066018f
C1249 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S 0.030434f
C1250 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.010898f
C1251 a_21402_28908# a_21402_28556# 0.010937f
C1252 SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR 1.20972f
C1253 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.056173f
C1254 SUNSAR_SAR8B_CV_0.XA4.CEIN a_13842_36828# 0.066018f
C1255 a_18882_31196# VPWR 0.44007f
C1256 a_8802_27148# a_8802_26796# 0.010937f
C1257 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.55251f
C1258 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_12710_41880# 0.072448f
C1259 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.026506f
C1260 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 0.021241f
C1261 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.098257f
C1262 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 4.45258f
C1263 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.13041f
C1264 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3a.A 0.530644f
C1265 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S VPWR 0.106927f
C1266 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S 0.077008f
C1267 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<1> 0.434706f
C1268 SUNSAR_SAR8B_CV_0.D<6> a_6302_41352# 0.079434f
C1269 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S 0.011542f
C1270 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR 0.101562f
C1271 SUNSAR_SAR8B_CV_0.XA20.CPO a_3762_27852# 0.067964f
C1272 SUNSAR_SAR8B_CV_0.XA20.CNO a_17730_27500# 0.066018f
C1273 a_7650_37532# a_7650_37180# 0.010937f
C1274 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_12690_34716# 0.070402f
C1275 SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR 2.65387f
C1276 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.744161f
C1277 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S 0.055627f
C1278 SUNSAR_SAR8B_CV_0.XA20.XA12.Y a_23922_35948# 0.033888f
C1279 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.066546f
C1280 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.023828f
C1281 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.098737f
C1282 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.026794f
C1283 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.504801f
C1284 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA20.CPO 0.057859f
C1285 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.010266f
C1286 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S 0.050207f
C1287 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_8822_43288# 0.031221f
C1288 ua[1] ua[3] 0.01847f
C1289 uio_in[5] uio_in[4] 0.023797f
C1290 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S 0.024386f
C1291 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.073013f
C1292 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA7.CEIN 0.019713f
C1293 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.021942f
C1294 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.SARN 0.034649f
C1295 SUNSAR_SAR8B_CV_0.XA4.XA11.A a_13842_36300# 0.091063f
C1296 SUNSAR_SAR8B_CV_0.D<6> a_5130_33836# 0.011975f
C1297 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G a_16542_5270# 0.073828f
C1298 SUNSAR_CAPT8B_CV_0.XF11.XA7.C uo_out[3] 0.249907f
C1299 SUNSAR_CAPT8B_CV_0.XG12.XA7.C VPWR 2.9722f
C1300 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.206292f
C1301 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_15230_41000# 0.156079f
C1302 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1303 SUNSAR_CAPT8B_CV_0.XA6.B a_23942_41352# 0.025015f
C1304 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18054_4848# 0.105547f
C1305 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C1306 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.149144f
C1307 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.030854f
C1308 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145339f
C1309 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_8822_42408# 0.09112f
C1310 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S 0.055045f
C1311 a_22790_43992# SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.071093f
C1312 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S 0.062799f
C1313 a_5150_41000# VPWR 0.38821f
C1314 SUNSAR_SAR8B_CV_0.XA7.EN a_21402_27500# 0.082231f
C1315 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_27500# 0.044989f
C1316 SUNSAR_SAR8B_CV_0.XA2.EN a_7650_27148# 0.071936f
C1317 a_22790_41352# a_22790_41000# 0.010937f
C1318 SUNSAR_SAR8B_CV_0.XA7.XA9.B VPWR 0.924613f
C1319 a_21402_37180# a_21402_36828# 0.010937f
C1320 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.05849f
C1321 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.056326f
C1322 SUNSAR_SAR8B_CV_0.XA4.CEIN a_12690_36828# 0.070731f
C1323 SUNSAR_SAR8B_CV_0.XA3.XA12.A a_11322_36828# 0.104051f
C1324 TIE_L TIE_L1 0.257767f
C1325 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_5150_42408# 0.015723f
C1326 a_10170_27852# VPWR 0.358413f
C1327 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.SARN 0.048717f
C1328 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.118161f
C1329 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C1330 a_16362_31196# SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.066018f
C1331 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.316693f
C1332 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.204048f
C1333 SUNSAR_SAR8B_CV_0.D<6> a_5150_41352# 0.06659f
C1334 SUNSAR_SAR8B_CV_0.XA20.CNO a_16362_27500# 0.067588f
C1335 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR 0.119314f
C1336 SUNSAR_SAR8B_CV_0.XB2.TIE_L ua[0] 1.52001f
C1337 SUNSAR_SAR8B_CV_0.XA20.CPO a_2610_27852# 0.072221f
C1338 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_11322_34716# 0.068905f
C1339 a_5130_27852# a_5130_27500# 0.010937f
C1340 SUNSAR_SAR8B_CV_0.SARP a_12582_2630# 0.023697f
C1341 SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR 2.65386f
C1342 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S 0.030221f
C1343 SUNSAR_SAR8B_CV_0.D<3> a_13842_32076# 0.020342f
C1344 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S 0.073313f
C1345 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.649845f
C1346 a_5130_28556# VPWR 0.406628f
C1347 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_2982# 0.158066f
C1348 a_12582_4038# a_12582_3686# 0.010937f
C1349 a_15390_4038# SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.071276f
C1350 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.SARN 0.591428f
C1351 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.419738f
C1352 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.058243f
C1353 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_23922_31724# 0.096918f
C1354 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CN1 0.466783f
C1355 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_43288# 0.069053f
C1356 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_8822_43288# 0.080718f
C1357 ua[1] ua[4] 0.01847f
C1358 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 0.63636f
C1359 tt_um_TT06_SAR_done_0.x3.MP1.G uio_out[0] 0.165429f
C1360 SUNSAR_SAR8B_CV_0.XA20.CPO a_17730_28908# 0.085247f
C1361 tt_um_TT06_SAR_done_0.DONE a_28727_39955# 0.067434f
C1362 a_16382_40648# a_16382_40296# 0.010937f
C1363 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_11142_3334# 0.071059f
C1364 SUNSAR_SAR8B_CV_0.XA4.XA11.A a_12690_36300# 0.13253f
C1365 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.028831f
C1366 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G a_15390_5270# 0.066018f
C1367 a_12582_5446# a_12582_5094# 0.010937f
C1368 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.010347f
C1369 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN VPWR 1.7759f
C1370 SUNSAR_CAPT8B_CV_0.XA6.B a_22790_41352# 0.036058f
C1371 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S 0.055045f
C1372 a_16542_5622# VPWR 0.472384f
C1373 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_5648# 0.049023f
C1374 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2502_2768# 0.0666f
C1375 a_22770_33132# SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.023111f
C1376 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA20.CNO 0.056065f
C1377 SUNSAR_SAR8B_CV_0.XA5.EN a_16362_30316# 0.06916f
C1378 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.022299f
C1379 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_8802_32956# 0.070763f
C1380 a_17750_42760# a_17750_42408# 0.010937f
C1381 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_7670_42408# 0.111909f
C1382 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.318734f
C1383 TIE_L SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.045419f
C1384 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S 0.050207f
C1385 a_3782_41000# VPWR 0.388305f
C1386 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S 0.050207f
C1387 a_20250_28908# a_20250_28556# 0.010937f
C1388 SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR 1.22023f
C1389 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 6.86675f
C1390 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.182595f
C1391 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.058943f
C1392 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.056173f
C1393 SUNSAR_SAR8B_CV_0.XA3.XA12.A a_10170_36828# 0.089492f
C1394 a_7650_27148# a_7650_26796# 0.010937f
C1395 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C1396 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_13842_35420# 0.133834f
C1397 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.054658f
C1398 SUNSAR_SAR8B_CV_0.EN a_20250_28908# 0.072887f
C1399 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.058243f
C1400 a_8802_27852# VPWR 0.358599f
C1401 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C1402 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.21623f
C1403 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.129613f
C1404 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.15005f
C1405 a_15210_31196# SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.067827f
C1406 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.025253f
C1407 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.126806f
C1408 SUNSAR_SAR8B_CV_0.XA20.CNO a_15210_27500# 0.066018f
C1409 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S 0.050207f
C1410 SUNSAR_SAR8B_CV_0.XA6.XA11.A VPWR 0.725614f
C1411 SUNSAR_SAR8B_CV_0.XB2.TIE_L ua[1] 0.845623f
C1412 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S 0.024478f
C1413 a_6282_37532# a_6282_37180# 0.010937f
C1414 SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR 2.65387f
C1415 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.062692f
C1416 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S 0.03516f
C1417 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_8822_42760# 0.031082f
C1418 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S 0.044855f
C1419 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.199522f
C1420 a_3762_28556# VPWR 0.406628f
C1421 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_22770_31724# 0.067834f
C1422 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_21402_32076# 0.089573f
C1423 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.SARP 0.524159f
C1424 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S 0.050207f
C1425 uio_in[6] uio_in[5] 0.023797f
C1426 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_7670_43288# 0.028213f
C1427 a_28727_40659# uio_out[0] 0.021625f
C1428 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.073013f
C1429 SUNSAR_SAR8B_CV_0.XA20.CPO a_16362_28908# 0.086948f
C1430 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N a_17730_29612# 0.031412f
C1431 a_10170_37532# VPWR 0.459696f
C1432 tt_um_TT06_SAR_done_0.DONE a_27575_39955# 0.069463f
C1433 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.179089f
C1434 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW a_9990_3334# 0.067588f
C1435 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S 0.050207f
C1436 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.078539f
C1437 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S a_20250_28204# 0.04865f
C1438 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_21402_28204# 0.067588f
C1439 a_15210_34716# VPWR 0.399819f
C1440 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S 0.028448f
C1441 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR 0.108436f
C1442 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S uo_out[4] 0.01183f
C1443 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S VPWR 0.106927f
C1444 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S 0.026506f
C1445 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S 0.089305f
C1446 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24678_5648# 0.024512f
C1447 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C1448 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_2768# 0.172147f
C1449 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> a_7650_32956# 0.101124f
C1450 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN 0.093019f
C1451 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43816# 0.129239f
C1452 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_27500# 0.054233f
C1453 SUNSAR_SAR8B_CV_0.XA1.EN a_6282_27148# 0.082474f
C1454 a_21422_41352# a_21422_41000# 0.010937f
C1455 a_20250_37180# a_20250_36828# 0.010937f
C1456 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA2.EN 0.493441f
C1457 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.061263f
C1458 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_21402_33836# 0.07476f
C1459 a_15210_31196# VPWR 0.44007f
C1460 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.301485f
C1461 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.DONE 0.076485f
C1462 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_12690_35420# 0.160931f
C1463 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S 0.036491f
C1464 SUNSAR_SAR8B_CV_0.EN a_18882_28908# 0.074323f
C1465 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.40619f
C1466 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.118226f
C1467 a_22790_44344# TIE_L 0.048319f
C1468 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S 0.076247f
C1469 SUNSAR_SAR8B_CV_0.XA20.XA3.CO a_23922_29964# 0.151031f
C1470 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S VPWR 0.106927f
C1471 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S 0.011494f
C1472 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<2> 2.9798f
C1473 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<1> 0.08537f
C1474 SUNSAR_SAR8B_CV_0.SARN a_12582_4390# 0.043858f
C1475 SUNSAR_SAR8B_CV_0.XA20.CNO a_13842_27500# 0.067588f
C1476 SUNSAR_SAR8B_CV_0.XA5.XA11.A VPWR 0.722887f
C1477 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.033333f
C1478 a_3762_27852# a_3762_27500# 0.010937f
C1479 SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR 2.65386f
C1480 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.205884f
C1481 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C1482 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.21461f
C1483 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_42760# 0.031591f
C1484 a_13950_2982# ua[0] 0.062855f
C1485 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.031784f
C1486 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.046398f
C1487 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_20250_32076# 0.066439f
C1488 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CN1 0.466783f
C1489 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_SAR8B_CV_0.D<2> 0.010401f
C1490 a_8802_37532# VPWR 0.45854f
C1491 a_27575_40659# uio_out[0] 0.046111f
C1492 tt_um_TT06_SAR_done_0.DONE a_28727_40307# 0.065834f
C1493 a_15230_40648# a_15230_40296# 0.010937f
C1494 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S 0.064105f
C1495 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_20250_28204# 0.096735f
C1496 a_13842_34716# VPWR 0.399819f
C1497 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.07478f
C1498 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S 0.016769f
C1499 SUNSAR_SAR8B_CV_0.XA3.XA11.A a_11322_36300# 0.13402f
C1500 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.SARN 0.034649f
C1501 a_16542_5622# a_16542_5270# 0.010937f
C1502 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N VPWR 0.279205f
C1503 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S uo_out[4] 0.023976f
C1504 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_SAR8B_CV_0.D<4> 0.018133f
C1505 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.093524f
C1506 a_16542_5974# VPWR 0.449888f
C1507 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18126_5808# 0.0666f
C1508 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_2928# 0.024512f
C1509 a_16382_42760# a_16382_42408# 0.010937f
C1510 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_6302_42408# 0.113479f
C1511 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.023976f
C1512 TIE_L2 uo_out[7] 0.099101f
C1513 SUNSAR_CAPT8B_CV_0.XI14.QN a_20270_43816# 0.089492f
C1514 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S 0.050207f
C1515 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.010898f
C1516 a_28727_41363# VPWR 0.440399f
C1517 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.375196f
C1518 SUNSAR_SAR8B_CV_0.XA1.EN a_5130_27148# 0.01235f
C1519 SUNSAR_SAR8B_CV_0.XA20.CNO a_21402_29612# 0.094795f
C1520 a_18882_28908# a_18882_28556# 0.010937f
C1521 SUNSAR_SAR8B_CV_0.XA6.XA9.B VPWR 0.930839f
C1522 SUNSAR_SAR8B_CV_0.XA3.CEIN a_11322_36828# 0.0733f
C1523 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.EN 0.064769f
C1524 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.324105f
C1525 a_13842_31196# VPWR 0.44007f
C1526 a_6282_27148# a_6282_26796# 0.010937f
C1527 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.2165f
C1528 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.026506f
C1529 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_SAR8B_CV_0.D<7> 0.241356f
C1530 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_11342_41880# 0.070877f
C1531 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.058243f
C1532 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C1533 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.13041f
C1534 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.72697f
C1535 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP 0.544952f
C1536 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.363295f
C1537 a_13842_31196# SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.066256f
C1538 SUNSAR_SAR8B_CV_0.XA20.XA3.CO a_22770_29964# 0.134249f
C1539 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S VPWR 0.106927f
C1540 SUNSAR_SAR8B_CV_0.XA20.CNO a_12690_27500# 0.066018f
C1541 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR 0.101979f
C1542 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.029317f
C1543 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_7650_34716# 0.070402f
C1544 a_5130_37532# a_5130_37180# 0.010937f
C1545 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR 2.75252f
C1546 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_20250_35948# 0.068853f
C1547 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S 0.028751f
C1548 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.215582f
C1549 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.107674f
C1550 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S 0.012065f
C1551 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S 0.050207f
C1552 uio_in[7] uio_in[6] 0.023797f
C1553 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.073013f
C1554 tt_um_TT06_SAR_done_0.x3.MP1.G ui_in[0] 0.02266f
C1555 tt_um_TT06_SAR_done_0.x4.MP0.G uio_out[0] 0.030222f
C1556 tt_um_TT06_SAR_done_0.DONE a_27575_40307# 0.071434f
C1557 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.027044f
C1558 a_28727_41011# a_28727_40659# 0.010937f
C1559 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.027995f
C1560 SUNSAR_SAR8B_CV_0.XA3.XA11.A a_10170_36300# 0.089492f
C1561 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN VPWR 1.7759f
C1562 SUNSAR_CAPT8B_CV_0.XE10.XA7.C uo_out[4] 0.246063f
C1563 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18054_5808# 0.105547f
C1564 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9054_2928# 0.024512f
C1565 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C1566 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_5150_42408# 0.08955f
C1567 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S 0.010488f
C1568 TIE_L2 VPWR 0.09991f
C1569 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S 0.055045f
C1570 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S 0.050207f
C1571 SUNSAR_SAR8B_CV_0.XA6.EN a_17730_27500# 0.085451f
C1572 SUNSAR_SAR8B_CV_0.XA20.CNO a_20250_29612# 0.011704f
C1573 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_27148# 0.010025f
C1574 a_20270_41352# a_20270_41000# 0.010937f
C1575 SUNSAR_SAR8B_CV_0.XA2.XA12.A a_8802_36828# 0.091063f
C1576 SUNSAR_SAR8B_CV_0.XA3.CEIN a_10170_36828# 0.07472f
C1577 a_18882_37180# a_18882_36828# 0.010937f
C1578 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.138f
C1579 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S 0.030434f
C1580 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_3782_42408# 0.015723f
C1581 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C1582 SUNSAR_SAR8B_CV_0.XA4.XA9.B a_12690_35420# 0.017683f
C1583 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S 0.021266f
C1584 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_SAR8B_CV_0.D<7> 0.393125f
C1585 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_11342_41880# 0.031087f
C1586 a_5130_27852# VPWR 0.358413f
C1587 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.118161f
C1588 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> a_8802_33836# 0.103403f
C1589 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 3.79361f
C1590 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.031841f
C1591 a_12690_31196# SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.067588f
C1592 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.057478f
C1593 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.204048f
C1594 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S 0.013533f
C1595 SUNSAR_SAR8B_CV_0.D<7> a_3782_41352# 0.06816f
C1596 SUNSAR_SAR8B_CV_0.XA20.CNO a_11322_27500# 0.067588f
C1597 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR 0.119314f
C1598 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.024478f
C1599 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_6282_34716# 0.068905f
C1600 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.082644f
C1601 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S a_23922_27148# 0.023111f
C1602 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S a_12690_27500# 0.036993f
C1603 a_2610_27852# a_2610_27500# 0.010937f
C1604 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR 2.75088f
C1605 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.062692f
C1606 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.178111f
C1607 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S 0.044234f
C1608 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_2982# 0.158066f
C1609 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.379175p
C1610 a_20250_28908# VPWR 0.395394f
C1611 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.175174f
C1612 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.046398f
C1613 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.031784f
C1614 a_12582_2982# ua[1] 0.062686f
C1615 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_18882_32076# 0.06801f
C1616 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.535113f
C1617 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S 0.050207f
C1618 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.060807f
C1619 tt_um_TT06_SAR_done_0.x4.MP0.G uio_oe[0] 0.073251f
C1620 SUNSAR_SAR8B_CV_0.XA20.CPO a_12690_28908# 0.085247f
C1621 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.178114f
C1622 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA6.CEIN 0.05126f
C1623 tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G 0.186749f
C1624 a_13862_40648# a_13862_40296# 0.010937f
C1625 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.064851f
C1626 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S 0.050207f
C1627 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S a_18882_28204# 0.04865f
C1628 SUNSAR_CAPT8B_CV_0.XF11.XA7.C VPWR 2.97211f
C1629 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN uo_out[4] 0.305131f
C1630 a_15390_5622# a_15390_5270# 0.010937f
C1631 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR 0.104609f
C1632 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1633 SUNSAR_SAR8B_CV_0.XA7.XA9.B a_21402_34716# 0.047651f
C1634 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S 0.055045f
C1635 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR 0.808658f
C1636 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_6608# 0.049023f
C1637 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2502_3728# 0.0666f
C1638 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_5130_32956# 0.069193f
C1639 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CN1 0.050135f
C1640 SUNSAR_SAR8B_CV_0.XA4.EN a_12690_30316# 0.070731f
C1641 a_15230_42760# a_15230_42408# 0.010937f
C1642 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.015882f
C1643 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S 0.076714f
C1644 SUNSAR_CAPT8B_CV_0.XH13.QN a_18902_43816# 0.091063f
C1645 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S 0.050207f
C1646 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S 0.050207f
C1647 a_23942_41352# VPWR 0.376408f
C1648 SUNSAR_SAR8B_CV_0.XA20.CNO a_18882_29612# 0.011248f
C1649 a_17730_28908# a_17730_28556# 0.010937f
C1650 SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR 1.2202f
C1651 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1615f
C1652 SUNSAR_SAR8B_CV_0.XA2.XA12.A a_7650_36828# 0.10248f
C1653 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.158152f
C1654 SUNSAR_SAR8B_CV_0.XA3.CEIN a_8802_36828# 0.015625f
C1655 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_17730_33836# 0.073189f
C1656 a_5130_27148# a_5130_26796# 0.010937f
C1657 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S 0.010335f
C1658 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S 0.021211f
C1659 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_41880# 0.100592f
C1660 SUNSAR_SAR8B_CV_0.EN a_15210_28908# 0.072753f
C1661 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.046398f
C1662 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.031784f
C1663 a_3762_27852# VPWR 0.358599f
C1664 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.129613f
C1665 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S 0.077008f
C1666 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_4742# 0.157637f
C1667 SUNSAR_SAR8B_CV_0.D<7> a_2630_41352# 0.077864f
C1668 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<2> 0.233744f
C1669 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C1670 SUNSAR_SAR8B_CV_0.XA20.CNO a_10170_27500# 0.066018f
C1671 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S 0.050207f
C1672 SUNSAR_SAR8B_CV_0.XA4.XA11.A VPWR 0.725614f
C1673 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.024423f
C1674 a_3762_37532# a_3762_37180# 0.010937f
C1675 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR 2.75432f
C1676 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S 0.044855f
C1677 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S 0.073313f
C1678 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_18882_35948# 0.070424f
C1679 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.50324f
C1680 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.038188f
C1681 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.26479f
C1682 a_11142_4038# SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.069705f
C1683 a_18882_28908# VPWR 0.395394f
C1684 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.070949f
C1685 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_17730_32076# 0.088002f
C1686 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.SARP 0.013998f
C1687 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S 0.012065f
C1688 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.026146f
C1689 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S 0.050207f
C1690 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_6302_43288# 0.028213f
C1691 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S 0.024386f
C1692 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.072852f
C1693 SUNSAR_SAR8B_CV_0.XA20.CPO a_11322_28908# 0.086948f
C1694 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S 0.030434f
C1695 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N a_16362_29612# 0.031412f
C1696 a_5130_37532# VPWR 0.459635f
C1697 a_27575_41011# a_27575_40659# 0.010937f
C1698 a_28727_41011# tt_um_TT06_SAR_done_0.x4.MP0.G 0.065834f
C1699 a_10170_34716# VPWR 0.399819f
C1700 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_18882_28204# 0.098305f
C1701 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S 0.064105f
C1702 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C1703 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.010335f
C1704 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.40916f
C1705 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.072622f
C1706 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_13862_41000# 0.15757f
C1707 SUNSAR_SAR8B_CV_0.XA7.XA9.B a_20250_34716# 0.023982f
C1708 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24678_6608# 0.024512f
C1709 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_3728# 0.172147f
C1710 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.303428f
C1711 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_3782_42408# 0.09112f
C1712 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.093019f
C1713 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43816# 0.127669f
C1714 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_23922_27148# 0.067588f
C1715 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S 0.050207f
C1716 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.383512f
C1717 SUNSAR_SAR8B_CV_0.XA5.EN a_16362_27500# 0.082231f
C1718 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_27500# 0.044989f
C1719 SUNSAR_SAR8B_CV_0.XA20.CNO a_17730_29612# 0.090551f
C1720 a_18902_41352# a_18902_41000# 0.010937f
C1721 SUNSAR_SAR8B_CV_0.XA5.XA9.B VPWR 0.93081f
C1722 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA1.EN 0.113413f
C1723 a_17730_37180# a_17730_36828# 0.010937f
C1724 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_16362_33836# 0.07476f
C1725 a_10170_31196# VPWR 0.44007f
C1726 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S 0.023798f
C1727 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.DONE 0.034185f
C1728 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.017528f
C1729 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.301485f
C1730 SUNSAR_SAR8B_CV_0.EN a_13842_28908# 0.074323f
C1731 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.118226f
C1732 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S 0.013533f
C1733 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_23922_28556# 0.067713f
C1734 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.316693f
C1735 a_11322_31196# SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.066018f
C1736 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S VPWR 0.106927f
C1737 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_4742# 0.157255f
C1738 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<3> 0.010193f
C1739 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.42282f
C1740 SUNSAR_SAR8B_CV_0.XA20.CNO a_8802_27500# 0.067588f
C1741 SUNSAR_SAR8B_CV_0.XA3.XA11.A VPWR 0.722887f
C1742 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S a_11322_27500# 0.036993f
C1743 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S a_21402_27852# 0.056787f
C1744 SUNSAR_SAR8B_CV_0.SARP a_12582_2982# 0.037284f
C1745 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S 0.030221f
C1746 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA6.A 0.649845f
C1747 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.205884f
C1748 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C1749 SUNSAR_SAR8B_CV_0.D<4> a_10170_32076# 0.020342f
C1750 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.669708f
C1751 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_3334# 0.114704f
C1752 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3334# 0.163985f
C1753 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.CP0 0.010925f
C1754 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.449584f
C1755 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 0.014291f
C1756 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.55953f
C1757 SUNSAR_SAR8B_CV_0.XA7.EN a_21402_29612# 0.073155f
C1758 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.015993f
C1759 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_SAR8B_CV_0.D<3> 0.010401f
C1760 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S 0.050207f
C1761 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_5150_43288# 0.082288f
C1762 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_6302_43288# 0.067482f
C1763 a_3762_37532# VPWR 0.458479f
C1764 a_12710_40648# a_12710_40296# 0.010937f
C1765 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CEIN 0.075193f
C1766 a_27575_41011# tt_um_TT06_SAR_done_0.x4.MP0.G 0.097391f
C1767 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.059546f
C1768 a_8802_34716# VPWR 0.399819f
C1769 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_17730_28204# 0.066018f
C1770 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.078539f
C1771 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S uo_out[5] 0.023976f
C1772 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S VPWR 0.106927f
C1773 a_16542_5622# SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G 0.096614f
C1774 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR 0.051878f
C1775 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_12710_41000# 0.114097f
C1776 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_21422_41352# 0.078431f
C1777 a_9990_5622# VPWR 0.470814f
C1778 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18126_6768# 0.0666f
C1779 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_3888# 0.024512f
C1780 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_3762_32956# 0.070763f
C1781 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.244517f
C1782 SUNSAR_SAR8B_CV_0.XA3.EN a_11322_30316# 0.06916f
C1783 a_13862_42760# a_13862_42408# 0.010937f
C1784 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_2630_42408# 0.111909f
C1785 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_22770_27148# 0.06916f
C1786 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.318734f
C1787 SUNSAR_SAR8B_CV_0.XA20.CNO a_16362_29612# 0.095246f
C1788 SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR 1.22023f
C1789 a_16362_28908# a_16362_28556# 0.010937f
C1790 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.220689f
C1791 SUNSAR_SAR8B_CV_0.XA2.CEIN a_8802_36828# 0.066018f
C1792 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.DONE 0.054848f
C1793 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.86675f
C1794 a_8802_31196# VPWR 0.44007f
C1795 a_3762_27148# a_3762_26796# 0.010937f
C1796 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_11322_35420# 0.160931f
C1797 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.527529f
C1798 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.031784f
C1799 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.046398f
C1800 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VPWR 0.045952f
C1801 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.394834f
C1802 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.SARN 0.048683f
C1803 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.13041f
C1804 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_22770_28556# 0.140127f
C1805 a_10170_31196# SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.067827f
C1806 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S VPWR 0.106927f
C1807 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.126806f
C1808 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.01291f
C1809 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.CPO 7.93512f
C1810 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.011542f
C1811 SUNSAR_SAR8B_CV_0.XA20.CNO a_7650_27500# 0.066018f
C1812 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR 0.101979f
C1813 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_2610_34716# 0.070402f
C1814 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.029312f
C1815 a_2610_37532# a_2610_37180# 0.010937f
C1816 a_20250_33836# VPWR 0.407174f
C1817 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.A 0.744161f
C1818 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.230084f
C1819 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S 0.03516f
C1820 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_3334# 0.118471f
C1821 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_16362_32076# 0.089573f
C1822 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.0264f
C1823 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S 0.050207f
C1824 clk ena 0.023797f
C1825 uio_out[2] uio_out[1] 0.023797f
C1826 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA6.A 0.040072f
C1827 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_43288# 0.031221f
C1828 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S 0.036094f
C1829 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.179089f
C1830 SUNSAR_SAR8B_CV_0.XA2.XA11.A a_8802_36300# 0.091063f
C1831 SUNSAR_CAPT8B_CV_0.XE10.XA7.C VPWR 2.97224f
C1832 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S uo_out[5] 0.01183f
C1833 a_15390_5622# SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G 0.067588f
C1834 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR 0.042834f
C1835 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_20270_41352# 0.077076f
C1836 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_21422_41352# 0.060327f
C1837 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1838 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_18054_6768# 0.105547f
C1839 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C1840 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9054_3888# 0.024512f
C1841 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> a_2610_32956# 0.101124f
C1842 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA20.CNO 0.05498f
C1843 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S 0.010488f
C1844 SUNSAR_CAPT8B_CV_0.XG12.QN a_16382_43816# 0.129239f
C1845 a_20270_41352# VPWR 0.394053f
C1846 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S 0.062799f
C1847 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_27500# 0.054233f
C1848 SUNSAR_SAR8B_CV_0.XA20.CNO a_15210_29612# 0.011704f
C1849 a_17750_41352# a_17750_41000# 0.010937f
C1850 SUNSAR_SAR8B_CV_0.XA1.XA12.A a_6282_36828# 0.104051f
C1851 SUNSAR_SAR8B_CV_0.XA2.CEIN a_7650_36828# 0.070731f
C1852 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA7.CEIN 0.033943f
C1853 a_16362_37180# a_16362_36828# 0.010937f
C1854 SUNSAR_SAR8B_CV_0.XA3.XA9.B a_11322_35420# 0.017683f
C1855 SUNSAR_SAR8B_CV_0.XA3.XA9.A a_10170_35420# 0.133834f
C1856 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.107823f
C1857 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S VPWR 0.065445f
C1858 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.118161f
C1859 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S 0.076247f
C1860 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<1> 0.081799f
C1861 a_23942_41880# SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.06668f
C1862 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.D<3> 3.07227f
C1863 SUNSAR_SAR8B_CV_0.XA20.CNO a_6282_27500# 0.067588f
C1864 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR 0.119314f
C1865 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.024478f
C1866 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.087347f
C1867 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_21402_27148# 0.023111f
C1868 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S a_20250_27852# 0.04865f
C1869 SUNSAR_SAR8B_CV_0.SARN ua[0] 1.03115f
C1870 a_18882_33836# VPWR 0.409601f
C1871 a_23922_36300# a_23922_35948# 0.010937f
C1872 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_16362_35948# 0.134161f
C1873 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_6302_42760# 0.031591f
C1874 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.038188f
C1875 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A a_16542_4038# 0.01736f
C1876 a_15210_28908# VPWR 0.395394f
C1877 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_23922_34540# 0.067821f
C1878 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.089055f
C1879 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.02157f
C1880 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.449584f
C1881 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B 0.014291f
C1882 a_16542_2630# VPWR 0.448756f
C1883 a_13950_3334# ua[0] 0.060151f
C1884 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_15210_32076# 0.066439f
C1885 clk rst_n 0.024358f
C1886 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S 0.050207f
C1887 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.63636f
C1888 SUNSAR_SAR8B_CV_0.XA20.CPO a_7650_28908# 0.085247f
C1889 a_28727_39955# VPWR 0.355584f
C1890 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.030806f
C1891 a_11342_40648# a_11342_40296# 0.010937f
C1892 tt_um_TT06_SAR_done_0.DONE a_23942_40296# 0.025759f
C1893 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.010675f
C1894 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.073269f
C1895 SUNSAR_SAR8B_CV_0.XA2.XA11.A a_7650_36300# 0.13253f
C1896 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN VPWR 1.7759f
C1897 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN uo_out[5] 0.30523f
C1898 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G a_11142_5270# 0.067588f
C1899 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N VPWR 0.271482f
C1900 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_41352# 0.058557f
C1901 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_SAR8B_CV_0.D<5> 0.018133f
C1902 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S 0.055045f
C1903 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S 0.026506f
C1904 a_9990_5974# VPWR 0.451043f
C1905 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2502_4688# 0.0666f
C1906 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3a.A 0.205975f
C1907 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.18462f
C1908 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.036749f
C1909 a_12710_42760# a_12710_42408# 0.010937f
C1910 a_23942_42760# SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.066018f
C1911 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.023976f
C1912 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.015882f
C1913 SUNSAR_CAPT8B_CV_0.XG12.QN a_15230_43816# 0.089492f
C1914 SUNSAR_CAPT8B_CV_0.XA7.MP0.G SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.060853f
C1915 a_18902_41352# VPWR 0.394053f
C1916 SUNSAR_SAR8B_CV_0.XA20.CNO a_13842_29612# 0.011248f
C1917 SUNSAR_SAR8B_CV_0.XA4.XA9.B VPWR 0.930839f
C1918 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6519f
C1919 a_15210_28908# a_15210_28556# 0.010937f
C1920 SUNSAR_SAR8B_CV_0.XA1.XA12.A a_5130_36828# 0.089492f
C1921 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.377598f
C1922 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_12690_33836# 0.073189f
C1923 a_2610_27148# a_2610_26796# 0.010937f
C1924 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_8822_41880# 0.099022f
C1925 SUNSAR_SAR8B_CV_0.EN a_10170_28908# 0.072753f
C1926 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S VPWR 0.066675f
C1927 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.014291f
C1928 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.449584f
C1929 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S 0.028026f
C1930 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 4.68155f
C1931 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S 0.011494f
C1932 a_8802_31196# SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.066256f
C1933 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.363295f
C1934 a_22790_41880# SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.071756f
C1935 SUNSAR_CAPT8B_CV_0.XA5.B a_23942_41352# 0.066018f
C1936 SUNSAR_SAR8B_CV_0.XA20.CNO a_5130_27500# 0.066018f
C1937 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S 0.050207f
C1938 SUNSAR_SAR8B_CV_0.XA2.XA11.A VPWR 0.725614f
C1939 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.175629f
C1940 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.024423f
C1941 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23922_34892# 0.010409f
C1942 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_20250_27148# 0.03422f
C1943 SUNSAR_SAR8B_CV_0.SARN ua[1] 0.806872f
C1944 SUNSAR_SAR8B_CV_0.XA5.XA10.A a_15210_35948# 0.068853f
C1945 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_42760# 0.031082f
C1946 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S 0.016689f
C1947 SUNSAR_SAR8B_CV_0.XB2.CKN a_16542_4038# 0.135393f
C1948 a_13842_28908# VPWR 0.395394f
C1949 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_22770_34540# 0.076663f
C1950 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.026455f
C1951 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S 0.050207f
C1952 ui_in[0] rst_n 0.023911f
C1953 uio_out[3] uio_out[2] 0.023797f
C1954 SUNSAR_SAR8B_CV_0.XA20.CPO a_6282_28908# 0.086948f
C1955 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.012223f
C1956 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA5.CEIN 0.019713f
C1957 tt_um_TT06_SAR_done_0.DONE a_22790_40296# 0.026542f
C1958 a_5130_34716# VPWR 0.399819f
C1959 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_16362_28204# 0.067588f
C1960 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S a_15210_28204# 0.04865f
C1961 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.078539f
C1962 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S 0.050207f
C1963 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S 0.016767f
C1964 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.127551f
C1965 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA20.CNO 2.96993f
C1966 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.010335f
C1967 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S VPWR 0.106927f
C1968 SUNSAR_CAPT8B_CV_0.XD09.XA7.C uo_out[5] 0.245678f
C1969 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G a_9990_5270# 0.072258f
C1970 a_11142_5622# a_11142_5270# 0.010937f
C1971 SUNSAR_SAR8B_CV_0.XA6.XA9.B a_18882_34716# 0.023982f
C1972 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S 0.055045f
C1973 a_23922_26796# VPWR 0.442318f
C1974 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C1975 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_4688# 0.172147f
C1976 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA20.CPO 0.328435f
C1977 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.145048f
C1978 a_22790_42760# SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.069971f
C1979 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S 0.050207f
C1980 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.024782f
C1981 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S 0.062799f
C1982 SUNSAR_SAR8B_CV_0.XA4.EN a_12690_27500# 0.085451f
C1983 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.SARP 0.046452f
C1984 SUNSAR_SAR8B_CV_0.XA20.CNO a_12690_29612# 0.090551f
C1985 a_16382_41352# a_16382_41000# 0.010937f
C1986 a_15210_37180# a_15210_36828# 0.010937f
C1987 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_11322_33836# 0.07476f
C1988 a_5130_31196# VPWR 0.44007f
C1989 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_41880# 0.031087f
C1990 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.301485f
C1991 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S 0.030434f
C1992 SUNSAR_SAR8B_CV_0.EN a_8802_28908# 0.074323f
C1993 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VPWR 0.036745f
C1994 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.SARN 0.056701f
C1995 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.031841f
C1996 a_7650_31196# SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.067588f
C1997 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S VPWR 0.106927f
C1998 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.01291f
C1999 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.075756f
C2000 SUNSAR_CAPT8B_CV_0.XA5.B a_22790_41352# 0.088634f
C2001 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S 0.010193f
C2002 SUNSAR_SAR8B_CV_0.XA20.CNO a_3762_27500# 0.067588f
C2003 SUNSAR_SAR8B_CV_0.XA1.XA11.A VPWR 0.722887f
C2004 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S a_18882_27852# 0.04865f
C2005 a_22770_36300# a_22770_35948# 0.010937f
C2006 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S 0.016683f
C2007 SUNSAR_SAR8B_CV_0.D<5> a_8802_32076# 0.020342f
C2008 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_3686# 0.16579f
C2009 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3334# 0.163985f
C2010 SUNSAR_SAR8B_CV_0.XB2.CKN a_15390_4038# 0.081275f
C2011 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.CP0 0.010925f
C2012 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.011022f
C2013 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.026917f
C2014 a_12582_3334# ua[1] 0.060039f
C2015 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_13842_32076# 0.06801f
C2016 SUNSAR_SAR8B_CV_0.XA6.EN a_17730_29612# 0.074595f
C2017 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_SAR8B_CV_0.D<4> 0.010401f
C2018 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S 0.050207f
C2019 ui_in[0] ui_in[1] 0.024013f
C2020 a_28727_40307# VPWR 0.410063f
C2021 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S 0.030434f
C2022 a_10190_40648# a_10190_40296# 0.010937f
C2023 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.178114f
C2024 tt_um_TT06_SAR_done_0.DONE a_21422_40296# 0.042653f
C2025 a_3762_34716# VPWR 0.399819f
C2026 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_15210_28204# 0.096735f
C2027 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S 0.064105f
C2028 SUNSAR_SAR8B_CV_0.XA1.XA11.A a_6282_36300# 0.13402f
C2029 SUNSAR_CAPT8B_CV_0.XD09.XA7.C uo_out[6] 0.010011f
C2030 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR 0.104609f
C2031 SUNSAR_SAR8B_CV_0.XA6.XA9.B a_17730_34716# 0.047651f
C2032 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_11342_41000# 0.115667f
C2033 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_4848# 0.024512f
C2034 SUNSAR_SAR8B_CV_0.XA2.EN a_7650_30316# 0.070731f
C2035 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.693521f
C2036 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA20.CNO 0.056065f
C2037 a_11342_42760# a_11342_42408# 0.010937f
C2038 SUNSAR_CAPT8B_CV_0.XF11.QN a_13862_43816# 0.091063f
C2039 a_21422_44168# a_21422_43816# 0.010937f
C2040 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S 0.050207f
C2041 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.SARP 0.062345f
C2042 SUNSAR_SAR8B_CV_0.XA20.CNO a_11322_29612# 0.095246f
C2043 SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR 1.2202f
C2044 a_13842_28908# a_13842_28556# 0.010937f
C2045 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.DONE 0.02194f
C2046 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.293159f
C2047 SUNSAR_SAR8B_CV_0.XA1.CEIN a_6282_36828# 0.0733f
C2048 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_7670_41880# 0.072448f
C2049 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1615f
C2050 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_13862_42760# 0.113305f
C2051 a_3762_31196# VPWR 0.44007f
C2052 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.026506f
C2053 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_8802_35420# 0.133834f
C2054 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.010335f
C2055 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VPWR 0.036745f
C2056 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.014291f
C2057 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.449584f
C2058 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C2059 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S 0.077008f
C2060 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S VPWR 0.106927f
C2061 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H 0.057478f
C2062 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.SARP 5.25248f
C2063 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C2064 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<1> 0.077821f
C2065 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S 0.011542f
C2066 SUNSAR_SAR8B_CV_0.XA20.CNO a_2610_27500# 0.066018f
C2067 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR 0.101979f
C2068 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.ENO 0.116058f
C2069 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.029317f
C2070 a_15210_33836# VPWR 0.409601f
C2071 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_13842_35948# 0.070424f
C2072 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S 0.03516f
C2073 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.230205f
C2074 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_12690_32076# 0.088002f
C2075 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S 0.050207f
C2076 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.040072f
C2077 uio_out[4] uio_out[3] 0.023797f
C2078 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_3782_43288# 0.031221f
C2079 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S 0.030434f
C2080 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S 0.030434f
C2081 tt_um_TT06_SAR_done_0.DONE a_20270_40296# 0.026182f
C2082 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31301f
C2083 SUNSAR_SAR8B_CV_0.XA1.XA11.A a_5130_36300# 0.089492f
C2084 SUNSAR_CAPT8B_CV_0.XA6.XA2.A clk 0.037336f
C2085 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN VPWR 1.7759f
C2086 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S uo_out[6] 0.01183f
C2087 a_16542_5974# a_16542_5622# 0.010937f
C2088 a_9990_5622# a_9990_5270# 0.010937f
C2089 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_10190_41000# 0.156079f
C2090 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N VPWR 0.271482f
C2091 a_21402_35420# a_21402_35068# 0.010937f
C2092 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9054_4848# 0.024512f
C2093 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.014291f
C2094 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C2095 a_21422_42760# SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.071391f
C2096 SUNSAR_CAPT8B_CV_0.XF11.QN a_12710_43816# 0.127669f
C2097 TIE_L SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.039224f
C2098 SUNSAR_SAR8B_CV_0.XA3.EN a_11322_27500# 0.082231f
C2099 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S 0.030434f
C2100 a_15230_41352# VPWR 0.394053f
C2101 SUNSAR_SAR8B_CV_0.XA20.CNO a_10170_29612# 0.011704f
C2102 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_27500# 0.044989f
C2103 a_15230_41352# a_15230_41000# 0.010937f
C2104 SUNSAR_SAR8B_CV_0.XA3.XA9.B VPWR 0.93081f
C2105 a_13842_37180# a_13842_36828# 0.010937f
C2106 SUNSAR_SAR8B_CV_0.XA0.XA12.A a_3762_36828# 0.091063f
C2107 SUNSAR_SAR8B_CV_0.XA1.CEIN a_5130_36828# 0.07472f
C2108 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA6.CEIN 0.432008f
C2109 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_12710_42760# 0.089774f
C2110 SUNSAR_SAR8B_CV_0.XA2.XA9.A a_7650_35420# 0.160931f
C2111 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.016772f
C2112 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.527529f
C2113 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S VPWR 0.065445f
C2114 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.204048f
C2115 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_28556# 0.073834f
C2116 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.316693f
C2117 a_6282_31196# SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.066018f
C2118 SUNSAR_SAR8B_CV_0.XA20.CNO a_21402_27852# 0.072527f
C2119 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR 0.119314f
C2120 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.024478f
C2121 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.849501f
C2122 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.EN 0.111173f
C2123 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_18882_27148# 0.03422f
C2124 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S a_7650_27500# 0.036993f
C2125 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S a_17730_27852# 0.056787f
C2126 SUNSAR_SAR8B_CV_0.SARP a_12582_3334# 0.038089f
C2127 a_13842_33836# VPWR 0.409601f
C2128 a_21402_36300# a_21402_35948# 0.010937f
C2129 SUNSAR_SAR8B_CV_0.XA4.XA10.A a_12690_35948# 0.132671f
C2130 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.016334f
C2131 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.26479f
C2132 a_10170_28908# VPWR 0.395394f
C2133 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.011022f
C2134 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.026917f
C2135 a_13950_3686# ua[0] 0.067632f
C2136 SUNSAR_SAR8B_CV_0.XA5.EN a_16362_29612# 0.073155f
C2137 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S 0.050207f
C2138 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.233892f
C2139 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_3782_43288# 0.080718f
C2140 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_43288# 0.069053f
C2141 tt_um_TT06_SAR_done_0.x3.MP1.G VPWR 0.695784f
C2142 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S 0.050207f
C2143 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.012023f
C2144 SUNSAR_SAR8B_CV_0.XA20.CPO a_2610_28908# 0.085247f
C2145 a_8822_40648# a_8822_40296# 0.010937f
C2146 tt_um_TT06_SAR_done_0.DONE a_18902_40296# 0.026182f
C2147 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR 3.91346f
C2148 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S a_13842_28204# 0.04865f
C2149 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S 0.050207f
C2150 SUNSAR_SAR8B_CV_0.SARN m1_14848_7490# 0.031022f
C2151 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.CN1 0.033978f
C2152 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.072558f
C2153 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.077804f
C2154 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.021174f
C2155 SUNSAR_CAPT8B_CV_0.XD09.XA7.C VPWR 2.97208f
C2156 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S uo_out[6] 0.023976f
C2157 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_18902_41352# 0.058557f
C2158 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C2159 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.093524f
C2160 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2502_5648# 0.0666f
C2161 a_20250_26796# VPWR 0.441753f
C2162 SUNSAR_SAR8B_CV_0.XA1.EN a_6282_30316# 0.06916f
C2163 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C2164 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.090222f
C2165 a_21402_33836# SUNSAR_SAR8B_CV_0.XA7.CP0 0.066219f
C2166 a_10190_42760# a_10190_42408# 0.010937f
C2167 a_20270_42760# SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.067588f
C2168 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.015882f
C2169 a_20270_44168# a_20270_43816# 0.010937f
C2170 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S 0.050207f
C2171 a_13862_41352# VPWR 0.394053f
C2172 SUNSAR_CAPT8B_CV_0.XA4.MP1.G clk 0.438597f
C2173 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S 0.050207f
C2174 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.375196f
C2175 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S 0.050207f
C2176 SUNSAR_SAR8B_CV_0.XA20.CNO a_8802_29612# 0.011248f
C2177 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.55251f
C2178 SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR 1.22023f
C2179 a_12690_28908# a_12690_28556# 0.010937f
C2180 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.158152f
C2181 SUNSAR_SAR8B_CV_0.XA0.XA12.A a_2610_36828# 0.10248f
C2182 SUNSAR_SAR8B_CV_0.XA1.CEIN a_3762_36828# 0.015625f
C2183 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_7650_33836# 0.073189f
C2184 SUNSAR_SAR8B_CV_0.XA20.CNO VPWR 6.94539f
C2185 a_21402_27500# a_21402_27148# 0.010937f
C2186 SUNSAR_SAR8B_CV_0.EN a_5130_28908# 0.072753f
C2187 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S 0.023798f
C2188 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S VPWR 0.066675f
C2189 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 0.026917f
C2190 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.126806f
C2191 a_5130_31196# SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.067827f
C2192 a_23942_42408# VPWR 0.3915f
C2193 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.702226f
C2194 SUNSAR_SAR8B_CV_0.XA20.CNO a_20250_27852# 0.067588f
C2195 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S 0.050207f
C2196 SUNSAR_SAR8B_CV_0.XA0.XA11.A VPWR 0.728421f
C2197 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.024423f
C2198 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.EN 0.893904f
C2199 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.EN 0.111217f
C2200 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_17730_27148# 0.023111f
C2201 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_3782_42760# 0.031082f
C2202 SUNSAR_SAR8B_CV_0.D<0> a_20250_32956# 0.017876f
C2203 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S 0.044153f
C2204 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.379175p
C2205 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.669708f
C2206 a_8802_28908# VPWR 0.395394f
C2207 a_13950_4390# a_13950_4038# 0.010937f
C2208 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.016471f
C2209 a_9990_2630# VPWR 0.447601f
C2210 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_11322_32076# 0.089573f
C2211 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S 0.050207f
C2212 uio_out[5] uio_out[4] 0.023797f
C2213 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S 0.036094f
C2214 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_2630_43288# 0.028213f
C2215 a_28727_40659# VPWR 0.39147f
C2216 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S 0.027953f
C2217 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.179089f
C2218 tt_um_TT06_SAR_done_0.DONE a_17750_40296# 0.042794f
C2219 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.027044f
C2220 a_23922_34892# VPWR 0.395601f
C2221 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_13842_28204# 0.098305f
C2222 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S 0.064105f
C2223 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.CN1 0.024218f
C2224 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S 0.028452f
C2225 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.010335f
C2226 SUNSAR_CAPT8B_CV_0.XC08.XA7.C uo_out[6] 0.251051f
C2227 a_15390_5974# a_15390_5622# 0.010937f
C2228 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_18902_41352# 0.075505f
C2229 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_41352# 0.060327f
C2230 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S 0.089305f
C2231 a_20250_35420# a_20250_35068# 0.010937f
C2232 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_5648# 0.172147f
C2233 a_18882_26796# VPWR 0.442908f
C2234 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.014291f
C2235 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C2236 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.041437f
C2237 a_20250_33836# SUNSAR_SAR8B_CV_0.XA7.CP0 0.067588f
C2238 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43816# 0.129239f
C2239 SUNSAR_SAR8B_CV_0.XA20.CNO a_7650_29612# 0.090551f
C2240 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_27500# 0.054233f
C2241 a_13862_41352# a_13862_41000# 0.010937f
C2242 tt_um_TT06_SAR_done_0.DONE a_23922_35948# 0.066018f
C2243 a_12690_37180# a_12690_36828# 0.010937f
C2244 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_6282_33836# 0.07476f
C2245 a_23922_31724# VPWR 0.412398f
C2246 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.301485f
C2247 SUNSAR_SAR8B_CV_0.EN a_3762_28908# 0.074323f
C2248 SUNSAR_SAR8B_CV_0.XA2.XA9.B a_7650_35420# 0.017683f
C2249 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VPWR 0.036745f
C2250 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C2251 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.15651f
C2252 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S 0.011494f
C2253 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_28556# 0.075865f
C2254 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S 0.076247f
C2255 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_5094# 0.16149f
C2256 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<2> 0.086175f
C2257 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.586025f
C2258 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<3> 0.083397f
C2259 SUNSAR_SAR8B_CV_0.XA20.CNO a_18882_27852# 0.066018f
C2260 SUNSAR_SAR8B_CV_0.XB2.TIE_L VPWR 11.0126f
C2261 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N a_21402_28908# 0.060353f
C2262 SUNSAR_SAR8B_CV_0.SARN a_12582_4742# 0.044957f
C2263 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.EN 0.952619f
C2264 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.EN 0.111173f
C2265 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S a_6282_27500# 0.036993f
C2266 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S a_16362_27852# 0.056787f
C2267 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_42760# 0.031591f
C2268 a_20250_36300# a_20250_35948# 0.010937f
C2269 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_11322_35948# 0.134161f
C2270 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S 0.044228f
C2271 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3686# 0.16579f
C2272 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.CP0 0.010925f
C2273 a_3762_34716# SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.068712f
C2274 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C2275 a_16542_2982# VPWR 0.490338f
C2276 a_12582_3686# ua[1] 0.067632f
C2277 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B ua[0] 0.241597f
C2278 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_10170_32076# 0.066439f
C2279 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_SAR8B_CV_0.D<5> 0.010401f
C2280 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S 0.050207f
C2281 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S 0.030434f
C2282 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.010898f
C2283 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S 0.0111f
C2284 a_7670_40648# a_7670_40296# 0.010937f
C2285 tt_um_TT06_SAR_done_0.DONE a_16382_40296# 0.042794f
C2286 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA4.CEIN 0.05126f
C2287 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_12690_28204# 0.066018f
C2288 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.078539f
C2289 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.CN1 0.024049f
C2290 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN uo_out[6] 0.306905f
C2291 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S VPWR 0.106927f
C2292 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR 0.104609f
C2293 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_17750_41352# 0.080002f
C2294 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_SAR8B_CV_0.D<6> 0.018133f
C2295 SUNSAR_SAR8B_CV_0.XA5.XA9.B a_16362_34716# 0.047651f
C2296 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_5808# 0.024512f
C2297 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.090222f
C2298 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C2299 a_8822_42760# a_8822_42408# 0.010937f
C2300 a_18902_42760# SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.066018f
C2301 SUNSAR_CAPT8B_CV_0.XE10.QN a_10190_43816# 0.089492f
C2302 a_18902_44168# a_18902_43816# 0.010937f
C2303 SUNSAR_SAR8B_CV_0.XA20.CNO a_6282_29612# 0.095246f
C2304 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S 0.050207f
C2305 SUNSAR_SAR8B_CV_0.D<0> clk 0.012554f
C2306 SUNSAR_SAR8B_CV_0.XA2.XA9.B VPWR 0.930839f
C2307 a_11322_28908# a_11322_28556# 0.010937f
C2308 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.220689f
C2309 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.DONE 0.054848f
C2310 tt_um_TT06_SAR_done_0.DONE a_22770_35948# 0.075373f
C2311 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6519f
C2312 a_20250_27500# a_20250_27148# 0.010937f
C2313 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.026506f
C2314 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_6302_41880# 0.070877f
C2315 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VPWR 0.036745f
C2316 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B 0.026917f
C2317 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C2318 SUNSAR_SAR8B_CV_0.XA7.EN a_17730_28556# 0.132757f
C2319 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.363295f
C2320 a_3762_31196# SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.066256f
C2321 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.702226f
C2322 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA20.CPO 0.255261f
C2323 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_5094# 0.161108f
C2324 SUNSAR_SAR8B_CV_0.XA20.CNO a_17730_27852# 0.074163f
C2325 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N a_20250_28908# 0.023475f
C2326 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.029312f
C2327 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.EN 1.02916f
C2328 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.EN 0.111217f
C2329 a_10170_33836# VPWR 0.409601f
C2330 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.230084f
C2331 SUNSAR_SAR8B_CV_0.XA3.XA10.A a_10170_35948# 0.068853f
C2332 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.038188f
C2333 a_12582_4390# a_12582_4038# 0.010937f
C2334 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.143148f
C2335 SUNSAR_SAR8B_CV_0.XA7.XA9.B a_20250_33836# 0.023316f
C2336 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S ua[0] 0.100365f
C2337 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S 0.050207f
C2338 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.040072f
C2339 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S 0.024386f
C2340 uio_out[6] uio_out[5] 0.023797f
C2341 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S 0.073313f
C2342 tt_um_TT06_SAR_done_0.x4.MP0.G VPWR 0.511762f
C2343 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N a_12690_29612# 0.031412f
C2344 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S 0.026417f
C2345 tt_um_TT06_SAR_done_0.DONE a_15230_40296# 0.026182f
C2346 SUNSAR_SAR8B_CV_0.XA7.ENO VPWR 4.77251f
C2347 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.CKN 0.169642f
C2348 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.55251f
C2349 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.CN1 0.024049f
C2350 SUNSAR_SAR8B_CV_0.XA0.XA11.A a_3762_36300# 0.091063f
C2351 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.073199f
C2352 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.075983f
C2353 a_20270_43816# uo_out[0] 0.022673f
C2354 SUNSAR_CAPT8B_CV_0.XC08.XA7.C VPWR 2.97221f
C2355 a_18882_35420# a_18882_35068# 0.010937f
C2356 SUNSAR_SAR8B_CV_0.XA5.XA9.B a_15210_34716# 0.023982f
C2357 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2502_2768# 0.024512f
C2358 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.026917f
C2359 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C2360 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9054_5808# 0.024512f
C2361 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.04064f
C2362 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C2363 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.59085f
C2364 a_18882_33836# SUNSAR_SAR8B_CV_0.XA6.CP0 0.066018f
C2365 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.28707f
C2366 a_17750_42760# SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.072962f
C2367 a_23942_43992# SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.033775f
C2368 SUNSAR_SAR8B_CV_0.XA20.CNO a_5130_29612# 0.011704f
C2369 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.010898f
C2370 a_10190_41352# VPWR 0.394053f
C2371 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S 0.050207f
C2372 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.383512f
C2373 SUNSAR_SAR8B_CV_0.XA2.EN a_7650_27500# 0.085451f
C2374 SUNSAR_SAR8B_CV_0.D<0> ui_in[0] 0.013f
C2375 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_27852# 0.024578f
C2376 a_12710_41352# a_12710_41000# 0.010937f
C2377 a_21402_37180# SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.069366f
C2378 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA5.CEIN 0.033943f
C2379 a_11322_37180# a_11322_36828# 0.010937f
C2380 SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR 2.62715f
C2381 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S 0.030434f
C2382 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_20270_42408# 0.076129f
C2383 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_21422_42408# 0.098561f
C2384 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_6302_41880# 0.031087f
C2385 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_11342_42760# 0.091344f
C2386 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S VPWR 0.065445f
C2387 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.380687f
C2388 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S 0.028026f
C2389 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S 0.013533f
C2390 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.204048f
C2391 a_20270_42408# VPWR 0.391292f
C2392 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.267238f
C2393 a_2610_31196# SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.067588f
C2394 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.024478f
C2395 SUNSAR_SAR8B_CV_0.XA20.CNO a_16362_27852# 0.072592f
C2396 a_20250_36828# VPWR 0.392512f
C2397 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.EN 0.111173f
C2398 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.EN 0.952619f
C2399 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_16362_27148# 0.023111f
C2400 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S a_15210_27852# 0.04865f
C2401 a_8802_33836# VPWR 0.409601f
C2402 SUNSAR_SAR8B_CV_0.SARP a_12582_3686# 0.045463f
C2403 SUNSAR_SAR8B_CV_0.D<6> a_5130_32076# 0.020342f
C2404 a_18882_36300# a_18882_35948# 0.010937f
C2405 a_5130_28908# VPWR 0.395394f
C2406 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_16542_4038# 0.034677f
C2407 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.161963f
C2408 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.40569f
C2409 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.440586f
C2410 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_8802_32076# 0.06801f
C2411 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.012886f
C2412 SUNSAR_SAR8B_CV_0.XA4.EN a_12690_29612# 0.074595f
C2413 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.CPO 0.096247f
C2414 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CNO 0.084573f
C2415 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S 0.050207f
C2416 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.63636f
C2417 VPWR ua[7] 0.010285f
C2418 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.B 0.342913f
C2419 a_23942_40296# VPWR 0.455498f
C2420 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S 0.050207f
C2421 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S 0.010745f
C2422 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CEIN 0.075193f
C2423 a_6302_40648# a_6302_40296# 0.010937f
C2424 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.178114f
C2425 tt_um_TT06_SAR_done_0.DONE a_13862_40296# 0.026182f
C2426 SUNSAR_SAR8B_CV_0.XA7.EN VPWR 5.54203f
C2427 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.CN1 0.024049f
C2428 SUNSAR_SAR8B_CV_0.XA0.XA11.A a_2610_36300# 0.13253f
C2429 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.010854f
C2430 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S uo_out[7] 0.024266f
C2431 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR 0.042839f
C2432 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN VPWR 1.7759f
C2433 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.SARP 0.05058f
C2434 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S 0.055045f
C2435 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2358_2768# 0.049023f
C2436 a_15210_26796# VPWR 0.441753f
C2437 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2502_6608# 0.0666f
C2438 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA20.CNO 0.056415f
C2439 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.090222f
C2440 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C2441 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.26071f
C2442 a_17730_33836# SUNSAR_SAR8B_CV_0.XA6.CP0 0.067789f
C2443 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.092023f
C2444 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_20270_42408# 0.015723f
C2445 a_7670_42760# a_7670_42408# 0.010937f
C2446 a_22790_43992# SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.030547f
C2447 SUNSAR_CAPT8B_CV_0.XD09.QN a_8822_43816# 0.091063f
C2448 TIE_L SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.039224f
C2449 a_17750_44168# a_17750_43816# 0.010937f
C2450 SUNSAR_SAR8B_CV_0.XA20.CNO a_3762_29612# 0.011248f
C2451 a_8822_41352# VPWR 0.394053f
C2452 SUNSAR_SAR8B_CV_0.D<0> tt_um_TT06_SAR_done_0.DONE 0.490252f
C2453 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B 3.55251f
C2454 SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR 1.2202f
C2455 a_10170_28908# a_10170_28556# 0.010937f
C2456 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_2610_33836# 0.073189f
C2457 a_20250_37180# SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.067588f
C2458 a_21402_37180# SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.033775f
C2459 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.377598f
C2460 SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR 2.62331f
C2461 a_18882_27500# a_18882_27148# 0.010937f
C2462 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_42408# 0.031125f
C2463 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_41880# 0.100592f
C2464 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_10190_42760# 0.111734f
C2465 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S 0.027192f
C2466 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S 0.010335f
C2467 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.046858f
C2468 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_6282_35420# 0.160931f
C2469 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C2470 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S VPWR 0.066675f
C2471 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.071907f
C2472 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.SARN 0.064384f
C2473 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.038766f
C2474 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_28556# 0.135353f
C2475 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_15390_5270# 0.012993f
C2476 a_18902_42408# VPWR 0.391292f
C2477 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.702226f
C2478 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.109021f
C2479 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<3> 0.073432f
C2480 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C2481 SUNSAR_SAR8B_CV_0.XA20.CPO a_21402_28204# 0.088691f
C2482 SUNSAR_SAR8B_CV_0.XA20.CNO a_15210_27852# 0.067588f
C2483 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S 0.050207f
C2484 a_18882_36828# VPWR 0.395703f
C2485 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.EN 1.02916f
C2486 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.EN 0.111217f
C2487 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_15210_27148# 0.03422f
C2488 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_8802_35948# 0.070424f
C2489 SUNSAR_SAR8B_CV_0.D<1> a_18882_32956# 0.017466f
C2490 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S 0.03516f
C2491 a_3762_28908# VPWR 0.395394f
C2492 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.CKN 0.011708f
C2493 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.016334f
C2494 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.059977f
C2495 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B ua[1] 0.241597f
C2496 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_7650_32076# 0.088002f
C2497 SUNSAR_SAR8B_CV_0.XA20.XA3.CO a_23922_31724# 0.010987f
C2498 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S 0.050207f
C2499 a_23942_42408# SUNSAR_CAPT8B_CV_0.XA5.B 0.066018f
C2500 uio_out[7] uio_out[6] 0.023797f
C2501 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_23942_43640# 0.070424f
C2502 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S 0.024389f
C2503 tt_um_TT06_SAR_done_0.DONE a_12710_40296# 0.042794f
C2504 SUNSAR_SAR8B_CV_0.XA6.EN VPWR 4.84607f
C2505 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_11322_28204# 0.067588f
C2506 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S a_10170_28204# 0.04865f
C2507 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S 0.028448f
C2508 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.099766f
C2509 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.010335f
C2510 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S uo_out[7] 0.012119f
C2511 a_18902_43816# uo_out[1] 0.022673f
C2512 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR 0.042839f
C2513 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S VPWR 0.106927f
C2514 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.300065f
C2515 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_8822_41000# 0.15757f
C2516 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.024853f
C2517 a_17730_35420# a_17730_35068# 0.010937f
C2518 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S 0.089305f
C2519 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S 0.026506f
C2520 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S 0.097398f
C2521 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_2928# 0.105547f
C2522 a_13842_26796# VPWR 0.442908f
C2523 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.026917f
C2524 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C2525 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_6608# 0.172147f
C2526 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 1.8915f
C2527 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.036726f
C2528 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.041437f
C2529 a_16382_42760# SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.071391f
C2530 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C2531 SUNSAR_SAR8B_CV_0.XA1.EN a_6282_27500# 0.082231f
C2532 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_27500# 0.044989f
C2533 SUNSAR_SAR8B_CV_0.XA20.CNO a_2610_29612# 0.090485f
C2534 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_27852# 0.025674f
C2535 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S 0.062799f
C2536 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S 0.050207f
C2537 a_11342_41352# a_11342_41000# 0.010937f
C2538 SUNSAR_SAR8B_CV_0.XA1.XA9.B VPWR 0.93081f
C2539 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.SARN 0.108405f
C2540 a_20250_37180# SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.030547f
C2541 a_10170_37180# a_10170_36828# 0.010937f
C2542 SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR 2.62344f
C2543 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S 0.023798f
C2544 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.126085f
C2545 SUNSAR_SAR8B_CV_0.XA1.XA9.B a_6282_35420# 0.017683f
C2546 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_5130_35420# 0.133834f
C2547 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VPWR 0.036745f
C2548 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C2549 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S 0.013533f
C2550 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_28556# 0.073834f
C2551 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_11142_5270# 0.012993f
C2552 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.SARP 0.036512f
C2553 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<5> 0.010193f
C2554 SUNSAR_SAR8B_CV_0.XA20.CPO a_20250_28204# 0.068716f
C2555 SUNSAR_SAR8B_CV_0.XA20.CNO a_13842_27852# 0.066018f
C2556 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.EN 0.111173f
C2557 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.EN 0.952619f
C2558 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S a_13842_27852# 0.04865f
C2559 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.EN 0.058308f
C2560 a_17730_36300# a_17730_35948# 0.010937f
C2561 SUNSAR_SAR8B_CV_0.XA2.XA10.A a_7650_35948# 0.132671f
C2562 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.038188f
C2563 SUNSAR_SAR8B_CV_0.XB2.XA4.GN a_13950_4038# 0.070815f
C2564 SUNSAR_SAR8B_CV_0.XB1.CKN a_11142_4038# 0.082845f
C2565 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.CP0 0.010925f
C2566 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.02165f
C2567 a_16542_4038# ua[0] 0.023111f
C2568 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S ua[1] 0.100365f
C2569 SUNSAR_SAR8B_CV_0.XA3.EN a_11322_29612# 0.073155f
C2570 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.034212f
C2571 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_SAR8B_CV_0.D<6> 0.010401f
C2572 a_22790_42408# SUNSAR_CAPT8B_CV_0.XA5.B 0.072519f
C2573 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S 0.050207f
C2574 SUNSAR_CAPT8B_CV_0.XA6.XA2.A a_22790_43640# 0.127669f
C2575 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S 0.026257f
C2576 a_5150_40648# a_5150_40296# 0.010937f
C2577 tt_um_TT06_SAR_done_0.DONE a_11342_40296# 0.042794f
C2578 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.030806f
C2579 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S 0.073693f
C2580 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_10170_28204# 0.096735f
C2581 a_21402_28556# a_21402_28204# 0.010937f
C2582 SUNSAR_SAR8B_CV_0.XA5.EN VPWR 5.52623f
C2583 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.081322f
C2584 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.077366f
C2585 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.09742f
C2586 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.019775f
C2587 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S 0.016769f
C2588 SUNSAR_SAR8B_CV_0.XA20.CK_CMP a_23922_36300# 0.066062f
C2589 a_11142_5622# SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G 0.066018f
C2590 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN uo_out[7] 0.308722f
C2591 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N VPWR 0.271482f
C2592 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_7670_41000# 0.114097f
C2593 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_13862_41880# 0.072658f
C2594 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_16382_41352# 0.078431f
C2595 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S 0.055045f
C2596 SUNSAR_SAR8B_CV_0.XA20.XA11.Y a_23922_34892# 0.067588f
C2597 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.023301f
C2598 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.093524f
C2599 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9054_2928# 0.0666f
C2600 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_6768# 0.024512f
C2601 a_16362_33836# SUNSAR_SAR8B_CV_0.XA5.CP0 0.066219f
C2602 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.090222f
C2603 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.431957f
C2604 a_15230_42760# SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.067588f
C2605 a_6302_42760# a_6302_42408# 0.010937f
C2606 a_16382_44168# a_16382_43816# 0.010937f
C2607 SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR 1.22398f
C2608 a_8802_28908# a_8802_28556# 0.010937f
C2609 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S 0.053284f
C2610 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.DONE 0.02194f
C2611 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.293159f
C2612 a_17730_27500# a_17730_27148# 0.010937f
C2613 SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR 2.62344f
C2614 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.55251f
C2615 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S 0.027192f
C2616 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.527529f
C2617 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C2618 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VPWR 0.036745f
C2619 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.113828f
C2620 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_21402_30316# 0.01727f
C2621 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.702226f
C2622 SUNSAR_SAR8B_CV_0.XA20.CPO a_18882_28204# 0.067146f
C2623 SUNSAR_SAR8B_CV_0.XA20.CNO a_12690_27852# 0.074163f
C2624 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.029317f
C2625 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.EN 1.04628f
C2626 a_5130_33836# VPWR 0.409601f
C2627 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S 0.016689f
C2628 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.230325f
C2629 SUNSAR_SAR8B_CV_0.XB1.CKN a_9990_4038# 0.135393f
C2630 SUNSAR_SAR8B_CV_0.XA6.XA9.B a_18882_33836# 0.023316f
C2631 a_15390_4038# ua[0] 0.043386f
C2632 a_9990_2982# VPWR 0.491909f
C2633 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_6282_32076# 0.089573f
C2634 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S 0.050207f
C2635 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_21422_41880# 0.035868f
C2636 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.040072f
C2637 SUNSAR_CAPT8B_CV_0.XI14.QN a_21422_43288# 0.03616f
C2638 a_20270_40296# VPWR 0.456842f
C2639 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N a_11322_29612# 0.031412f
C2640 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S 0.026117f
C2641 tt_um_TT06_SAR_done_0.DONE a_10190_40296# 0.026182f
C2642 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA3.CEIN 0.019713f
C2643 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 54.2165f
C2644 SUNSAR_SAR8B_CV_0.XA4.EN VPWR 4.84607f
C2645 SUNSAR_SAR8B_CV_0.XA20.CK_CMP a_22770_36300# 0.078456f
C2646 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN VPWR 1.7759f
C2647 a_9990_5622# SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G 0.098184f
C2648 SUNSAR_CAPT8B_CV_0.XB07.XA7.C uo_out[7] 0.248979f
C2649 SUNSAR_SAR8B_CV_0.XA20.XA11.Y a_22770_34892# 0.069969f
C2650 a_16362_35420# a_16362_35068# 0.010937f
C2651 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.SARP 0.046484f
C2652 SUNSAR_SAR8B_CV_0.XA4.XA9.B a_13842_34716# 0.023982f
C2653 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_12710_41880# 0.066018f
C2654 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_16382_41352# 0.060327f
C2655 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_15230_41352# 0.077076f
C2656 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2502_3728# 0.024512f
C2657 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.021241f
C2658 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.098257f
C2659 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9054_6768# 0.024512f
C2660 a_15210_33836# SUNSAR_SAR8B_CV_0.XA5.CP0 0.067588f
C2661 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.04064f
C2662 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.07159f
C2663 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C2664 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_27500# 0.054233f
C2665 a_5150_41352# VPWR 0.394053f
C2666 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.018975f
C2667 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S 0.062799f
C2668 a_10190_41352# a_10190_41000# 0.010937f
C2669 SUNSAR_SAR8B_CV_0.D<1> tt_um_TT06_SAR_done_0.DONE 0.295407f
C2670 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S 0.022628f
C2671 a_18882_37180# SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.066018f
C2672 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA4.CEIN 0.432008f
C2673 a_8802_37180# a_8802_36828# 0.010937f
C2674 SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR 2.62344f
C2675 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S VPWR 0.065445f
C2676 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C2677 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_28556# 0.075865f
C2678 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G 0.08427f
C2679 a_15230_42408# VPWR 0.391292f
C2680 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<4> 0.073463f
C2681 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<5> 1.62763f
C2682 SUNSAR_SAR8B_CV_0.XA20.CPO a_17730_28204# 0.09022f
C2683 SUNSAR_SAR8B_CV_0.XA20.CNO a_11322_27852# 0.072592f
C2684 a_15210_36828# VPWR 0.395582f
C2685 a_3762_33836# VPWR 0.409601f
C2686 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_13842_27148# 0.03422f
C2687 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S a_2610_27500# 0.036993f
C2688 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S a_12690_27852# 0.056787f
C2689 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S 0.016683f
C2690 a_16362_36300# a_16362_35948# 0.010937f
C2691 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_6282_35948# 0.134161f
C2692 SUNSAR_SAR8B_CV_0.D<7> a_3762_32076# 0.066018f
C2693 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR 0.104609f
C2694 SUNSAR_CAPT8B_CV_0.XF11.XA6.A uo_out[3] 0.016067f
C2695 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A a_9990_4038# 0.01736f
C2696 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.089055f
C2697 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_34716# 0.067815f
C2698 a_13950_4038# ua[0] 0.056243f
C2699 a_16542_3334# VPWR 0.380282f
C2700 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_5130_32076# 0.066439f
C2701 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<0> 0.18344f
C2702 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_20270_41880# 0.024901f
C2703 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.060807f
C2704 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S 0.050207f
C2705 SUNSAR_CAPT8B_CV_0.XI14.QN a_20270_43288# 0.024901f
C2706 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S 0.027953f
C2707 a_18902_40296# VPWR 0.458821f
C2708 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S 0.050207f
C2709 a_3782_40648# a_3782_40296# 0.010937f
C2710 tt_um_TT06_SAR_done_0.DONE a_8822_40296# 0.026182f
C2711 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB1.CKN 0.169642f
C2712 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S a_8802_28204# 0.04865f
C2713 a_20250_28556# a_20250_28204# 0.010937f
C2714 SUNSAR_SAR8B_CV_0.XA3.EN VPWR 5.52623f
C2715 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.073962f
C2716 SUNSAR_CAPT8B_CV_0.XB07.XA7.C VPWR 2.97213f
C2717 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR 0.104609f
C2718 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_SAR8B_CV_0.D<7> 0.018133f
C2719 SUNSAR_SAR8B_CV_0.XA4.XA9.B a_12690_34716# 0.047651f
C2720 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_41352# 0.058557f
C2721 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2358_3728# 0.049023f
C2722 a_10170_26796# VPWR 0.441753f
C2723 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.090222f
C2724 a_5150_42760# a_5150_42408# 0.010937f
C2725 a_13862_42760# SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.066018f
C2726 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_18902_42408# 0.015723f
C2727 a_15230_44168# a_15230_43816# 0.010937f
C2728 SUNSAR_CAPT8B_CV_0.XC08.QN a_5150_43816# 0.089492f
C2729 a_3782_41352# VPWR 0.394053f
C2730 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_27852# 0.010898f
C2731 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 54.2173f
C2732 SUNSAR_SAR8B_CV_0.XA0.XA9.B VPWR 0.94014f
C2733 a_7650_28908# a_7650_28556# 0.010937f
C2734 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.090118f
C2735 a_17730_37180# SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.070936f
C2736 a_18882_37180# SUNSAR_SAR8B_CV_0.XA7.CEIN 0.040807f
C2737 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.158152f
C2738 a_16362_27500# a_16362_27148# 0.010937f
C2739 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR 2.62395f
C2740 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_3782_41880# 0.099022f
C2741 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S 0.027192f
C2742 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_8822_42760# 0.113305f
C2743 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_18902_42408# 0.031125f
C2744 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.DONE 0.049573f
C2745 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_3762_35420# 0.133834f
C2746 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S VPWR 0.066675f
C2747 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C2748 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.702226f
C2749 SUNSAR_CAPT8B_CV_0.XA5.XA2.A clk 0.024024f
C2750 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S 0.011494f
C2751 SUNSAR_SAR8B_CV_0.XA5.EN a_12690_28556# 0.132757f
C2752 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_13950_5446# 0.104059f
C2753 a_13862_42408# VPWR 0.391292f
C2754 SUNSAR_SAR8B_CV_0.XA20.CPO a_16362_28204# 0.088673f
C2755 SUNSAR_SAR8B_CV_0.XA20.CNO a_10170_27852# 0.067588f
C2756 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S 0.050207f
C2757 a_13842_36828# VPWR 0.395703f
C2758 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_12690_27148# 0.023111f
C2759 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S 0.03516f
C2760 SUNSAR_SAR8B_CV_0.XA1.XA10.A a_5130_35948# 0.068853f
C2761 SUNSAR_SAR8B_CV_0.D<7> a_2610_32076# 0.073183f
C2762 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_34716# 0.075712f
C2763 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 0.635098f
C2764 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<0> 0.315965f
C2765 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S 0.050207f
C2766 uio_oe[2] uio_oe[1] 0.023797f
C2767 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S 0.024386f
C2768 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S 0.0111f
C2769 tt_um_TT06_SAR_done_0.DONE a_7670_40296# 0.042794f
C2770 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_8802_28204# 0.098305f
C2771 SUNSAR_SAR8B_CV_0.XA2.EN VPWR 4.84607f
C2772 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.010335f
C2773 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.073275f
C2774 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 2.40935f
C2775 a_15230_43816# uo_out[2] 0.022673f
C2776 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR 0.765792f
C2777 a_11142_5974# a_11142_5622# 0.010937f
C2778 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N VPWR 0.271482f
C2779 a_15210_35420# a_15210_35068# 0.010937f
C2780 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_3888# 0.105547f
C2781 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.021241f
C2782 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.098257f
C2783 a_8802_26796# VPWR 0.442908f
C2784 a_13842_33836# SUNSAR_SAR8B_CV_0.XA4.CP0 0.066018f
C2785 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.041437f
C2786 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.036749f
C2787 a_12710_42760# SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.072962f
C2788 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S 0.013794f
C2789 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_27852# 0.024578f
C2790 a_8822_41352# a_8822_41000# 0.010937f
C2791 a_23922_35948# VPWR 0.390687f
C2792 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.CN0 0.075315f
C2793 a_17730_37180# SUNSAR_SAR8B_CV_0.XA7.CEIN 0.023111f
C2794 a_7650_37180# a_7650_36828# 0.010937f
C2795 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR 2.62405f
C2796 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_41880# 0.031087f
C2797 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA20.CPO 0.074326f
C2798 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S 0.027192f
C2799 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_7670_42760# 0.089774f
C2800 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S 0.030434f
C2801 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_18902_42408# 0.074559f
C2802 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_42408# 0.100131f
C2803 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_2610_35420# 0.160931f
C2804 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.034924f
C2805 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VPWR 0.036745f
C2806 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C2807 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.CP0 0.08098f
C2808 SUNSAR_SAR8B_CV_0.XA7.CN1 a_20250_31196# 0.069193f
C2809 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_12582_5446# 0.102489f
C2810 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S 0.010193f
C2811 SUNSAR_SAR8B_CV_0.XA20.CPO a_15210_28204# 0.068716f
C2812 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N a_18882_28908# 0.023475f
C2813 SUNSAR_SAR8B_CV_0.XA20.CNO a_8802_27852# 0.066018f
C2814 SUNSAR_SAR8B_CV_0.SARN VPWR 0.148723f
C2815 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S a_11322_27852# 0.056787f
C2816 a_21402_28204# a_21402_27852# 0.010937f
C2817 a_15210_36300# a_15210_35948# 0.010937f
C2818 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR 0.104609f
C2819 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_4038# 0.068974f
C2820 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.250503f
C2821 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.CP0 0.010925f
C2822 a_12582_4038# ua[1] 0.056243f
C2823 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.082663f
C2824 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_3762_32076# 0.06801f
C2825 SUNSAR_SAR8B_CV_0.XA2.EN a_7650_29612# 0.074595f
C2826 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_18902_41880# 0.024901f
C2827 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_SAR8B_CV_0.D<7> 0.010401f
C2828 uio_out[0] uio_out[1] 0.023797f
C2829 a_21422_43816# SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.071553f
C2830 SUNSAR_CAPT8B_CV_0.XH13.QN a_18902_43288# 0.024901f
C2831 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S 0.050207f
C2832 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S 0.030434f
C2833 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S 0.025128f
C2834 tt_um_TT06_SAR_done_0.DONE a_6302_40296# 0.042794f
C2835 a_2630_40648# a_2630_40296# 0.010937f
C2836 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S 0.073693f
C2837 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_7650_28204# 0.066018f
C2838 a_18882_28556# a_18882_28204# 0.010937f
C2839 SUNSAR_SAR8B_CV_0.XA1.EN VPWR 5.52718f
C2840 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.079158f
C2841 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.010854f
C2842 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S 0.055045f
C2843 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_6302_41000# 0.115667f
C2844 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C2845 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.SARP 0.049542f
C2846 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9054_3888# 0.0666f
C2847 a_12690_33836# SUNSAR_SAR8B_CV_0.XA4.CP0 0.067789f
C2848 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.090222f
C2849 a_3782_42760# a_3782_42408# 0.010937f
C2850 a_13862_44168# a_13862_43816# 0.010937f
C2851 SUNSAR_CAPT8B_CV_0.XB07.QN a_3782_43816# 0.091063f
C2852 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR 0.635621f
C2853 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S 0.050207f
C2854 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.375196f
C2855 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S 0.050207f
C2856 SUNSAR_SAR8B_CV_0.D<2> tt_um_TT06_SAR_done_0.DONE 0.295646f
C2857 a_6282_28908# a_6282_28556# 0.010937f
C2858 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S 0.022425f
C2859 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.CN0 0.02493f
C2860 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.DONE 0.054848f
C2861 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.220689f
C2862 a_15210_27500# a_15210_27148# 0.010937f
C2863 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.55251f
C2864 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_2630_41880# 0.072448f
C2865 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.026506f
C2866 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.010335f
C2867 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.DONE 0.048717f
C2868 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.74594f
C2869 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_17730_30316# 0.01727f
C2870 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_28556# 0.135353f
C2871 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<5> 0.073518f
C2872 SUNSAR_SAR8B_CV_0.SARN a_12582_5094# 0.049641f
C2873 SUNSAR_SAR8B_CV_0.XA20.CPO a_13842_28204# 0.067146f
C2874 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N a_17730_28908# 0.060353f
C2875 SUNSAR_SAR8B_CV_0.XA20.CNO a_7650_27852# 0.074163f
C2876 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.029312f
C2877 SUNSAR_SAR8B_CV_0.SARP a_13950_4038# 0.025713f
C2878 SUNSAR_SAR8B_CV_0.D<2> a_15210_32956# 0.017466f
C2879 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S 0.044153f
C2880 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_3762_35948# 0.070424f
C2881 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.229239f
C2882 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S VPWR 0.097536f
C2883 a_16542_4566# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.011545f
C2884 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.CKN 0.41624f
C2885 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.016774f
C2886 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_34716# 0.077282f
C2887 a_11142_4038# ua[1] 0.043386f
C2888 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_2610_32076# 0.088002f
C2889 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA20.CPO 0.068386f
C2890 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S 0.050207f
C2891 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_17750_41880# 0.035868f
C2892 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<1> 0.180769f
C2893 uio_oe[3] uio_oe[2] 0.023797f
C2894 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43288# 0.03616f
C2895 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S 0.036094f
C2896 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA6.A 0.040072f
C2897 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S 0.030434f
C2898 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S 0.026188f
C2899 a_15230_40296# VPWR 0.457171f
C2900 tt_um_TT06_SAR_done_0.DONE a_5150_40296# 0.026182f
C2901 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.027044f
C2902 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B 6.86675f
C2903 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.074269f
C2904 a_20270_43816# VPWR 0.391817f
C2905 a_13862_43816# uo_out[3] 0.024759f
C2906 a_9990_5974# a_9990_5622# 0.010937f
C2907 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_11342_41880# 0.067588f
C2908 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S 0.089305f
C2909 a_13842_35420# a_13842_35068# 0.010937f
C2910 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_5150_41000# 0.156079f
C2911 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.ENO 0.051732f
C2912 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S 0.021211f
C2913 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.419738f
C2914 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2502_4688# 0.024512f
C2915 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.058243f
C2916 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.04064f
C2917 a_11342_42760# SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.071391f
C2918 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43816# 0.127669f
C2919 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.294852f
C2920 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_27852# 0.025674f
C2921 a_7670_41352# a_7670_41000# 0.010937f
C2922 a_16362_37180# SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.069366f
C2923 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA3.CEIN 0.033943f
C2924 a_6282_37180# a_6282_36828# 0.010937f
C2925 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S 0.050648f
C2926 a_20250_32076# VPWR 0.433941f
C2927 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S 0.027192f
C2928 SUNSAR_SAR8B_CV_0.XA0.XA9.B a_2610_35420# 0.017683f
C2929 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.527529f
C2930 a_20250_28204# VPWR 0.361706f
C2931 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> a_3762_33836# 0.011483f
C2932 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.071571f
C2933 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.CP0 0.08098f
C2934 SUNSAR_SAR8B_CV_0.XA6.CN1 a_18882_31196# 0.070763f
C2935 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.204048f
C2936 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_28556# 0.073834f
C2937 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_15390_5622# 0.03948f
C2938 a_10190_42408# VPWR 0.391292f
C2939 SUNSAR_SAR8B_CV_0.XA20.CPO a_12690_28204# 0.09022f
C2940 SUNSAR_SAR8B_CV_0.XA20.CNO a_6282_27852# 0.072592f
C2941 a_10170_36828# VPWR 0.396003f
C2942 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.301665f
C2943 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR 0.09699f
C2944 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_11322_27148# 0.023111f
C2945 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S a_10170_27852# 0.04865f
C2946 a_20250_28204# a_20250_27852# 0.010937f
C2947 SUNSAR_SAR8B_CV_0.SARP a_12582_4038# 0.016299f
C2948 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S 0.044228f
C2949 a_13842_36300# a_13842_35948# 0.010937f
C2950 SUNSAR_SAR8B_CV_0.XA0.XA10.A a_2610_35948# 0.132671f
C2951 SUNSAR_CAPT8B_CV_0.XE10.XA6.A uo_out[4] 0.014139f
C2952 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S VPWR 0.097536f
C2953 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR 0.035055f
C2954 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_9990_4038# 0.034677f
C2955 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S 0.101001f
C2956 SUNSAR_SAR8B_CV_0.XA7.EN a_17730_34716# 0.066245f
C2957 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 0.635098f
C2958 a_9990_4038# ua[1] 0.023111f
C2959 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA20.CNO 0.053965f
C2960 SUNSAR_SAR8B_CV_0.XA1.EN a_6282_29612# 0.073155f
C2961 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<1> 0.07415f
C2962 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.63636f
C2963 a_20270_43816# SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.071475f
C2964 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S 0.050207f
C2965 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S 0.010745f
C2966 a_13862_40296# VPWR 0.458821f
C2967 tt_um_TT06_SAR_done_0.DONE a_3782_40296# 0.026182f
C2968 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA2.CEIN 0.05126f
C2969 a_17730_28556# a_17730_28204# 0.010937f
C2970 a_20250_35068# VPWR 0.391458f
C2971 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.070556f
C2972 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.019775f
C2973 a_18902_43816# VPWR 0.391817f
C2974 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[0] 0.453892f
C2975 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR 0.104609f
C2976 SUNSAR_SAR8B_CV_0.XA3.XA9.B a_11322_34716# 0.047651f
C2977 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_10190_41880# 0.071088f
C2978 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.039903f
C2979 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_13862_41352# 0.058557f
C2980 SUNSAR_CAPT8B_CV_0.XA6.A a_23942_41880# 0.091053f
C2981 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_SAR8B_CV_0.D<0> 0.393578f
C2982 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S 0.021266f
C2983 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2358_4688# 0.049023f
C2984 a_5130_26796# VPWR 0.441753f
C2985 a_11322_33836# SUNSAR_SAR8B_CV_0.XA3.CP0 0.066219f
C2986 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.26537f
C2987 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.090222f
C2988 a_10190_42760# SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.067588f
C2989 a_2630_42760# a_2630_42408# 0.010937f
C2990 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.02398f
C2991 SUNSAR_SAR8B_CV_0.D<0> VPWR 5.69368f
C2992 a_12710_44168# a_12710_43816# 0.010937f
C2993 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S 0.050207f
C2994 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S 0.050207f
C2995 a_20250_35948# VPWR 0.414756f
C2996 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 6.86675f
C2997 a_5130_28908# a_5130_28556# 0.010937f
C2998 a_15210_37180# SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.067588f
C2999 a_16362_37180# SUNSAR_SAR8B_CV_0.XA6.CEIN 0.024074f
C3000 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.377598f
C3001 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.074964f
C3002 a_13842_27500# a_13842_27148# 0.010937f
C3003 a_18882_32076# VPWR 0.436368f
C3004 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA20.CPO 0.074065f
C3005 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.DONE 0.049573f
C3006 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S 0.023798f
C3007 a_18882_28204# VPWR 0.36179f
C3008 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.085036f
C3009 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C3010 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C3011 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.748719f
C3012 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S 0.013533f
C3013 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_16362_30316# 0.01727f
C3014 a_8822_42408# VPWR 0.391292f
C3015 SUNSAR_SAR8B_CV_0.XA20.CPO a_11322_28204# 0.088673f
C3016 SUNSAR_SAR8B_CV_0.XA20.CNO a_5130_27852# 0.067588f
C3017 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S 0.050207f
C3018 a_8802_36828# VPWR 0.396052f
C3019 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR 0.405511f
C3020 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_10170_27148# 0.03422f
C3021 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_20250_27500# 0.033843f
C3022 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.038188f
C3023 SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR 1.63909f
C3024 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR 0.035055f
C3025 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.011708f
C3026 SUNSAR_SAR8B_CV_0.XA5.XA9.B a_15210_33836# 0.023316f
C3027 a_9990_3334# VPWR 0.380282f
C3028 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.175642f
C3029 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA20.CNO 0.053594f
C3030 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.310451f
C3031 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_16382_41880# 0.035868f
C3032 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_SAR8B_CV_0.D<0> 0.018133f
C3033 uio_oe[4] uio_oe[3] 0.023797f
C3034 uo_out[0] uio_in[7] 0.030841f
C3035 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S 0.024389f
C3036 a_23942_40648# ui_in[0] 0.068184f
C3037 SUNSAR_CAPT8B_CV_0.XG12.QN a_16382_43288# 0.03616f
C3038 tt_um_TT06_SAR_done_0.DONE a_2630_40296# 0.042653f
C3039 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S a_5130_28204# 0.04865f
C3040 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_6282_28204# 0.067588f
C3041 a_18882_35068# VPWR 0.394528f
C3042 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.010335f
C3043 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.08276f
C3044 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S 0.016767f
C3045 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.232115f
C3046 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[1] 0.238239f
C3047 SUNSAR_SAR8B_CV_0.XA3.XA9.B a_10170_34716# 0.023982f
C3048 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_41352# 0.060327f
C3049 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_13862_41352# 0.075505f
C3050 SUNSAR_CAPT8B_CV_0.XA6.A a_22790_41880# 0.111538f
C3051 a_12690_35420# a_12690_35068# 0.010937f
C3052 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.SARP 0.050902f
C3053 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_SAR8B_CV_0.D<0> 0.241356f
C3054 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN 0.144331f
C3055 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.419738f
C3056 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_4848# 0.105547f
C3057 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.058243f
C3058 a_3762_26796# VPWR 0.442908f
C3059 a_10170_33836# SUNSAR_SAR8B_CV_0.XA3.CP0 0.067588f
C3060 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.268769f
C3061 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.058755f
C3062 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.041437f
C3063 SUNSAR_CAPT8B_CV_0.XA7.MP0.G SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.031791f
C3064 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S VPWR 0.106927f
C3065 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.029914f
C3066 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.383512f
C3067 a_6302_41352# a_6302_41000# 0.010937f
C3068 SUNSAR_SAR8B_CV_0.D<3> tt_um_TT06_SAR_done_0.DONE 0.295397f
C3069 a_18882_35948# VPWR 0.417826f
C3070 a_15210_37180# SUNSAR_SAR8B_CV_0.XA6.CEIN 0.029627f
C3071 a_5130_37180# a_5130_36828# 0.010937f
C3072 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23922_34540# 0.017541f
C3073 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.073805f
C3074 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.134182f
C3075 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.038658f
C3076 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_6302_42760# 0.091344f
C3077 SUNSAR_SAR8B_CV_0.XA20.XA12.Y a_23922_35420# 0.098978f
C3078 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.SARN 0.041877f
C3079 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.CP0 0.08098f
C3080 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_28556# 0.075865f
C3081 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.SARP 0.032416f
C3082 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.D<6> 0.075797f
C3083 SUNSAR_SAR8B_CV_0.XA20.CPO a_10170_28204# 0.068716f
C3084 SUNSAR_SAR8B_CV_0.XA20.CNO a_3762_27852# 0.066018f
C3085 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.CEIN 0.03012f
C3086 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR 1.70987f
C3087 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S a_8802_27852# 0.04865f
C3088 a_18882_28204# a_18882_27852# 0.010937f
C3089 a_12690_36300# a_12690_35948# 0.010937f
C3090 a_23922_36300# SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.034234f
C3091 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_34716# 0.067815f
C3092 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.42639f
C3093 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.010925f
C3094 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.012886f
C3095 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA20.CNO 0.054464f
C3096 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.082663f
C3097 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.058669f
C3098 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.15234f
C3099 SUNSAR_CAPT8B_CV_0.XG12.XA5.A a_15230_41880# 0.024901f
C3100 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<2> 0.18141f
C3101 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S 0.050207f
C3102 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S 0.030434f
C3103 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S 0.026257f
C3104 a_22790_40648# ui_in[0] 0.076643f
C3105 SUNSAR_CAPT8B_CV_0.XG12.QN a_15230_43288# 0.024901f
C3106 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.CEIN 0.075193f
C3107 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S 0.073693f
C3108 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_5130_28204# 0.096735f
C3109 a_16362_28556# a_16362_28204# 0.010937f
C3110 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW uio_out[0] 0.088825f
C3111 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR 0.042839f
C3112 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_12710_41352# 0.080002f
C3113 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S 0.036491f
C3114 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9054_4848# 0.0666f
C3115 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.090222f
C3116 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.239611f
C3117 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_15230_42408# 0.015723f
C3118 a_8822_42760# SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.066018f
C3119 SUNSAR_CAPT8B_CV_0.XA7.MP0.G a_23942_43992# 0.073828f
C3120 a_11342_44168# a_11342_43816# 0.010937f
C3121 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_27852# 0.010898f
C3122 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S 0.011062f
C3123 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S VPWR 0.106927f
C3124 a_3762_28908# a_3762_28556# 0.010937f
C3125 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.293159f
C3126 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.DONE 0.02194f
C3127 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22770_34540# 0.012281f
C3128 a_12690_27500# a_12690_27148# 0.010937f
C3129 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.2165f
C3130 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.026506f
C3131 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S 0.027192f
C3132 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_5150_42760# 0.111734f
C3133 a_23922_35948# SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.023111f
C3134 SUNSAR_SAR8B_CV_0.XA20.XA12.Y a_22770_35420# 0.067834f
C3135 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.DONE 0.048717f
C3136 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.165965f
C3137 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA3a.A 0.136678f
C3138 SUNSAR_SAR8B_CV_0.XA3.EN a_7650_28556# 0.132757f
C3139 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C3140 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28908# 0.066932f
C3141 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G 0.08427f
C3142 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.138433f
C3143 SUNSAR_SAR8B_CV_0.XA20.CPO a_8802_28204# 0.067146f
C3144 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N a_16362_28908# 0.060353f
C3145 SUNSAR_SAR8B_CV_0.XA20.CNO a_2610_27852# 0.074097f
C3146 a_28727_40307# a_28727_39955# 0.010937f
C3147 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.029317f
C3148 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR 0.097407f
C3149 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.228208f
C3150 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S 0.03516f
C3151 SUNSAR_SAR8B_CV_0.D<3> a_13842_32956# 0.017466f
C3152 a_22770_36300# SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.023111f
C3153 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XB1.CKN 0.143148f
C3154 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR 0.104609f
C3155 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_34716# 0.075712f
C3156 SUNSAR_SAR8B_CV_0.EN a_20250_27148# 0.066018f
C3157 a_13950_4390# ua[0] 0.05387f
C3158 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.036102f
C3159 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.340491f
C3160 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<2> 0.074634f
C3161 uio_oe[5] uio_oe[4] 0.023797f
C3162 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S 0.026117f
C3163 a_10190_40296# VPWR 0.457269f
C3164 a_23942_41000# a_23942_40648# 0.010937f
C3165 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 27.1615f
C3166 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.725407f
C3167 a_15230_43816# VPWR 0.391817f
C3168 a_10190_43816# uo_out[4] 0.022673f
C3169 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW uio_oe[0] 0.135493f
C3170 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR 0.042839f
C3171 a_11322_35420# a_11322_35068# 0.010937f
C3172 a_22770_35420# SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.031543f
C3173 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA7.EN 0.051732f
C3174 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2502_5648# 0.024512f
C3175 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.046398f
C3176 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.031784f
C3177 a_23922_27148# VPWR 0.483246f
C3178 SUNSAR_SAR8B_CV_0.SARN a_22770_33132# 0.022743f
C3179 a_8802_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.066018f
C3180 a_7670_42760# SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.072962f
C3181 SUNSAR_CAPT8B_CV_0.XA7.MP0.G a_22790_43992# 0.066018f
C3182 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_27852# 0.024578f
C3183 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP 0.435464f
C3184 SUNSAR_SAR8B_CV_0.D<1> VPWR 5.47059f
C3185 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S 0.062799f
C3186 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S 0.050207f
C3187 a_5150_41352# a_5150_41000# 0.010937f
C3188 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.252966f
C3189 a_3762_37180# a_3762_36828# 0.010937f
C3190 a_13842_37180# SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.066018f
C3191 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA2.CEIN 0.432008f
C3192 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S 0.031338f
C3193 a_15210_32076# VPWR 0.436368f
C3194 SUNSAR_CAPT8B_CV_0.XG12.XA7.C a_15230_42408# 0.076129f
C3195 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_16382_42408# 0.098561f
C3196 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S 0.030434f
C3197 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA20.CPO 0.074326f
C3198 a_15210_28204# VPWR 0.361706f
C3199 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.069846f
C3200 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.CP0 0.08098f
C3201 SUNSAR_SAR8B_CV_0.XA5.CN1 a_15210_31196# 0.069193f
C3202 a_5150_42408# VPWR 0.391292f
C3203 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_28908# 0.073535f
C3204 SUNSAR_SAR8B_CV_0.XB2.TIE_L a_11142_5622# 0.03948f
C3205 SUNSAR_SAR8B_CV_0.XA20.CPO a_7650_28204# 0.09022f
C3206 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N a_15210_28908# 0.023475f
C3207 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S 0.064851f
C3208 a_5130_36828# VPWR 0.395767f
C3209 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_8802_27148# 0.03422f
C3210 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_18882_27500# 0.033843f
C3211 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S a_7650_27852# 0.056787f
C3212 a_17730_28204# a_17730_27852# 0.010937f
C3213 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.038188f
C3214 a_11322_36300# a_11322_35948# 0.010937f
C3215 SUNSAR_CAPT8B_CV_0.XD09.XA6.A uo_out[5] 0.014139f
C3216 SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR 1.63909f
C3217 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.017546f
C3218 a_21402_35068# a_21402_34716# 0.010937f
C3219 SUNSAR_SAR8B_CV_0.EN a_18882_27148# 0.067588f
C3220 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR 1.50074f
C3221 a_21402_32956# SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.066679f
C3222 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S 0.010423f
C3223 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_13862_41880# 0.024901f
C3224 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.233892f
C3225 a_18902_43816# SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 0.069905f
C3226 SUNSAR_CAPT8B_CV_0.XF11.QN a_13862_43288# 0.024901f
C3227 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S 0.027953f
C3228 a_8822_40296# VPWR 0.458821f
C3229 tt_um_TT06_SAR_done_0.DONE a_21422_40648# 0.08452f
C3230 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.025287f
C3231 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S a_3762_28204# 0.04865f
C3232 a_15210_28556# a_15210_28204# 0.010937f
C3233 a_15210_35068# VPWR 0.394528f
C3234 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.071417f
C3235 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.099137f
C3236 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.010854f
C3237 a_13862_43816# VPWR 0.391817f
C3238 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW clk 0.044089f
C3239 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N VPWR 0.271482f
C3240 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.SARP 0.102632f
C3241 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_8822_41880# 0.072658f
C3242 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2358_5648# 0.049023f
C3243 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.095491f
C3244 a_7650_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.067789f
C3245 a_10190_44168# a_10190_43816# 0.010937f
C3246 SUNSAR_SAR8B_CV_0.D<4> tt_um_TT06_SAR_done_0.DONE 0.295493f
C3247 a_2610_28908# a_2610_28556# 0.010937f
C3248 a_15210_35948# VPWR 0.417826f
C3249 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B 27.1632f
C3250 a_12690_37180# SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.070936f
C3251 a_13842_37180# SUNSAR_SAR8B_CV_0.XA5.CEIN 0.040807f
C3252 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.158152f
C3253 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S 0.053284f
C3254 a_11322_27500# a_11322_27148# 0.010937f
C3255 a_13842_32076# VPWR 0.436368f
C3256 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_42408# 0.031125f
C3257 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S 0.010335f
C3258 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.046858f
C3259 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S 0.027192f
C3260 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.DONE 0.049573f
C3261 a_13842_28204# VPWR 0.36179f
C3262 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S 0.028026f
C3263 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_12690_30316# 0.01727f
C3264 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.SARP 0.032416f
C3265 a_3782_42408# VPWR 0.391292f
C3266 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_28556# 0.135353f
C3267 SUNSAR_SAR8B_CV_0.XA20.CPO a_6282_28204# 0.088673f
C3268 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S 0.050207f
C3269 a_3762_36828# VPWR 0.395857f
C3270 a_27575_40307# a_27575_39955# 0.010937f
C3271 tt_um_TT06_SAR_done_0.x3.MP1.G a_28727_39955# 0.021508f
C3272 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR 4.36142f
C3273 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_7650_27148# 0.023111f
C3274 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S 0.016689f
C3275 a_21402_36300# SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.066704f
C3276 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S VPWR 0.097536f
C3277 SUNSAR_CAPT8B_CV_0.XA6.A clk 0.206733f
C3278 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.CKN 0.200119f
C3279 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_34716# 0.077282f
C3280 SUNSAR_SAR8B_CV_0.XA4.XA9.B a_13842_33836# 0.023316f
C3281 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR 0.183853f
C3282 a_12582_4390# ua[1] 0.05387f
C3283 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.437693f
C3284 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.SARP 0.506551f
C3285 a_20250_32956# SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.067588f
C3286 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<3> 0.180769f
C3287 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_12710_41880# 0.035868f
C3288 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S 0.036094f
C3289 uio_oe[0] uio_out[7] 0.03074f
C3290 SUNSAR_CAPT8B_CV_0.XF11.QN a_12710_43288# 0.03616f
C3291 uio_oe[6] uio_oe[5] 0.023797f
C3292 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S 0.030434f
C3293 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.010898f
C3294 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N a_7650_29612# 0.031412f
C3295 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S 0.0111f
C3296 a_22790_41000# a_22790_40648# 0.010937f
C3297 tt_um_TT06_SAR_done_0.DONE a_20270_40648# 0.066617f
C3298 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_3762_28204# 0.098305f
C3299 a_13842_35068# VPWR 0.394528f
C3300 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.010335f
C3301 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S 0.028452f
C3302 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ui_in[0] 0.097118f
C3303 SUNSAR_CAPT8B_CV_0.XI14.QN uio_out[0] 0.021018f
C3304 a_8822_43816# uo_out[5] 0.022673f
C3305 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_3782_41000# 0.15757f
C3306 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_7670_41880# 0.066018f
C3307 SUNSAR_SAR8B_CV_0.XA2.XA9.B a_8802_34716# 0.023982f
C3308 a_10170_35420# a_10170_35068# 0.010937f
C3309 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_5808# 0.105547f
C3310 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.046398f
C3311 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.031784f
C3312 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S a_23922_33132# 0.023111f
C3313 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.036726f
C3314 a_6302_42760# SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.071391f
C3315 a_21422_44168# SUNSAR_CAPT8B_CV_0.XI14.QN 0.069523f
C3316 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S 0.050207f
C3317 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S 0.062799f
C3318 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.276413f
C3319 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_27852# 0.025674f
C3320 a_3782_41352# a_3782_41000# 0.010937f
C3321 a_13842_35948# VPWR 0.417826f
C3322 a_2610_37180# a_2610_36828# 0.010937f
C3323 a_12690_37180# SUNSAR_SAR8B_CV_0.XA5.CEIN 0.023111f
C3324 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S 0.022628f
C3325 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A 0.011542f
C3326 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S 0.023798f
C3327 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.038846f
C3328 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S 0.027192f
C3329 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.CP0 0.08098f
C3330 SUNSAR_SAR8B_CV_0.XA4.CN1 a_13842_31196# 0.070763f
C3331 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_28908# 0.072087f
C3332 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_28556# 0.073834f
C3333 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<7> 0.010193f
C3334 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S 0.030434f
C3335 SUNSAR_SAR8B_CV_0.XA20.CPO a_5130_28204# 0.068716f
C3336 tt_um_TT06_SAR_done_0.x3.MP1.G a_27575_39955# 0.034104f
C3337 a_23922_34540# VPWR 0.502044f
C3338 a_16362_28204# a_16362_27852# 0.010937f
C3339 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S a_6282_27852# 0.056787f
C3340 SUNSAR_SAR8B_CV_0.SARP a_13950_4390# 0.039425f
C3341 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S 0.016683f
C3342 a_10170_36300# a_10170_35948# 0.010937f
C3343 a_20250_36300# SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.067588f
C3344 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S VPWR 0.097536f
C3345 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR 0.104609f
C3346 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.101001f
C3347 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S 0.011382f
C3348 SUNSAR_SAR8B_CV_0.XA5.EN a_12690_34716# 0.066245f
C3349 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.010925f
C3350 a_20250_35068# a_20250_34716# 0.010937f
C3351 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VPWR 1.50269f
C3352 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.082663f
C3353 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<3> 0.07415f
C3354 a_17750_43816# SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.073123f
C3355 uio_oe[0] uio_oe[1] 0.023797f
C3356 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S 0.025128f
C3357 tt_um_TT06_SAR_done_0.DONE a_18902_40648# 0.068187f
C3358 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S 0.073693f
C3359 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_2610_28204# 0.066018f
C3360 a_13842_28556# a_13842_28204# 0.010937f
C3361 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.019775f
C3362 SUNSAR_SAR8B_CV_0.D<0> a_20250_34716# 0.070775f
C3363 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.074602f
C3364 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR 0.104609f
C3365 SUNSAR_CAPT8B_CV_0.XH13.QN uio_out[0] 0.021018f
C3366 SUNSAR_CAPT8B_CV_0.XI14.QN uio_oe[0] 0.032f
C3367 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_2630_41000# 0.114097f
C3368 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S 0.036491f
C3369 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_11342_41352# 0.078431f
C3370 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW tt_um_TT06_SAR_done_0.DONE 0.094851f
C3371 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN 0.144331f
C3372 SUNSAR_SAR8B_CV_0.XA2.XA9.B a_7650_34716# 0.047651f
C3373 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_21402_35068# 0.129098f
C3374 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9054_5808# 0.0666f
C3375 a_20250_27148# VPWR 0.470364f
C3376 a_6282_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.066219f
C3377 a_5150_42760# SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.067588f
C3378 a_8822_44168# a_8822_43816# 0.010937f
C3379 a_20270_44168# SUNSAR_CAPT8B_CV_0.XI14.QN 0.067588f
C3380 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_21402_29612# 0.040867f
C3381 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S 0.041902f
C3382 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S 0.011178f
C3383 SUNSAR_SAR8B_CV_0.D<2> VPWR 5.45923f
C3384 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.CEIN 0.075291f
C3385 a_10170_27500# a_10170_27148# 0.010937f
C3386 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.86675f
C3387 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_3782_42760# 0.113305f
C3388 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.527529f
C3389 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA20.CPO 0.075237f
C3390 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.048717f
C3391 a_16542_2982# a_16542_2630# 0.010937f
C3392 SUNSAR_SAR8B_CV_0.XA4.CN1 a_12690_31196# 0.107567f
C3393 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR 0.686731f
C3394 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_11322_30316# 0.01727f
C3395 SUNSAR_SAR8B_CV_0.XA7.EN a_17730_28908# 0.068502f
C3396 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S 0.055627f
C3397 SUNSAR_SAR8B_CV_0.XA20.CPO a_3762_28204# 0.067146f
C3398 SUNSAR_SAR8B_CV_0.XA7.XA12.A VPWR 0.714341f
C3399 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.064851f
C3400 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.022538f
C3401 tt_um_TT06_SAR_done_0.x3.MP1.G a_28727_40307# 0.070033f
C3402 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.021955f
C3403 a_22770_34540# VPWR 0.024886f
C3404 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CP0 0.320252f
C3405 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S 0.03516f
C3406 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.638363f
C3407 a_16542_4566# SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.071041f
C3408 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.CKN 0.41624f
C3409 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.018669f
C3410 SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR 1.63909f
C3411 SUNSAR_SAR8B_CV_0.EN a_15210_27148# 0.066018f
C3412 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S 0.026506f
C3413 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR 0.183853f
C3414 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.175642f
C3415 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA20.CPO 0.068426f
C3416 a_18882_32956# SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.066018f
C3417 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_SAR8B_CV_0.D<1> 0.018133f
C3418 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_11342_41880# 0.035868f
C3419 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S 0.024386f
C3420 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43288# 0.03616f
C3421 uio_oe[7] uio_oe[6] 0.023797f
C3422 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S 0.050207f
C3423 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S 0.026188f
C3424 a_5150_40296# VPWR 0.457199f
C3425 a_21422_41000# a_21422_40648# 0.010937f
C3426 tt_um_TT06_SAR_done_0.DONE a_17750_40648# 0.083091f
C3427 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6519f
C3428 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.085086f
C3429 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.070567f
C3430 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N VPWR 0.271482f
C3431 a_10190_43816# VPWR 0.391817f
C3432 SUNSAR_CAPT8B_CV_0.XG12.QN uio_out[0] 0.021018f
C3433 SUNSAR_CAPT8B_CV_0.XH13.QN uio_oe[0] 0.032f
C3434 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_SAR8B_CV_0.D<1> 0.241356f
C3435 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_10190_41352# 0.077076f
C3436 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_11342_41352# 0.060327f
C3437 SUNSAR_SAR8B_CV_0.XA7.XA9.B a_21402_35068# 0.011912f
C3438 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_20250_35068# 0.089492f
C3439 a_18882_35420# SUNSAR_SAR8B_CV_0.XA6.DONE 0.023111f
C3440 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA6.EN 0.051732f
C3441 a_8802_35420# a_8802_35068# 0.010937f
C3442 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.SARP 0.081546f
C3443 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2502_6608# 0.024512f
C3444 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.449584f
C3445 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B 0.014291f
C3446 a_18882_27148# VPWR 0.471462f
C3447 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.386137f
C3448 a_5130_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.067588f
C3449 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_20250_29612# 0.023777f
C3450 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S 0.152518f
C3451 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S 0.041456f
C3452 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S VPWR 0.106927f
C3453 SUNSAR_SAR8B_CV_0.D<5> tt_um_TT06_SAR_done_0.DONE 0.295822f
C3454 a_2630_41352# a_2630_41000# 0.010937f
C3455 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.018236f
C3456 a_11322_37180# SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.069366f
C3457 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.030459f
C3458 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.050524f
C3459 a_10170_32076# VPWR 0.436368f
C3460 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.12241f
C3461 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_2630_42760# 0.089774f
C3462 a_21402_35948# SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.071154f
C3463 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S 0.027192f
C3464 a_10170_28204# VPWR 0.361706f
C3465 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.092293f
C3466 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.110078f
C3467 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR 0.898003f
C3468 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_28556# 0.075865f
C3469 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S 0.026885f
C3470 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S 0.030434f
C3471 SUNSAR_SAR8B_CV_0.XA20.CPO a_2610_28204# 0.09022f
C3472 SUNSAR_SAR8B_CV_0.XA20.CK_CMP VPWR 1.1111f
C3473 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.064851f
C3474 tt_um_TT06_SAR_done_0.x3.MP1.G a_27575_40307# 0.099188f
C3475 a_28727_40659# a_28727_40307# 0.010937f
C3476 a_15210_28204# a_15210_27852# 0.010937f
C3477 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S a_5130_27852# 0.04865f
C3478 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_6282_27148# 0.023111f
C3479 a_18882_36300# SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.066018f
C3480 a_8802_36300# a_8802_35948# 0.010937f
C3481 SUNSAR_CAPT8B_CV_0.XC08.XA6.A uo_out[6] 0.014938f
C3482 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR 0.035055f
C3483 a_21422_43288# uo_out[0] 0.067687f
C3484 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.250503f
C3485 a_15390_4566# SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.036098f
C3486 a_13950_4742# a_13950_4390# 0.010937f
C3487 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.CKN 0.015687f
C3488 SUNSAR_SAR8B_CV_0.EN a_13842_27148# 0.067588f
C3489 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_34716# 0.067815f
C3490 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S 0.055045f
C3491 a_18882_35068# a_18882_34716# 0.010937f
C3492 a_16542_4038# VPWR 0.379979f
C3493 SUNSAR_SAR8B_CV_0.XB2.XA4.GN ua[0] 0.765539f
C3494 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.437693f
C3495 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.116333f
C3496 a_17730_32956# SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.06825f
C3497 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<4> 0.18141f
C3498 SUNSAR_CAPT8B_CV_0.XE10.XA5.A a_10190_41880# 0.024901f
C3499 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.63636f
C3500 SUNSAR_CAPT8B_CV_0.XE10.QN a_10190_43288# 0.024901f
C3501 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 a_23922_28556# 0.023111f
C3502 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S 0.010745f
C3503 a_3782_40296# VPWR 0.458821f
C3504 tt_um_TT06_SAR_done_0.DONE a_16382_40648# 0.084662f
C3505 a_10170_35068# VPWR 0.394528f
C3506 a_12690_28556# a_12690_28204# 0.010937f
C3507 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.010772f
C3508 SUNSAR_CAPT8B_CV_0.XG12.QN uio_oe[0] 0.031059f
C3509 a_8822_43816# VPWR 0.391817f
C3510 SUNSAR_CAPT8B_CV_0.XF11.QN uio_out[0] 0.021018f
C3511 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_SAR8B_CV_0.D<1> 0.393049f
C3512 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S 0.021266f
C3513 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_41352# 0.058557f
C3514 a_17730_35420# SUNSAR_SAR8B_CV_0.XA6.DONE 0.030547f
C3515 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_2358_6608# 0.049023f
C3516 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 0.671839f
C3517 a_3782_42760# SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.066018f
C3518 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.301485f
C3519 a_7670_44168# a_7670_43816# 0.010937f
C3520 a_18902_44168# SUNSAR_CAPT8B_CV_0.XH13.QN 0.066018f
C3521 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.375025f
C3522 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S 0.050207f
C3523 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S VPWR 0.106927f
C3524 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_27852# 0.010898f
C3525 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.284482f
C3526 a_10170_35948# VPWR 0.417826f
C3527 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 13.652401f
C3528 a_10170_37180# SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.067588f
C3529 a_11322_37180# SUNSAR_SAR8B_CV_0.XA4.CEIN 0.024074f
C3530 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.098006f
C3531 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.075315f
C3532 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.078716f
C3533 a_8802_27500# a_8802_27148# 0.010937f
C3534 a_8802_32076# VPWR 0.436368f
C3535 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.432466f
C3536 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_13862_42408# 0.031125f
C3537 a_20250_35948# SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.067588f
C3538 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.049573f
C3539 a_8802_28204# VPWR 0.36179f
C3540 a_15390_2982# a_15390_2630# 0.010937f
C3541 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_28908# 0.06753f
C3542 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.CPO 0.131536f
C3543 SUNSAR_SAR8B_CV_0.XA3.CN1 a_11322_31196# 0.109137f
C3544 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR 0.898003f
C3545 SUNSAR_SAR8B_CV_0.XA1.EN a_2610_28556# 0.132757f
C3546 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA6.A 0.011748f
C3547 SUNSAR_SAR8B_CV_0.XA6.XA12.A VPWR 0.723713f
C3548 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S 0.050207f
C3549 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_15210_27500# 0.033843f
C3550 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_5130_27148# 0.03422f
C3551 SUNSAR_SAR8B_CV_0.D<4> a_10170_32956# 0.017466f
C3552 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S 0.044153f
C3553 a_17730_36300# SUNSAR_SAR8B_CV_0.XA6.XA10.A 0.068275f
C3554 a_20270_43288# uo_out[0] 0.071088f
C3555 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.017476f
C3556 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR 0.035055f
C3557 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_34716# 0.075712f
C3558 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.014021f
C3559 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.014291f
C3560 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.065837f
C3561 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.143633f
C3562 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.152052f
C3563 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<4> 0.074691f
C3564 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.B 0.012998f
C3565 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.010898f
C3566 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N a_6282_29612# 0.031412f
C3567 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S 0.024389f
C3568 a_20270_41000# a_20270_40648# 0.010937f
C3569 tt_um_TT06_SAR_done_0.DONE a_15230_40648# 0.066617f
C3570 a_8802_35068# VPWR 0.394528f
C3571 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.075181f
C3572 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S 0.028448f
C3573 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.010335f
C3574 SUNSAR_CAPT8B_CV_0.XI14.QN uo_out[0] 0.24816f
C3575 SUNSAR_CAPT8B_CV_0.XF11.QN uio_oe[0] 0.018103f
C3576 a_5150_43816# uo_out[6] 0.022673f
C3577 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S 0.021211f
C3578 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_6302_41880# 0.067588f
C3579 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN 0.144331f
C3580 a_7650_35420# a_7650_35068# 0.010937f
C3581 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_6768# 0.105547f
C3582 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.449584f
C3583 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 0.014291f
C3584 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.034649f
C3585 a_3762_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.066018f
C3586 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.035717f
C3587 a_2630_42760# SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.072962f
C3588 a_17750_44168# SUNSAR_CAPT8B_CV_0.XH13.QN 0.071093f
C3589 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_18882_29612# 0.023777f
C3590 SUNSAR_SAR8B_CV_0.D<3> VPWR 5.44876f
C3591 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S 0.150467f
C3592 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_27852# 0.024578f
C3593 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.019052f
C3594 a_8802_35948# VPWR 0.417826f
C3595 a_10170_37180# SUNSAR_SAR8B_CV_0.XA4.CEIN 0.029627f
C3596 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S 0.022425f
C3597 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.07371f
C3598 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S 0.030434f
C3599 SUNSAR_CAPT8B_CV_0.XF11.XA7.C a_13862_42408# 0.074559f
C3600 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_42408# 0.100131f
C3601 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.038658f
C3602 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA20.CPO 0.067023f
C3603 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.168325f
C3604 SUNSAR_SAR8B_CV_0.XA6.EN a_15210_28908# 0.073535f
C3605 SUNSAR_SAR8B_CV_0.XA3.CN1 a_10170_31196# 0.069193f
C3606 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR 0.898003f
C3607 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.A 0.504864f
C3608 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S 0.010682f
C3609 SUNSAR_SAR8B_CV_0.XA7.CEIN VPWR 2.28789f
C3610 a_28727_40659# tt_um_TT06_SAR_done_0.x3.MP1.G 0.065834f
C3611 a_27575_40659# a_27575_40307# 0.010937f
C3612 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 1.62434f
C3613 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR 0.097407f
C3614 a_13842_28204# a_13842_27852# 0.010937f
C3615 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S a_3762_27852# 0.04865f
C3616 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.01255f
C3617 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S 0.044297f
C3618 a_7650_36300# a_7650_35948# 0.010937f
C3619 SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR 1.63909f
C3620 a_9990_4566# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.011545f
C3621 a_12582_4742# a_12582_4390# 0.010937f
C3622 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.010925f
C3623 a_17730_35068# a_17730_34716# 0.010937f
C3624 a_23922_34892# SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.023111f
C3625 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.CN0 0.093524f
C3626 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.144751f
C3627 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.181018f
C3628 a_16362_32956# SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.066679f
C3629 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA20.CPO 0.068386f
C3630 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.339883f
C3631 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.054448f
C3632 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_8822_41880# 0.024901f
C3633 SUNSAR_CAPT8B_CV_0.XD09.QN a_8822_43288# 0.024901f
C3634 a_16382_43816# SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.071553f
C3635 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S 0.026257f
C3636 a_23942_40648# VPWR 0.490244f
C3637 tt_um_TT06_SAR_done_0.DONE a_13862_40648# 0.068187f
C3638 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S 0.073693f
C3639 a_11322_28556# a_11322_28204# 0.010937f
C3640 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.077963f
C3641 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.06386f
C3642 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S 0.016769f
C3643 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.010502f
C3644 SUNSAR_SAR8B_CV_0.D<1> a_18882_34716# 0.069204f
C3645 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR 0.104609f
C3646 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_5150_41880# 0.071088f
C3647 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_18882_35068# 0.091063f
C3648 a_16362_35420# SUNSAR_SAR8B_CV_0.XA5.DONE 0.031235f
C3649 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARP 0.187721f
C3650 SUNSAR_SAR8B_CV_0.XA1.XA9.B a_6282_34716# 0.047651f
C3651 a_15210_27148# VPWR 0.470364f
C3652 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9054_6768# 0.0666f
C3653 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_23922_31724# 0.067588f
C3654 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.CPO 0.372599f
C3655 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.034649f
C3656 a_2610_33836# SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.067789f
C3657 a_6302_44168# a_6302_43816# 0.010937f
C3658 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S 0.050207f
C3659 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S 0.050207f
C3660 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_17730_29612# 0.040867f
C3661 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.040976f
C3662 SUNSAR_SAR8B_CV_0.D<6> tt_um_TT06_SAR_done_0.DONE 0.2961f
C3663 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S 0.050648f
C3664 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1615f
C3665 a_7650_27500# a_7650_27148# 0.010937f
C3666 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.026506f
C3667 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.105906f
C3668 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.010335f
C3669 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S 0.027192f
C3670 a_13950_2982# a_13950_2630# 0.010937f
C3671 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.059183f
C3672 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.067025f
C3673 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 3.45828f
C3674 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C3675 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR 0.898003f
C3676 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 a_22770_30844# 0.030757f
C3677 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_7650_30316# 0.01727f
C3678 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.033659f
C3679 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.143023f
C3680 SUNSAR_SAR8B_CV_0.XA5.XA12.A VPWR 0.720096f
C3681 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S 0.050207f
C3682 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.064851f
C3683 a_27575_40659# tt_um_TT06_SAR_done_0.x3.MP1.G 0.070359f
C3684 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR 0.112098f
C3685 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.020332f
C3686 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.37807f
C3687 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CP0 0.31626f
C3688 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.EN 0.227503f
C3689 a_16362_36300# SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.066704f
C3690 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S VPWR 0.097536f
C3691 a_18902_43288# uo_out[1] 0.072658f
C3692 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR 0.104609f
C3693 SUNSAR_SAR8B_CV_0.XA3.XA9.B a_10170_33836# 0.023316f
C3694 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_34716# 0.077282f
C3695 SUNSAR_SAR8B_CV_0.EN a_10170_27148# 0.066018f
C3696 a_22770_34892# SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.036577f
C3697 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.139425f
C3698 a_15210_32956# SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.067588f
C3699 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.B 0.297144f
C3700 SUNSAR_CAPT8B_CV_0.XD09.XA5.A a_7670_41880# 0.035868f
C3701 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<5> 0.180769f
C3702 ua[1] ua[0] 3.85017f
C3703 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43288# 0.03616f
C3704 a_23942_43992# a_23942_43640# 0.010937f
C3705 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S 0.050207f
C3706 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S 0.026117f
C3707 a_18902_41000# a_18902_40648# 0.010937f
C3708 tt_um_TT06_SAR_done_0.DONE a_12710_40648# 0.083091f
C3709 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA12.Y 0.151003f
C3710 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.55251f
C3711 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.300886f
C3712 SUNSAR_CAPT8B_CV_0.XH13.QN uo_out[1] 0.248827f
C3713 a_5150_43816# VPWR 0.391817f
C3714 a_3782_43816# uo_out[7] 0.02434f
C3715 SUNSAR_SAR8B_CV_0.XA6.XA9.A a_17730_35068# 0.127528f
C3716 a_15210_35420# SUNSAR_SAR8B_CV_0.XA5.DONE 0.023111f
C3717 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA5.EN 0.051732f
C3718 SUNSAR_SAR8B_CV_0.XA1.XA9.B a_5130_34716# 0.023982f
C3719 a_6282_35420# a_6282_35068# 0.010937f
C3720 a_13842_27148# VPWR 0.471462f
C3721 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.011022f
C3722 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.026917f
C3723 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.107427f
C3724 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_22770_31724# 0.071657f
C3725 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.034649f
C3726 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23942_42760# 0.101843f
C3727 a_16382_44168# SUNSAR_CAPT8B_CV_0.XG12.QN 0.069523f
C3728 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S 0.062799f
C3729 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.030034f
C3730 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_27852# 0.025674f
C3731 SUNSAR_CAPT8B_CV_0.XA4.MP1.G a_23942_41352# 0.023111f
C3732 a_8802_37180# SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.066018f
C3733 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.074964f
C3734 a_5130_32076# VPWR 0.436368f
C3735 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.527529f
C3736 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_SAR8B_CV_0.EN 0.03206f
C3737 a_5130_28204# VPWR 0.361706f
C3738 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.110246f
C3739 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S 0.028026f
C3740 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.033149f
C3741 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.SARP 0.032416f
C3742 SUNSAR_SAR8B_CV_0.XA5.EN a_13842_28908# 0.072087f
C3743 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR 0.898003f
C3744 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_8802_31196# 0.070763f
C3745 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S 0.026885f
C3746 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S 0.010682f
C3747 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N a_13842_28908# 0.023475f
C3748 SUNSAR_SAR8B_CV_0.XA6.CEIN VPWR 1.06023f
C3749 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.064851f
C3750 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.268016f
C3751 tt_um_TT06_SAR_done_0.x4.MP0.G tt_um_TT06_SAR_done_0.x3.MP1.G 0.071481f
C3752 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR 0.112858f
C3753 a_12690_28204# a_12690_27852# 0.010937f
C3754 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S a_2610_27852# 0.056787f
C3755 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G a_13842_27500# 0.033843f
C3756 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_3762_27148# 0.03422f
C3757 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S 0.027112f
C3758 a_15210_36300# SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.067588f
C3759 a_6282_36300# a_6282_35948# 0.010937f
C3760 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.224309f
C3761 a_17750_43288# uo_out[1] 0.066117f
C3762 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S VPWR 0.097536f
C3763 SUNSAR_CAPT8B_CV_0.XB07.XA6.A uo_out[7] 0.015483f
C3764 SUNSAR_SAR8B_CV_0.XA3.EN a_7650_34716# 0.066245f
C3765 SUNSAR_SAR8B_CV_0.EN a_8802_27148# 0.067588f
C3766 a_16362_35068# a_16362_34716# 0.010937f
C3767 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.014291f
C3768 SUNSAR_SAR8B_CV_0.XB1.XA4.GN ua[1] 0.762388f
C3769 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.036057f
C3770 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.012886f
C3771 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<5> 0.067851f
C3772 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.060807f
C3773 a_15230_43816# SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 0.071475f
C3774 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S 0.027953f
C3775 tt_um_TT06_SAR_done_0.DONE a_11342_40648# 0.084662f
C3776 a_5130_35068# VPWR 0.394528f
C3777 a_21402_28556# SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.066018f
C3778 a_10170_28556# a_10170_28204# 0.010937f
C3779 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR 0.042839f
C3780 a_3782_43816# VPWR 0.391817f
C3781 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.023976f
C3782 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_8822_41352# 0.058557f
C3783 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 0.803963f
C3784 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA20.CNO 0.252047f
C3785 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.301485f
C3786 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22790_42760# 0.13379f
C3787 a_5150_44168# a_5150_43816# 0.010937f
C3788 a_15230_44168# SUNSAR_CAPT8B_CV_0.XG12.QN 0.067588f
C3789 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S 0.050207f
C3790 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_16362_29612# 0.040867f
C3791 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.104122f
C3792 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S 0.011062f
C3793 SUNSAR_SAR8B_CV_0.D<4> VPWR 5.44394f
C3794 SUNSAR_CAPT8B_CV_0.XA4.MP1.G a_22790_41352# 0.036766f
C3795 a_5130_35948# VPWR 0.417826f
C3796 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B 3.57461f
C3797 a_7650_37180# SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.070936f
C3798 a_8802_37180# SUNSAR_SAR8B_CV_0.XA3.CEIN 0.040807f
C3799 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.030446f
C3800 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.073779f
C3801 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S 0.028011f
C3802 a_6282_27500# a_6282_27148# 0.010937f
C3803 a_3762_32076# VPWR 0.436368f
C3804 a_18882_35948# SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.066018f
C3805 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.432466f
C3806 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S 0.023798f
C3807 SUNSAR_CAPT8B_CV_0.XA6.A a_23942_43112# 0.067943f
C3808 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S 0.027192f
C3809 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA20.CPO 0.06466f
C3810 a_12582_2982# a_12582_2630# 0.010937f
C3811 a_3762_28204# VPWR 0.36179f
C3812 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.03343f
C3813 SUNSAR_SAR8B_CV_0.XA5.EN a_12690_28908# 0.068502f
C3814 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> a_7650_31196# 0.110962f
C3815 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR 0.898003f
C3816 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA20.CNO 0.024154f
C3817 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_6282_30316# 0.01727f
C3818 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.A 0.744161f
C3819 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S 0.055627f
C3820 SUNSAR_SAR8B_CV_0.XA4.XA12.A VPWR 0.723728f
C3821 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.142977f
C3822 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N a_12690_28908# 0.060353f
C3823 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.023017f
C3824 tt_um_TT06_SAR_done_0.x4.MP0.G a_28727_40659# 0.067434f
C3825 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR 4.24813f
C3826 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G a_2610_27148# 0.023111f
C3827 SUNSAR_SAR8B_CV_0.D<5> a_8802_32956# 0.017466f
C3828 a_11142_4566# SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.036098f
C3829 SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR 1.63909f
C3830 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.694484f
C3831 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.026917f
C3832 a_9990_4038# VPWR 0.379979f
C3833 a_13842_32956# SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.066018f
C3834 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.154232f
C3835 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_SAR8B_CV_0.D<2> 0.018133f
C3836 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S 0.089305f
C3837 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_6302_41880# 0.035868f
C3838 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43288# 0.03616f
C3839 a_22790_43992# a_22790_43640# 0.010937f
C3840 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S 0.024386f
C3841 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S 0.0111f
C3842 a_20270_40648# VPWR 0.493179f
C3843 a_17750_41000# a_17750_40648# 0.010937f
C3844 tt_um_TT06_SAR_done_0.DONE a_10190_40648# 0.066617f
C3845 a_3762_35068# VPWR 0.394528f
C3846 a_20250_28556# SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.071498f
C3847 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.098057f
C3848 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.061061f
C3849 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.057445f
C3850 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.788486f
C3851 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR 0.042839f
C3852 SUNSAR_CAPT8B_CV_0.XG12.QN uo_out[2] 0.249322f
C3853 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S 0.010488f
C3854 SUNSAR_SAR8B_CV_0.XA6.XA9.B a_17730_35068# 0.011912f
C3855 a_13842_35420# SUNSAR_SAR8B_CV_0.XA4.DONE 0.023111f
C3856 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S 0.021211f
C3857 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_41352# 0.060327f
C3858 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_8822_41352# 0.075505f
C3859 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.145483f
C3860 a_5130_35420# a_5130_35068# 0.010937f
C3861 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.026917f
C3862 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.011022f
C3863 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.11884f
C3864 a_23942_43112# a_23942_42760# 0.010937f
C3865 SUNSAR_SAR8B_CV_0.XA7.XA2.A a_21402_30316# 0.091063f
C3866 SUNSAR_SAR8B_CV_0.XA5.XA4.A a_15210_29612# 0.023777f
C3867 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S 0.155821f
C3868 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.038148f
C3869 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S VPWR 0.106927f
C3870 SUNSAR_SAR8B_CV_0.D<7> tt_um_TT06_SAR_done_0.DONE 0.292137f
C3871 a_3762_35948# VPWR 0.417826f
C3872 a_7650_37180# SUNSAR_SAR8B_CV_0.XA3.CEIN 0.023111f
C3873 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S 0.028011f
C3874 a_17730_35948# SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.072725f
C3875 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.12241f
C3876 SUNSAR_CAPT8B_CV_0.XA6.A a_22790_43112# 0.076609f
C3877 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S 0.027192f
C3878 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.038862f
C3879 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C3880 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.033149f
C3881 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.133602f
C3882 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR 0.898003f
C3883 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA6.A 0.649845f
C3884 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S 0.030221f
C3885 SUNSAR_SAR8B_CV_0.XA5.CEIN VPWR 2.30385f
C3886 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S 0.010682f
C3887 tt_um_TT06_SAR_done_0.x4.MP0.G a_27575_40659# 0.071058f
C3888 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR 0.097407f
C3889 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.3191f
C3890 a_11322_28204# a_11322_27852# 0.010937f
C3891 SUNSAR_SAR8B_CV_0.EN a_20250_30316# 0.076987f
C3892 a_13842_36300# SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.066018f
C3893 a_5130_36300# a_5130_35948# 0.010937f
C3894 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H a_15390_4566# 0.091934f
C3895 a_9990_4566# SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.072612f
C3896 SUNSAR_SAR8B_CV_0.SARP ua[1] 1.03265f
C3897 a_16382_43288# uo_out[2] 0.067687f
C3898 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR 0.104609f
C3899 a_15210_35068# a_15210_34716# 0.010937f
C3900 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.012236f
C3901 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_34716# 0.067815f
C3902 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S 0.055045f
C3903 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H ua[0] 0.023477f
C3904 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C3905 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A VPWR 2.50679f
C3906 a_12690_32956# SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.06825f
C3907 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.3401f
C3908 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S 0.010423f
C3909 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<6> 0.18141f
C3910 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.055045f
C3911 SUNSAR_CAPT8B_CV_0.XC08.XA5.A a_5150_41880# 0.024901f
C3912 SUNSAR_CAPT8B_CV_0.XC08.QN a_5150_43288# 0.024901f
C3913 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S 0.025128f
C3914 a_18902_40648# VPWR 0.491776f
C3915 tt_um_TT06_SAR_done_0.DONE a_8822_40648# 0.068187f
C3916 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S 0.073693f
C3917 a_8802_28556# a_8802_28204# 0.010937f
C3918 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.55251f
C3919 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S 0.054448f
C3920 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.015913f
C3921 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.112859f
C3922 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N VPWR 0.271482f
C3923 SUNSAR_CAPT8B_CV_0.XA7.MP0.G uio_oe[0] 0.064035f
C3924 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR 16.813599f
C3925 a_12690_35420# SUNSAR_SAR8B_CV_0.XA4.DONE 0.030547f
C3926 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S 0.021266f
C3927 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_SAR8B_CV_0.D<2> 0.393063f
C3928 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_3782_41880# 0.072658f
C3929 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_7670_41352# 0.080002f
C3930 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN 0.144331f
C3931 a_10170_27148# VPWR 0.470364f
C3932 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C3933 a_3782_44168# a_3782_43816# 0.010937f
C3934 a_13862_44168# SUNSAR_CAPT8B_CV_0.XF11.QN 0.066018f
C3935 SUNSAR_SAR8B_CV_0.XA7.XA2.A a_20250_30316# 0.127528f
C3936 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.019336f
C3937 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S VPWR 0.106927f
C3938 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.097975f
C3939 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S 0.053284f
C3940 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6519f
C3941 a_5130_27500# a_5130_27148# 0.010937f
C3942 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR 0.618979f
C3943 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.026506f
C3944 a_11142_2982# a_11142_2630# 0.010937f
C3945 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR 0.429492f
C3946 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.03343f
C3947 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_28908# 0.06753f
C3948 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C3949 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.SARP 0.032416f
C3950 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR 0.898003f
C3951 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S 0.044855f
C3952 SUNSAR_SAR8B_CV_0.XA3.XA12.A VPWR 0.720133f
C3953 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.142956f
C3954 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.064851f
C3955 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.316879f
C3956 SUNSAR_SAR8B_CV_0.EN a_18882_30316# 0.078124f
C3957 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.011917f
C3958 a_12690_36300# SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.068275f
C3959 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.036274f
C3960 SUNSAR_CAPT8B_CV_0.XA6.A VPWR 1.18734f
C3961 a_15230_43288# uo_out[2] 0.071088f
C3962 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S 0.026506f
C3963 SUNSAR_SAR8B_CV_0.XA2.XA9.B a_8802_33836# 0.023316f
C3964 SUNSAR_SAR8B_CV_0.EN a_5130_27148# 0.066018f
C3965 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_34716# 0.075712f
C3966 a_13950_4742# ua[0] 0.05378f
C3967 SUNSAR_SAR8B_CV_0.XB2.CKN VPWR 2.34497f
C3968 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<6> 0.064919f
C3969 uio_oe[0] uio_out[0] 1.55761f
C3970 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S 0.076714f
C3971 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S 0.036094f
C3972 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S 0.026188f
C3973 a_16382_41000# a_16382_40648# 0.010937f
C3974 tt_um_TT06_SAR_done_0.DONE a_7670_40648# 0.083091f
C3975 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.11263f
C3976 SUNSAR_CAPT8B_CV_0.XA7.MP0.G clk 0.030582f
C3977 SUNSAR_CAPT8B_CV_0.XF11.QN uo_out[3] 0.267395f
C3978 a_23942_43992# VPWR 0.388156f
C3979 SUNSAR_SAR8B_CV_0.XA0.XA9.B a_3762_34716# 0.023982f
C3980 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_SAR8B_CV_0.D<2> 0.241356f
C3981 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_2630_41880# 0.066018f
C3982 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA4.EN 0.051732f
C3983 a_3762_35420# a_3762_35068# 0.010937f
C3984 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.145483f
C3985 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C3986 a_8802_27148# VPWR 0.471462f
C3987 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.386137f
C3988 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03123f
C3989 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.CN1 0.083897f
C3990 a_22790_43112# a_22790_42760# 0.010937f
C3991 a_12710_44168# SUNSAR_CAPT8B_CV_0.XF11.QN 0.071093f
C3992 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S 0.050207f
C3993 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_13842_29612# 0.023777f
C3994 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S 0.150467f
C3995 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.276413f
C3996 SUNSAR_SAR8B_CV_0.D<5> VPWR 5.39174f
C3997 SUNSAR_SAR8B_CV_0.D<0> a_21422_41352# 0.079434f
C3998 SUNSAR_SAR8B_CV_0.XA20.XA12.Y VPWR 1.13456f
C3999 a_6282_37180# SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.069366f
C4000 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S 0.022628f
C4001 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR 0.324111f
C4002 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.01042f
C4003 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S 0.030434f
C4004 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.240612f
C4005 SUNSAR_CAPT8B_CV_0.XE10.XA7.C a_10190_42408# 0.076129f
C4006 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_11342_42408# 0.098561f
C4007 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S 0.027192f
C4008 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR 0.137646f
C4009 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.033149f
C4010 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.133602f
C4011 SUNSAR_SAR8B_CV_0.XA4.EN a_10170_28908# 0.073535f
C4012 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_5130_31196# 0.069193f
C4013 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.012661f
C4014 a_23942_42760# VPWR 0.388156f
C4015 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_21422_43288# 0.028213f
C4016 SUNSAR_SAR8B_CV_0.XA4.CEIN VPWR 1.06023f
C4017 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S 0.030434f
C4018 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S 0.010682f
C4019 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.064851f
C4020 a_10170_28204# a_10170_27852# 0.010937f
C4021 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR 4.25548f
C4022 SUNSAR_SAR8B_CV_0.D<0> a_20250_33836# 0.011975f
C4023 a_3762_36300# a_3762_35948# 0.010937f
C4024 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.011382f
C4025 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G a_16542_4566# 0.067588f
C4026 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.CKN 0.015687f
C4027 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR 0.035055f
C4028 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S 0.089305f
C4029 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.093524f
C4030 SUNSAR_SAR8B_CV_0.EN a_3762_27148# 0.067588f
C4031 a_13842_35068# a_13842_34716# 0.010937f
C4032 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.ENO 0.793076f
C4033 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C4034 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.026917f
C4035 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S 0.010423f
C4036 a_11322_32956# SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.066679f
C4037 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.036102f
C4038 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_3782_41880# 0.024901f
C4039 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.055045f
C4040 clk uio_out[0] 0.120689f
C4041 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S 0.055045f
C4042 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.63636f
C4043 SUNSAR_CAPT8B_CV_0.XB07.QN a_3782_43288# 0.024901f
C4044 a_13862_43816# SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.069905f
C4045 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S 0.050207f
C4046 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S 0.010745f
C4047 tt_um_TT06_SAR_done_0.DONE a_6302_40648# 0.084662f
C4048 a_18882_28556# SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.069927f
C4049 a_7650_28556# a_7650_28204# 0.010937f
C4050 SUNSAR_SAR8B_CV_0.XA20.XA10.Y VPWR 2.1352f
C4051 SUNSAR_SAR8B_CV_0.D<2> a_15210_34716# 0.070775f
C4052 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.112859f
C4053 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.381914f
C4054 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.060418f
C4055 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.078434f
C4056 SUNSAR_SAR8B_CV_0.XA0.XA9.B a_2610_34716# 0.047651f
C4057 a_11322_35420# SUNSAR_SAR8B_CV_0.XA3.DONE 0.031235f
C4058 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S 0.036491f
C4059 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_16362_35068# 0.129098f
C4060 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.018085f
C4061 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C4062 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> a_3762_32076# 0.02026f
C4063 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.301485f
C4064 a_2630_44168# a_2630_43816# 0.010937f
C4065 SUNSAR_SAR8B_CV_0.XA6.XA2.A a_18882_30316# 0.129098f
C4066 SUNSAR_SAR8B_CV_0.XA4.XA4.A a_12690_29612# 0.040867f
C4067 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.040976f
C4068 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S 0.011178f
C4069 SUNSAR_SAR8B_CV_0.D<0> a_20270_41352# 0.06659f
C4070 SUNSAR_SAR8B_CV_0.SARN a_13950_2630# 0.023457f
C4071 SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR 0.774301f
C4072 a_5130_37180# SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.067588f
C4073 a_6282_37180# SUNSAR_SAR8B_CV_0.XA2.CEIN 0.024074f
C4074 SUNSAR_SAR8B_CV_0.XA7.XA4.A VPWR 2.30002f
C4075 a_3762_27500# a_3762_27148# 0.010937f
C4076 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S 0.010335f
C4077 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.046858f
C4078 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN a_10190_42408# 0.031125f
C4079 a_9990_2982# a_9990_2630# 0.010937f
C4080 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VPWR 1.06002f
C4081 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.03343f
C4082 SUNSAR_SAR8B_CV_0.XA0.XA4.A a_2610_30316# 0.01727f
C4083 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_21422_43288# 0.067482f
C4084 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_20270_43288# 0.082288f
C4085 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.142977f
C4086 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N a_11322_28908# 0.060353f
C4087 SUNSAR_SAR8B_CV_0.XA2.XA12.A VPWR 0.723762f
C4088 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.021955f
C4089 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G a_20250_27852# 0.028807f
C4090 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G a_10170_27500# 0.033843f
C4091 a_11322_36300# SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.066704f
C4092 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S 0.050207f
C4093 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.088197f
C4094 a_13862_43288# uo_out[3] 0.073588f
C4095 a_20270_43288# VPWR 0.394205f
C4096 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.CKN 0.200119f
C4097 a_16542_4918# a_16542_4566# 0.010937f
C4098 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.018669f
C4099 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR 0.035055f
C4100 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G a_15390_4566# 0.071837f
C4101 SUNSAR_SAR8B_CV_0.EN a_2610_27148# 0.071606f
C4102 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_34716# 0.077282f
C4103 a_12582_4742# ua[1] 0.05378f
C4104 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.021241f
C4105 a_10170_32956# SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.067588f
C4106 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA20.CPO 0.068426f
C4107 SUNSAR_CAPT8B_CV_0.XB07.XA5.A a_2630_41880# 0.035868f
C4108 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S 0.089305f
C4109 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.D<7> 0.174845f
C4110 clk uio_oe[0] 0.260056f
C4111 ui_in[0] uio_out[0] 0.01872f
C4112 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.318734f
C4113 SUNSAR_CAPT8B_CV_0.XB07.QN a_2630_43288# 0.03616f
C4114 a_28727_41011# uio_oe[0] 0.051915f
C4115 a_15230_40648# VPWR 0.493179f
C4116 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S 0.024389f
C4117 a_15230_41000# a_15230_40648# 0.010937f
C4118 tt_um_TT06_SAR_done_0.DONE a_5150_40648# 0.066617f
C4119 a_17730_28556# SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.067588f
C4120 SUNSAR_SAR8B_CV_0.XA6.DONE VPWR 0.246222f
C4121 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.11263f
C4122 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S 0.034383f
C4123 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.054448f
C4124 SUNSAR_CAPT8B_CV_0.XI14.QN VPWR 0.901631f
C4125 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[4] 0.248612f
C4126 a_20250_30316# VPWR 0.403745f
C4127 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN 0.144331f
C4128 a_10170_35420# SUNSAR_SAR8B_CV_0.XA3.DONE 0.023111f
C4129 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S 0.010488f
C4130 SUNSAR_SAR8B_CV_0.XA5.XA9.B a_16362_35068# 0.011912f
C4131 SUNSAR_SAR8B_CV_0.XA5.XA9.A a_15210_35068# 0.089492f
C4132 a_2610_35420# a_2610_35068# 0.010937f
C4133 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.145483f
C4134 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C4135 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.0357f
C4136 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.CN1 0.083897f
C4137 SUNSAR_SAR8B_CV_0.XA7.CN0 a_20250_33836# 0.101833f
C4138 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03123f
C4139 a_11342_44168# SUNSAR_CAPT8B_CV_0.XE10.QN 0.069523f
C4140 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S 0.050207f
C4141 SUNSAR_SAR8B_CV_0.XA6.XA2.A a_17730_30316# 0.089492f
C4142 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S 0.030034f
C4143 SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR 0.780003f
C4144 a_5130_37180# SUNSAR_SAR8B_CV_0.XA2.CEIN 0.029627f
C4145 SUNSAR_SAR8B_CV_0.XA6.XA4.A VPWR 2.31167f
C4146 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S 0.023798f
C4147 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.12241f
C4148 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.032042f
C4149 a_16362_35948# SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.071154f
C4150 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR 0.138148f
C4151 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.068314f
C4152 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.033149f
C4153 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.133602f
C4154 SUNSAR_SAR8B_CV_0.XA3.EN a_8802_28908# 0.072087f
C4155 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA20.CNO 0.189429f
C4156 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_43288# 0.031221f
C4157 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S 0.010682f
C4158 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N a_10170_28908# 0.023475f
C4159 SUNSAR_SAR8B_CV_0.XA3.CEIN VPWR 2.30393f
C4160 SUNSAR_SAR8B_CV_0.SARP a_13950_4742# 0.041839f
C4161 a_8802_28204# a_8802_27852# 0.010937f
C4162 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.016387f
C4163 SUNSAR_SAR8B_CV_0.EN a_15210_30316# 0.078934f
C4164 a_10170_36300# SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.067588f
C4165 a_2610_36300# a_2610_35948# 0.010937f
C4166 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.013922f
C4167 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.040072f
C4168 a_18902_43288# VPWR 0.394205f
C4169 a_12710_43288# uo_out[3] 0.0663f
C4170 a_12690_35068# a_12690_34716# 0.010937f
C4171 SUNSAR_SAR8B_CV_0.XA1.EN a_2610_34716# 0.066245f
C4172 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA7.EN 0.026181f
C4173 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.098257f
C4174 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.290432f
C4175 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.016772f
C4176 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<7> 0.343916f
C4177 ui_in[0] uio_oe[0] 0.038407f
C4178 uo_out[0] uio_out[0] 0.201579f
C4179 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.093019f
C4180 tt_um_TT06_SAR_done_0.DONE uio_out[0] 0.058964f
C4181 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S 0.030434f
C4182 a_12710_43816# SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.073123f
C4183 a_13862_40648# VPWR 0.491776f
C4184 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S 0.026257f
C4185 tt_um_TT06_SAR_done_0.DONE a_3782_40648# 0.068187f
C4186 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S 0.073693f
C4187 a_6282_28556# a_6282_28204# 0.010937f
C4188 SUNSAR_SAR8B_CV_0.XA5.DONE VPWR 0.245452f
C4189 tt_um_TT06_SAR_done_0.DONE a_21402_35420# 0.038844f
C4190 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.112859f
C4191 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.010609f
C4192 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.098057f
C4193 a_21422_44168# uo_out[0] 0.040621f
C4194 SUNSAR_CAPT8B_CV_0.XH13.QN VPWR 0.901622f
C4195 a_18882_30316# VPWR 0.403802f
C4196 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.023976f
C4197 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_6302_41352# 0.078431f
C4198 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.011105f
C4199 a_5130_27148# VPWR 0.470364f
C4200 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C4201 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_21422_42760# 0.091344f
C4202 SUNSAR_SAR8B_CV_0.D<6> VPWR 5.42967f
C4203 a_10190_44168# SUNSAR_CAPT8B_CV_0.XE10.QN 0.067588f
C4204 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_11322_29612# 0.040867f
C4205 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.104122f
C4206 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.284482f
C4207 SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR 0.779986f
C4208 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.075315f
C4209 SUNSAR_SAR8B_CV_0.XA5.XA4.A VPWR 2.31167f
C4210 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.55251f
C4211 a_2610_27500# a_2610_27148# 0.010937f
C4212 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S 0.027563f
C4213 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.432466f
C4214 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_21422_42760# 0.031591f
C4215 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.527529f
C4216 a_15210_35948# SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.067588f
C4217 a_16542_3334# a_16542_2982# 0.010937f
C4218 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VPWR 1.06875f
C4219 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.SARN 0.64474f
C4220 SUNSAR_SAR8B_CV_0.XA20.XA3a.A SUNSAR_SAR8B_CV_0.XA20.CPO 0.11826f
C4221 a_20270_42760# VPWR 0.391454f
C4222 SUNSAR_SAR8B_CV_0.XA3.EN a_7650_28908# 0.068502f
C4223 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA6.CN1 0.024265f
C4224 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA20.CNO 0.191868f
C4225 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S 0.044855f
C4226 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.142956f
C4227 SUNSAR_SAR8B_CV_0.XA1.XA12.A VPWR 0.720114f
C4228 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S 0.064851f
C4229 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.019092f
C4230 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.010239f
C4231 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.31626f
C4232 SUNSAR_SAR8B_CV_0.D<6> a_5130_32956# 0.017466f
C4233 SUNSAR_SAR8B_CV_0.EN a_13842_30316# 0.077363f
C4234 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S 0.050207f
C4235 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR 0.104609f
C4236 a_15390_4918# a_15390_4566# 0.010937f
C4237 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S 0.055045f
C4238 SUNSAR_SAR8B_CV_0.EN a_20250_27500# 0.073293f
C4239 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.146492f
C4240 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.CNO 0.092221f
C4241 a_8802_32956# SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.066018f
C4242 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S 0.089305f
C4243 ui_in[0] clk 0.25248f
C4244 uo_out[1] uio_out[0] 0.064738f
C4245 uo_out[0] uio_oe[0] 0.670799f
C4246 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N a_2610_29612# 0.031412f
C4247 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S 0.026117f
C4248 a_13862_41000# a_13862_40648# 0.010937f
C4249 tt_um_TT06_SAR_done_0.DONE a_2630_40648# 0.08295f
C4250 SUNSAR_SAR8B_CV_0.XA4.DONE VPWR 0.246222f
C4251 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.2165f
C4252 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C4253 tt_um_TT06_SAR_done_0.DONE a_20250_35420# 0.024133f
C4254 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S 0.028452f
C4255 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38424f
C4256 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.11263f
C4257 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.02121f
C4258 SUNSAR_CAPT8B_CV_0.XG12.QN VPWR 0.901622f
C4259 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[5] 0.248535f
C4260 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[6] 0.029694f
C4261 a_20270_44168# uo_out[0] 0.035586f
C4262 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA3.EN 0.051732f
C4263 a_8802_35420# SUNSAR_SAR8B_CV_0.XA2.DONE 0.023111f
C4264 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_6302_41352# 0.060327f
C4265 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_5150_41352# 0.077076f
C4266 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.B 0.545186f
C4267 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.145483f
C4268 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.028261f
C4269 a_3762_27148# VPWR 0.471462f
C4270 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.107427f
C4271 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.CN1 0.083897f
C4272 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03107f
C4273 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_20270_42760# 0.111734f
C4274 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S 0.050207f
C4275 SUNSAR_SAR8B_CV_0.XA5.XA2.A a_16362_30316# 0.091063f
C4276 SUNSAR_SAR8B_CV_0.XA3.XA4.A a_10170_29612# 0.023777f
C4277 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S 0.155821f
C4278 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.038148f
C4279 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S VPWR 0.106927f
C4280 SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR 0.780003f
C4281 a_3762_37180# SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.066018f
C4282 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S 0.022425f
C4283 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.073665f
C4284 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.030459f
C4285 SUNSAR_SAR8B_CV_0.XA4.XA4.A VPWR 2.31167f
C4286 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.026506f
C4287 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN a_20270_42760# 0.031082f
C4288 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR 0.137646f
C4289 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.137745f
C4290 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_23922_30844# 0.100515f
C4291 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.XA2.A 0.133602f
C4292 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.012782f
C4293 a_18902_42760# VPWR 0.391454f
C4294 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S 0.030221f
C4295 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.649845f
C4296 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S 0.010682f
C4297 SUNSAR_SAR8B_CV_0.XA2.CEIN VPWR 1.06023f
C4298 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_23922_35420# 0.079313f
C4299 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G a_8802_27500# 0.033843f
C4300 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G a_18882_27852# 0.028807f
C4301 a_7650_28204# a_7650_27852# 0.010937f
C4302 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR 0.097407f
C4303 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.089645f
C4304 a_8802_36300# SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.066018f
C4305 SUNSAR_SAR8B_CV_0.D<1> a_18882_33836# 0.011974f
C4306 a_11342_43288# uo_out[4] 0.067687f
C4307 SUNSAR_SAR8B_CV_0.EN a_18882_27500# 0.071722f
C4308 a_11322_35068# a_11322_34716# 0.010937f
C4309 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA6.EN 1.2771f
C4310 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.098257f
C4311 SUNSAR_SAR8B_CV_0.XB1.CKN VPWR 2.34497f
C4312 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.021241f
C4313 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.031163f
C4314 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA20.CPO 0.058427f
C4315 a_7650_32956# SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.06825f
C4316 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.055045f
C4317 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S 0.055045f
C4318 uo_out[2] uio_out[0] 0.052955f
C4319 uo_out[1] uio_oe[0] 0.432144f
C4320 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.233892f
C4321 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S 0.025128f
C4322 a_16362_28556# SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.066018f
C4323 a_5130_28556# a_5130_28204# 0.010937f
C4324 SUNSAR_SAR8B_CV_0.XA3.DONE VPWR 0.245452f
C4325 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.242472f
C4326 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.010771f
C4327 SUNSAR_SAR8B_CV_0.D<3> a_13842_34716# 0.069204f
C4328 SUNSAR_CAPT8B_CV_0.XF11.QN VPWR 0.901622f
C4329 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[6] 0.029694f
C4330 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[7] 0.010491f
C4331 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S 0.036491f
C4332 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S 0.036164f
C4333 a_7650_35420# SUNSAR_SAR8B_CV_0.XA2.DONE 0.030547f
C4334 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN 0.381205f
C4335 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_13842_35068# 0.091063f
C4336 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_41352# 0.058557f
C4337 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.020079f
C4338 a_8822_44168# SUNSAR_CAPT8B_CV_0.XD09.QN 0.066018f
C4339 a_23942_44344# a_23942_43992# 0.010937f
C4340 SUNSAR_SAR8B_CV_0.XA5.XA2.A a_15210_30316# 0.127528f
C4341 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.474658f
C4342 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S VPWR 0.106927f
C4343 SUNSAR_SAR8B_CV_0.D<1> a_18902_41352# 0.06816f
C4344 SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR 0.779986f
C4345 a_2610_37180# SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.070936f
C4346 a_3762_37180# SUNSAR_SAR8B_CV_0.XA1.CEIN 0.040807f
C4347 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.098006f
C4348 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S 0.050648f
C4349 SUNSAR_SAR8B_CV_0.XA3.XA4.A VPWR 2.31167f
C4350 a_21402_27852# a_21402_27500# 0.010937f
C4351 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S 0.027192f
C4352 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.412143f
C4353 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_8822_42408# 0.031125f
C4354 a_15390_3334# a_15390_2982# 0.010937f
C4355 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B a_16542_2630# 0.015402f
C4356 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VPWR 1.05322f
C4357 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_23922_33132# 0.067588f
C4358 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C4359 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.162703f
C4360 SUNSAR_SAR8B_CV_0.XA20.XA3a.A a_22770_30844# 0.066264f
C4361 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_28908# 0.06753f
C4362 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S 0.055627f
C4363 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.744161f
C4364 SUNSAR_SAR8B_CV_0.XA0.XA12.A VPWR 0.728492f
C4365 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.142977f
C4366 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S 0.030434f
C4367 SUNSAR_SAR8B_CV_0.CK_SAMPLE a_22770_35420# 0.067244f
C4368 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S 0.050207f
C4369 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR 0.112858f
C4370 a_7650_36300# SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.068275f
C4371 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.032857f
C4372 a_15230_43288# VPWR 0.394205f
C4373 a_10190_43288# uo_out[4] 0.071088f
C4374 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.22339f
C4375 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.036274f
C4376 SUNSAR_SAR8B_CV_0.XA1.XA9.B a_5130_33836# 0.023316f
C4377 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A VPWR 2.50679f
C4378 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.152052f
C4379 uo_out[3] uio_out[0] 0.057862f
C4380 uo_out[2] uio_oe[0] 0.267754f
C4381 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S 0.076714f
C4382 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S 0.036094f
C4383 a_10190_40648# VPWR 0.493224f
C4384 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.SARP 0.054401f
C4385 tt_um_TT06_SAR_done_0.DONE ui_in[0] 0.201929f
C4386 a_12710_41000# a_12710_40648# 0.010937f
C4387 a_15210_28556# SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.071498f
C4388 SUNSAR_SAR8B_CV_0.XA2.DONE VPWR 0.246222f
C4389 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.303978f
C4390 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.098057f
C4391 a_18902_44168# uo_out[1] 0.035338f
C4392 SUNSAR_CAPT8B_CV_0.XE10.QN VPWR 0.901622f
C4393 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[6] 0.258218f
C4394 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.55251f
C4395 a_23922_27148# a_23922_26796# 0.010937f
C4396 a_15210_30316# VPWR 0.404384f
C4397 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_SAR8B_CV_0.D<3> 0.241356f
C4398 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.321724f
C4399 SUNSAR_SAR8B_CV_0.XA4.XA9.A a_12690_35068# 0.127528f
C4400 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.145483f
C4401 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C4402 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.CN1 0.083897f
C4403 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 0.803935f
C4404 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.038099f
C4405 TIE_L SUNSAR_CAPT8B_CV_0.XI14.QN 0.013038f
C4406 a_7670_44168# SUNSAR_CAPT8B_CV_0.XD09.QN 0.071093f
C4407 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_8802_29612# 0.023777f
C4408 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S 0.150467f
C4409 SUNSAR_SAR8B_CV_0.D<7> VPWR 3.7939f
C4410 SUNSAR_SAR8B_CV_0.D<1> a_17750_41352# 0.077864f
C4411 SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR 0.780003f
C4412 SUNSAR_SAR8B_CV_0.SARP a_22770_28556# 0.023717f
C4413 a_2610_37180# SUNSAR_SAR8B_CV_0.XA1.CEIN 0.023111f
C4414 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.074964f
C4415 SUNSAR_SAR8B_CV_0.XA2.XA4.A VPWR 2.31167f
C4416 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_8822_42408# 0.074559f
C4417 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN a_7670_42408# 0.100131f
C4418 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S 0.027664f
C4419 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.031231f
C4420 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR 0.138148f
C4421 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S 0.03027f
C4422 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.021464f
C4423 SUNSAR_SAR8B_CV_0.XA20.XA10.Y a_22770_33132# 0.073025f
C4424 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.133602f
C4425 SUNSAR_SAR8B_CV_0.XA7.XA4.A a_21402_31196# 0.010411f
C4426 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.01601f
C4427 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S 0.012065f
C4428 SUNSAR_SAR8B_CV_0.XA2.EN a_5130_28908# 0.073535f
C4429 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.SARP 0.032814f
C4430 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S 0.026885f
C4431 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_18902_43288# 0.031221f
C4432 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S 0.030434f
C4433 SUNSAR_SAR8B_CV_0.XA1.CEIN VPWR 2.30575f
C4434 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S 0.010682f
C4435 a_6282_28204# a_6282_27852# 0.010937f
C4436 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR 0.112858f
C4437 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.040072f
C4438 SUNSAR_SAR8B_CV_0.EN a_10170_30316# 0.078934f
C4439 a_13862_43288# VPWR 0.394205f
C4440 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR 0.104609f
C4441 a_16542_4918# SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.030771f
C4442 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G a_11142_4566# 0.073407f
C4443 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.224309f
C4444 a_10170_35068# a_10170_34716# 0.010937f
C4445 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA5.EN 0.026181f
C4446 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H ua[1] 0.023477f
C4447 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.419738f
C4448 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR 0.665179f
C4449 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.058243f
C4450 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.339883f
C4451 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA7.CN1 0.010488f
C4452 a_6282_32956# SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.066679f
C4453 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.055045f
C4454 uo_out[4] uio_out[0] 0.013711f
C4455 a_11342_43816# SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.071553f
C4456 uo_out[3] uio_oe[0] 0.212351f
C4457 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 0.093019f
C4458 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S 0.050207f
C4459 a_8822_40648# VPWR 0.491776f
C4460 a_23942_41000# ui_in[0] 0.066166f
C4461 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S 0.073693f
C4462 a_3762_28556# a_3762_28204# 0.010937f
C4463 SUNSAR_SAR8B_CV_0.XA1.DONE VPWR 0.245452f
C4464 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.56958f
C4465 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.054448f
C4466 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.13078f
C4467 a_17750_44168# uo_out[1] 0.041262f
C4468 SUNSAR_CAPT8B_CV_0.XD09.QN VPWR 0.901622f
C4469 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[7] 0.016809f
C4470 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_SAR8B_CV_0.D<3> 0.393049f
C4471 a_13842_30316# VPWR 0.404384f
C4472 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.023976f
C4473 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S 0.021266f
C4474 a_6282_35420# SUNSAR_SAR8B_CV_0.XA1.DONE 0.031235f
C4475 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN 0.144331f
C4476 a_20250_27500# VPWR 0.382397f
C4477 TIE_L SUNSAR_CAPT8B_CV_0.XH13.QN 0.013038f
C4478 a_22790_44344# a_22790_43992# 0.010937f
C4479 SUNSAR_SAR8B_CV_0.XA4.XA2.A a_13842_30316# 0.129098f
C4480 SUNSAR_SAR8B_CV_0.XA2.XA4.A a_7650_29612# 0.040867f
C4481 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S 0.011062f
C4482 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 a_22770_29964# 0.031884f
C4483 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.040976f
C4484 SUNSAR_SAR8B_CV_0.SARN a_13950_2982# 0.037174f
C4485 SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR 0.779986f
C4486 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S 0.028011f
C4487 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.064969f
C4488 SUNSAR_SAR8B_CV_0.XA1.XA4.A VPWR 2.31167f
C4489 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.55251f
C4490 a_20250_27852# a_20250_27500# 0.010937f
C4491 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.432466f
C4492 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S 0.012357f
C4493 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S 0.073313f
C4494 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.010335f
C4495 a_13842_35948# SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.066018f
C4496 a_13950_3334# a_13950_2982# 0.010937f
C4497 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VPWR 1.06875f
C4498 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA7.CP0 0.017772f
C4499 a_15230_42760# VPWR 0.391454f
C4500 a_21402_32076# SUNSAR_SAR8B_CV_0.XA7.CN1 0.06792f
C4501 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA4.CN1 0.024265f
C4502 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_43288# 0.069053f
C4503 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_18902_43288# 0.080718f
C4504 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.142956f
C4505 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.023017f
C4506 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR 4.249f
C4507 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S 0.050207f
C4508 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A 0.201839f
C4509 a_6282_36300# SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.066704f
C4510 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.316879f
C4511 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.090136f
C4512 SUNSAR_SAR8B_CV_0.EN a_8802_30316# 0.077363f
C4513 a_8822_43288# uo_out[5] 0.072658f
C4514 SUNSAR_CAPT8B_CV_0.XA6.B clk 0.07088f
C4515 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G a_9990_4566# 0.066018f
C4516 a_15390_4918# SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.015779f
C4517 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H a_11142_4566# 0.090364f
C4518 a_21402_35068# SUNSAR_SAR8B_CV_0.XA7.ENO 0.066018f
C4519 SUNSAR_SAR8B_CV_0.EN a_15210_27500# 0.073293f
C4520 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S 0.055045f
C4521 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S 0.026506f
C4522 a_16542_4566# VPWR 0.413433f
C4523 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.724892f
C4524 a_5130_32956# SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.067588f
C4525 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S 0.089305f
C4526 uo_out[5] uio_out[0] 0.109219f
C4527 uo_out[4] uio_oe[0] 0.550054f
C4528 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.318734f
C4529 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S 0.024386f
C4530 uo_out[1] uo_out[0] 0.355472f
C4531 a_22790_41000# ui_in[0] 0.074344f
C4532 a_11342_41000# a_11342_40648# 0.010937f
C4533 SUNSAR_SAR8B_CV_0.XA0.DONE VPWR 0.247527f
C4534 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.86675f
C4535 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.012048f
C4536 a_22770_27148# a_22770_26796# 0.010937f
C4537 SUNSAR_CAPT8B_CV_0.XC08.QN VPWR 0.901622f
C4538 SUNSAR_CAPT8B_CV_0.XB07.QN uo_out[7] 0.263255f
C4539 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S 0.010488f
C4540 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S 0.021211f
C4541 a_5130_35420# SUNSAR_SAR8B_CV_0.XA1.DONE 0.023111f
C4542 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA2.EN 0.051732f
C4543 SUNSAR_SAR8B_CV_0.XA4.XA9.B a_12690_35068# 0.011912f
C4544 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.145483f
C4545 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C4546 a_18882_27500# VPWR 0.382189f
C4547 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.016209f
C4548 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.CN1 0.083897f
C4549 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_18902_42760# 0.113305f
C4550 a_6302_44168# SUNSAR_CAPT8B_CV_0.XC08.QN 0.069523f
C4551 SUNSAR_SAR8B_CV_0.XA4.XA2.A a_12690_30316# 0.089492f
C4552 SUNSAR_SAR8B_CV_0.XA7.ENO a_20250_28204# 0.016912f
C4553 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S 0.030034f
C4554 a_23942_41880# VPWR 0.398828f
C4555 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.015927f
C4556 SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR 0.784656f
C4557 a_21402_37532# a_21402_37180# 0.010937f
C4558 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S 0.028011f
C4559 SUNSAR_SAR8B_CV_0.XA0.XA4.A VPWR 2.31167f
C4560 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.12241f
C4561 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_18902_42760# 0.031082f
C4562 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.062692f
C4563 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.527529f
C4564 a_12690_35948# SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.072725f
C4565 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR 0.137646f
C4566 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C4567 SUNSAR_SAR8B_CV_0.EN uio_oe[0] 0.010306f
C4568 SUNSAR_SAR8B_CV_0.CK_SAMPLE clk 0.031633f
C4569 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.133602f
C4570 SUNSAR_SAR8B_CV_0.XA1.EN a_3762_28908# 0.072087f
C4571 a_13862_42760# VPWR 0.391454f
C4572 a_20250_32076# SUNSAR_SAR8B_CV_0.XA7.CN1 0.067588f
C4573 ui_in[2] ui_in[1] 0.023797f
C4574 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_17750_43288# 0.028213f
C4575 a_20250_37180# VPWR 0.469114f
C4576 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S 0.010682f
C4577 a_5130_28204# a_5130_27852# 0.010937f
C4578 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR 0.097407f
C4579 a_5130_36300# SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.067588f
C4580 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.09968f
C4581 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR 0.035055f
C4582 a_7670_43288# uo_out[5] 0.066117f
C4583 a_11142_4918# a_11142_4566# 0.010937f
C4584 a_20250_35068# SUNSAR_SAR8B_CV_0.XA7.ENO 0.071277f
C4585 a_8802_35068# a_8802_34716# 0.010937f
C4586 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA4.EN 1.2771f
C4587 SUNSAR_SAR8B_CV_0.EN a_13842_27500# 0.071722f
C4588 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S 0.055045f
C4589 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_25610_2722# 0.029253f
C4590 a_13950_5094# ua[0] 0.053744f
C4591 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.419738f
C4592 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.058243f
C4593 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.036057f
C4594 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.63636f
C4595 uo_out[6] uio_out[0] 0.010745f
C4596 VPWR ua[0] 0.629451f
C4597 a_10190_43816# SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.071475f
C4598 uo_out[5] uio_oe[0] 1.55329f
C4599 a_13842_28556# SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.069927f
C4600 a_2610_28556# a_2610_28204# 0.010937f
C4601 a_23922_35420# VPWR 0.416528f
C4602 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.ENO 0.409849f
C4603 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.352238f
C4604 a_16382_44168# uo_out[2] 0.040603f
C4605 SUNSAR_CAPT8B_CV_0.XB07.QN VPWR 0.901622f
C4606 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_3782_41352# 0.058557f
C4607 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.030426f
C4608 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_17750_42760# 0.089774f
C4609 a_5150_44168# SUNSAR_CAPT8B_CV_0.XC08.QN 0.067588f
C4610 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_6282_29612# 0.040867f
C4611 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.104122f
C4612 a_23922_36300# VPWR 0.472384f
C4613 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S 0.050207f
C4614 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S 0.053284f
C4615 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.030446f
C4616 SUNSAR_SAR8B_CV_0.XA20.XA3a.A VPWR 4.6743f
C4617 a_18882_27852# a_18882_27500# 0.010937f
C4618 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_42760# 0.031591f
C4619 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA20.CNO 0.066214f
C4620 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.205884f
C4621 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S 0.023798f
C4622 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 0.59598f
C4623 a_12582_3334# a_12582_2982# 0.010937f
C4624 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VPWR 1.05322f
C4625 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S 0.028026f
C4626 SUNSAR_SAR8B_CV_0.CK_SAMPLE ui_in[0] 0.079428f
C4627 SUNSAR_SAR8B_CV_0.XA1.EN a_2610_28908# 0.068502f
C4628 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARP 0.033467f
C4629 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S 0.030434f
C4630 a_18882_37180# VPWR 0.473682f
C4631 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.142977f
C4632 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G a_5130_27500# 0.033843f
C4633 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G a_15210_27852# 0.028807f
C4634 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S 0.050207f
C4635 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.175332f
C4636 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR 0.035055f
C4637 a_10190_43288# VPWR 0.394205f
C4638 a_16542_4918# SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.066018f
C4639 SUNSAR_SAR8B_CV_0.XA0.XA9.B a_3762_33836# 0.023316f
C4640 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24750_2768# 0.172147f
C4641 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR 0.665179f
C4642 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.154232f
C4643 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.723071f
C4644 a_3762_32956# SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.066018f
C4645 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S 0.089305f
C4646 uo_out[7] uio_out[0] 0.07272f
C4647 VPWR ua[1] 0.349347f
C4648 uo_out[2] uo_out[1] 0.06895f
C4649 uo_out[6] uio_oe[0] 0.057603f
C4650 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S 0.076714f
C4651 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S 0.030434f
C4652 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.010898f
C4653 a_5150_40648# VPWR 0.493192f
C4654 a_21422_41000# tt_um_TT06_SAR_done_0.DONE 0.06916f
C4655 a_10190_41000# a_10190_40648# 0.010937f
C4656 a_12690_28556# SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.067588f
C4657 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.42106f
C4658 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.054448f
C4659 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.033093f
C4660 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 54.2165f
C4661 a_21402_27148# a_21402_26796# 0.010937f
C4662 a_10170_30316# VPWR 0.404384f
C4663 a_15230_44168# uo_out[2] 0.035338f
C4664 SUNSAR_CAPT8B_CV_0.XA7.MP0.G VPWR 0.667429f
C4665 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN a_2630_41352# 0.060327f
C4666 SUNSAR_CAPT8B_CV_0.XB07.XA7.C a_3782_41352# 0.075505f
C4667 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_21422_41880# 0.070877f
C4668 a_3762_35420# SUNSAR_SAR8B_CV_0.XA0.DONE 0.023111f
C4669 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN 0.144331f
C4670 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.145483f
C4671 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C4672 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 0.803963f
C4673 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.101323f
C4674 SUNSAR_SAR8B_CV_0.XA3.XA2.A a_11322_30316# 0.091063f
C4675 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S 0.011494f
C4676 SUNSAR_SAR8B_CV_0.XA1.XA4.A a_5130_29612# 0.023777f
C4677 SUNSAR_SAR8B_CV_0.XA7.EN a_18882_28204# 0.017441f
C4678 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S 0.155821f
C4679 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.038148f
C4680 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.276413f
C4681 SUNSAR_SAR8B_CV_0.D<2> a_16382_41352# 0.079434f
C4682 a_20250_37532# a_20250_37180# 0.010937f
C4683 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S 0.022628f
C4684 SUNSAR_SAR8B_CV_0.EN a_20250_29612# 0.142592f
C4685 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.746324f
C4686 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR 0.138148f
C4687 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.026794f
C4688 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.CN0 0.036885f
C4689 SUNSAR_SAR8B_CV_0.EN ui_in[0] 0.968121f
C4690 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.133602f
C4691 SUNSAR_SAR8B_CV_0.XA6.XA4.A a_17730_31196# 0.010411f
C4692 a_18882_32076# SUNSAR_SAR8B_CV_0.XA6.CN1 0.066018f
C4693 SUNSAR_SAR8B_CV_0.CK_SAMPLE tt_um_TT06_SAR_done_0.DONE 0.403015f
C4694 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S 0.026885f
C4695 ui_in[3] ui_in[2] 0.023797f
C4696 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N a_8802_28908# 0.023475f
C4697 a_3762_28204# a_3762_27852# 0.010937f
C4698 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR 4.26707f
C4699 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA6.A 0.040072f
C4700 a_3762_36300# SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.066018f
C4701 SUNSAR_SAR8B_CV_0.D<2> a_15210_33836# 0.011975f
C4702 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.297124f
C4703 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.021942f
C4704 SUNSAR_SAR8B_CV_0.EN a_5130_30316# 0.078934f
C4705 a_8822_43288# VPWR 0.394205f
C4706 a_15390_4918# SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.099734f
C4707 a_9990_4918# a_9990_4566# 0.010937f
C4708 a_6302_43288# uo_out[6] 0.068411f
C4709 a_18882_35068# SUNSAR_SAR8B_CV_0.XA7.EN 0.069707f
C4710 a_7650_35068# a_7650_34716# 0.010937f
C4711 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA3.EN 0.026181f
C4712 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B m3_24678_2768# 0.0666f
C4713 a_12582_5094# ua[1] 0.053744f
C4714 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.046398f
C4715 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.031784f
C4716 a_2610_32956# SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.06825f
C4717 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S 0.010423f
C4718 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA20.CNO 0.066819f
C4719 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.3401f
C4720 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.055045f
C4721 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_21422_41880# 0.067588f
C4722 uo_out[7] uio_oe[0] 0.43252f
C4723 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S 0.055045f
C4724 VPWR uio_out[0] 0.408488f
C4725 a_3782_40648# VPWR 0.491776f
C4726 a_20270_41000# tt_um_TT06_SAR_done_0.DONE 0.067588f
C4727 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.018236f
C4728 ua[2] VGND 0.117454f
C4729 ua[3] VGND 0.117454f
C4730 ua[4] VGND 0.118698f
C4731 ua[5] VGND 0.120088f
C4732 ua[6] VGND 0.120088f
C4733 ua[7] VGND 0.111009f
C4734 ena VGND 0.073297f
C4735 rst_n VGND 0.048301f
C4736 ui_in[1] VGND 0.048271f
C4737 ui_in[2] VGND 0.048424f
C4738 ui_in[3] VGND 0.043149f
C4739 ui_in[4] VGND 0.047461f
C4740 ui_in[5] VGND 0.047747f
C4741 ui_in[6] VGND 0.044024f
C4742 ui_in[7] VGND 0.044024f
C4743 uio_in[0] VGND 0.047253f
C4744 uio_in[1] VGND 0.045497f
C4745 uio_in[2] VGND 0.047751f
C4746 uio_in[3] VGND 0.046379f
C4747 uio_in[4] VGND 0.044575f
C4748 uio_in[5] VGND 0.044575f
C4749 uio_in[6] VGND 0.044575f
C4750 uio_in[7] VGND 0.046165f
C4751 uio_out[1] VGND 0.037696f
C4752 uio_out[2] VGND 0.037696f
C4753 uio_out[3] VGND 0.037696f
C4754 uio_out[4] VGND 0.037696f
C4755 uio_out[5] VGND 0.037696f
C4756 uio_out[6] VGND 0.037822f
C4757 uio_out[7] VGND 0.037696f
C4758 uio_oe[1] VGND 0.037696f
C4759 uio_oe[2] VGND 0.037696f
C4760 uio_oe[3] VGND 0.037696f
C4761 uio_oe[4] VGND 0.03773f
C4762 uio_oe[5] VGND 0.037932f
C4763 uio_oe[6] VGND 0.037696f
C4764 uio_oe[7] VGND 0.062293f
C4765 ua[0] VGND 7.65072f
C4766 ua[1] VGND 7.01222f
C4767 uio_out[0] VGND 8.429111f
C4768 uio_oe[0] VGND 7.8235f
C4769 clk VGND 7.0308f
C4770 ui_in[0] VGND 6.39197f
C4771 uo_out[0] VGND 2.40292f
C4772 uo_out[1] VGND 1.50319f
C4773 uo_out[2] VGND 1.42895f
C4774 uo_out[3] VGND 1.68048f
C4775 uo_out[4] VGND 1.55276f
C4776 uo_out[5] VGND 1.75883f
C4777 uo_out[6] VGND 2.73387f
C4778 uo_out[7] VGND 3.23518f
C4779 VPWR VGND 0.955234p
C4780 m4_6696_44772# VGND 0.016293f $ **FLOATING
C4781 m4_5739_44772# VGND 0.016293f $ **FLOATING
C4782 TIE_L1 VGND 1.33513f
C4783 TIE_L2 VGND 1.65212f
C4784 m4_798_44892# VGND 0.015387f $ **FLOATING
C4785 m3_25610_2722# VGND 0.186542f $ **FLOATING
C4786 m1_14848_7490# VGND 0.145299f $ **FLOATING
C4787 li_16096_7824# VGND 0.039377f $ **FLOATING
C4788 li_11088_7824# VGND 0.039377f $ **FLOATING
C4789 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93682f
C4790 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93682f
C4791 li_16096_8428# VGND 0.0355f $ **FLOATING
C4792 li_11088_8428# VGND 0.0355f $ **FLOATING
C4793 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.555001f
C4794 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.555001f
C4795 li_16096_9032# VGND 0.0355f $ **FLOATING
C4796 li_11088_9032# VGND 0.0355f $ **FLOATING
C4797 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.335569f
C4798 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.335569f
C4799 li_16096_9636# VGND 0.035528f $ **FLOATING
C4800 li_11088_9636# VGND 0.035528f $ **FLOATING
C4801 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.4697f
C4802 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.4697f
C4803 li_16096_10240# VGND 0.035574f $ **FLOATING
C4804 li_11088_10240# VGND 0.035574f $ **FLOATING
C4805 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43607f
C4806 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43607f
C4807 li_16096_10844# VGND 0.033763f $ **FLOATING
C4808 li_11088_10844# VGND 0.033763f $ **FLOATING
C4809 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67818f
C4810 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67818f
C4811 li_16096_11224# VGND 0.037139f $ **FLOATING
C4812 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.66914f
C4813 li_11088_11224# VGND 0.037139f $ **FLOATING
C4814 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.66914f
C4815 li_16096_11828# VGND 0.035704f $ **FLOATING
C4816 li_11088_11828# VGND 0.035704f $ **FLOATING
C4817 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.5762f
C4818 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.5762f
C4819 li_16096_12432# VGND 0.035549f $ **FLOATING
C4820 li_11088_12432# VGND 0.035549f $ **FLOATING
C4821 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33485f
C4822 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33485f
C4823 li_16096_13036# VGND 0.0355f $ **FLOATING
C4824 li_11088_13036# VGND 0.0355f $ **FLOATING
C4825 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.4697f
C4826 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.4697f
C4827 li_16096_13640# VGND 0.0355f $ **FLOATING
C4828 li_11088_13640# VGND 0.0355f $ **FLOATING
C4829 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43607f
C4830 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43607f
C4831 li_16096_14244# VGND 0.033227f $ **FLOATING
C4832 li_11088_14244# VGND 0.033227f $ **FLOATING
C4833 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67818f
C4834 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67818f
C4835 li_16096_14624# VGND 0.033227f $ **FLOATING
C4836 li_11088_14624# VGND 0.033227f $ **FLOATING
C4837 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.66914f
C4838 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.66914f
C4839 li_16096_15228# VGND 0.0355f $ **FLOATING
C4840 li_11088_15228# VGND 0.0355f $ **FLOATING
C4841 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.5768f
C4842 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.5768f
C4843 li_16096_15832# VGND 0.0355f $ **FLOATING
C4844 li_11088_15832# VGND 0.0355f $ **FLOATING
C4845 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33485f
C4846 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33485f
C4847 li_16096_16436# VGND 0.0355f $ **FLOATING
C4848 li_11088_16436# VGND 0.0355f $ **FLOATING
C4849 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.4697f
C4850 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.4697f
C4851 li_16096_17040# VGND 0.0355f $ **FLOATING
C4852 li_11088_17040# VGND 0.0355f $ **FLOATING
C4853 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43607f
C4854 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43607f
C4855 li_16096_17644# VGND 0.033227f $ **FLOATING
C4856 li_11088_17644# VGND 0.033227f $ **FLOATING
C4857 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67818f
C4858 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67818f
C4859 li_16096_18024# VGND 0.033227f $ **FLOATING
C4860 li_11088_18024# VGND 0.033227f $ **FLOATING
C4861 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.66914f
C4862 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.66914f
C4863 li_16096_18628# VGND 0.0355f $ **FLOATING
C4864 li_11088_18628# VGND 0.0355f $ **FLOATING
C4865 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.5735f
C4866 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.5735f
C4867 li_16096_19232# VGND 0.0355f $ **FLOATING
C4868 li_11088_19232# VGND 0.0355f $ **FLOATING
C4869 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33485f
C4870 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33485f
C4871 li_16096_19836# VGND 0.0355f $ **FLOATING
C4872 li_11088_19836# VGND 0.0355f $ **FLOATING
C4873 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.472599f
C4874 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.472599f
C4875 li_16096_20440# VGND 0.0355f $ **FLOATING
C4876 li_11088_20440# VGND 0.0355f $ **FLOATING
C4877 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.44327f
C4878 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44327f
C4879 li_16096_21044# VGND 0.039377f $ **FLOATING
C4880 li_11088_21044# VGND 0.039377f $ **FLOATING
C4881 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.38664f
C4882 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.3834f
C4883 a_16542_2630# VGND 0.096631f $ **FLOATING
C4884 a_15390_2630# VGND 0.543325f $ **FLOATING
C4885 a_13950_2630# VGND 0.428911f $ **FLOATING
C4886 a_12582_2630# VGND 0.428496f $ **FLOATING
C4887 a_11142_2630# VGND 0.544481f $ **FLOATING
C4888 a_9990_2630# VGND 0.096631f $ **FLOATING
C4889 a_15390_2982# VGND 0.492315f $ **FLOATING
C4890 a_13950_2982# VGND 0.352955f $ **FLOATING
C4891 a_12582_2982# VGND 0.352955f $ **FLOATING
C4892 a_11142_2982# VGND 0.490744f $ **FLOATING
C4893 a_15390_3334# VGND 0.375184f $ **FLOATING
C4894 a_13950_3334# VGND 0.352694f $ **FLOATING
C4895 a_12582_3334# VGND 0.352694f $ **FLOATING
C4896 a_11142_3334# VGND 0.375184f $ **FLOATING
C4897 a_13950_3686# VGND 0.352463f $ **FLOATING
C4898 a_12582_3686# VGND 0.352463f $ **FLOATING
C4899 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND 41.6715f
C4900 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.702101f
C4901 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VGND 41.754498f
C4902 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.702101f
C4903 a_15390_4038# VGND 0.397033f $ **FLOATING
C4904 a_13950_4038# VGND 0.354407f $ **FLOATING
C4905 a_12582_4038# VGND 0.354407f $ **FLOATING
C4906 a_11142_4038# VGND 0.397033f $ **FLOATING
C4907 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A VGND 37.783802f
C4908 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.38663f
C4909 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND 0.103625f
C4910 a_13950_4390# VGND 0.352432f $ **FLOATING
C4911 a_12582_4390# VGND 0.352432f $ **FLOATING
C4912 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND 0.103625f
C4913 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.38663f
C4914 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A VGND 37.790997f
C4915 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VGND 3.12067f
C4916 a_15390_4566# VGND 0.389036f $ **FLOATING
C4917 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VGND 3.08351f
C4918 a_11142_4566# VGND 0.389036f $ **FLOATING
C4919 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VGND 0.970036f
C4920 a_13950_4742# VGND 0.352456f $ **FLOATING
C4921 a_12582_4742# VGND 0.352456f $ **FLOATING
C4922 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND 0.7964f
C4923 a_15390_4918# VGND 0.470144f $ **FLOATING
C4924 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND 0.7964f
C4925 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VGND 0.970036f
C4926 a_11142_4918# VGND 0.471715f $ **FLOATING
C4927 a_13950_5094# VGND 0.353103f $ **FLOATING
C4928 a_12582_5094# VGND 0.353103f $ **FLOATING
C4929 a_15390_5270# VGND 0.492927f $ **FLOATING
C4930 a_11142_5270# VGND 0.491356f $ **FLOATING
C4931 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND 0.596866f
C4932 a_13950_5446# VGND 0.433341f $ **FLOATING
C4933 a_12582_5446# VGND 0.433756f $ **FLOATING
C4934 a_15390_5622# VGND 0.47219f $ **FLOATING
C4935 a_16542_5974# VGND 0.09029f $ **FLOATING
C4936 a_15390_5974# VGND 0.541341f $ **FLOATING
C4937 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND 0.596866f
C4938 a_11142_5622# VGND 0.47376f $ **FLOATING
C4939 a_11142_5974# VGND 0.540186f $ **FLOATING
C4940 a_9990_5974# VGND 0.09029f $ **FLOATING
C4941 a_23922_26796# VGND 0.090673f $ **FLOATING
C4942 a_22770_26796# VGND 0.529341f $ **FLOATING
C4943 a_21402_26796# VGND 0.531659f $ **FLOATING
C4944 a_20250_26796# VGND 0.088963f $ **FLOATING
C4945 a_18882_26796# VGND 0.088807f $ **FLOATING
C4946 a_17730_26796# VGND 0.530818f $ **FLOATING
C4947 a_16362_26796# VGND 0.531974f $ **FLOATING
C4948 a_15210_26796# VGND 0.088807f $ **FLOATING
C4949 a_13842_26796# VGND 0.088807f $ **FLOATING
C4950 a_12690_26796# VGND 0.530818f $ **FLOATING
C4951 a_11322_26796# VGND 0.531974f $ **FLOATING
C4952 a_10170_26796# VGND 0.088807f $ **FLOATING
C4953 a_8802_26796# VGND 0.088807f $ **FLOATING
C4954 a_7650_26796# VGND 0.530197f $ **FLOATING
C4955 a_6282_26796# VGND 0.530964f $ **FLOATING
C4956 a_5130_26796# VGND 0.088807f $ **FLOATING
C4957 a_3762_26796# VGND 0.088807f $ **FLOATING
C4958 a_2610_26796# VGND 0.531651f $ **FLOATING
C4959 a_22770_27148# VGND 0.499848f $ **FLOATING
C4960 a_21402_27148# VGND 0.467094f $ **FLOATING
C4961 a_17730_27148# VGND 0.471477f $ **FLOATING
C4962 a_16362_27148# VGND 0.467695f $ **FLOATING
C4963 a_12690_27148# VGND 0.471477f $ **FLOATING
C4964 a_11322_27148# VGND 0.467695f $ **FLOATING
C4965 a_7650_27148# VGND 0.470234f $ **FLOATING
C4966 a_6282_27148# VGND 0.465706f $ **FLOATING
C4967 a_2610_27148# VGND 0.471688f $ **FLOATING
C4968 a_21402_27500# VGND 0.385968f $ **FLOATING
C4969 a_17730_27500# VGND 0.387712f $ **FLOATING
C4970 a_16362_27500# VGND 0.386249f $ **FLOATING
C4971 a_12690_27500# VGND 0.387712f $ **FLOATING
C4972 a_11322_27500# VGND 0.386249f $ **FLOATING
C4973 a_7650_27500# VGND 0.38671f $ **FLOATING
C4974 a_6282_27500# VGND 0.384229f $ **FLOATING
C4975 a_2610_27500# VGND 0.387692f $ **FLOATING
C4976 a_21402_27852# VGND 0.370125f $ **FLOATING
C4977 a_17730_27852# VGND 0.370785f $ **FLOATING
C4978 a_16362_27852# VGND 0.368771f $ **FLOATING
C4979 a_12690_27852# VGND 0.370785f $ **FLOATING
C4980 a_11322_27852# VGND 0.368771f $ **FLOATING
C4981 a_7650_27852# VGND 0.369543f $ **FLOATING
C4982 a_6282_27852# VGND 0.366751f $ **FLOATING
C4983 a_2610_27852# VGND 0.370525f $ **FLOATING
C4984 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND 0.506947f
C4985 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND 0.501154f
C4986 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND 0.476152f
C4987 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND 0.501154f
C4988 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND 0.476152f
C4989 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND 0.501154f
C4990 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND 0.476152f
C4991 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND 0.501154f
C4992 a_21402_28204# VGND 0.405715f $ **FLOATING
C4993 a_17730_28204# VGND 0.406253f $ **FLOATING
C4994 a_16362_28204# VGND 0.406253f $ **FLOATING
C4995 a_12690_28204# VGND 0.406253f $ **FLOATING
C4996 a_11322_28204# VGND 0.406253f $ **FLOATING
C4997 a_7650_28204# VGND 0.405102f $ **FLOATING
C4998 a_6282_28204# VGND 0.404324f $ **FLOATING
C4999 a_2610_28204# VGND 0.406084f $ **FLOATING
C5000 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND 0.609217f
C5001 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND 0.741242f
C5002 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND 0.749084f
C5003 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND 0.735365f
C5004 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND 0.749084f
C5005 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND 0.735365f
C5006 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND 0.746424f
C5007 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND 0.730432f
C5008 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND 0.749031f
C5009 a_22770_28556# VGND 0.401649f $ **FLOATING
C5010 a_21402_28556# VGND 0.387558f $ **FLOATING
C5011 a_17730_28556# VGND 0.388096f $ **FLOATING
C5012 a_16362_28556# VGND 0.388096f $ **FLOATING
C5013 a_12690_28556# VGND 0.388096f $ **FLOATING
C5014 a_11322_28556# VGND 0.388096f $ **FLOATING
C5015 a_7650_28556# VGND 0.386945f $ **FLOATING
C5016 a_6282_28556# VGND 0.386167f $ **FLOATING
C5017 a_2610_28556# VGND 0.387927f $ **FLOATING
C5018 a_21402_28908# VGND 0.394283f $ **FLOATING
C5019 a_17730_28908# VGND 0.394821f $ **FLOATING
C5020 a_16362_28908# VGND 0.394821f $ **FLOATING
C5021 a_12690_28908# VGND 0.394821f $ **FLOATING
C5022 a_11322_28908# VGND 0.394821f $ **FLOATING
C5023 a_7650_28908# VGND 0.39367f $ **FLOATING
C5024 a_6282_28908# VGND 0.392892f $ **FLOATING
C5025 a_2610_28908# VGND 0.394652f $ **FLOATING
C5026 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND 0.09754f
C5027 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND 0.025702f
C5028 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND 0.09754f
C5029 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND 0.09754f
C5030 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND 0.025702f
C5031 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND 0.025702f
C5032 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND 0.09754f
C5033 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND 0.09754f
C5034 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND 0.025702f
C5035 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND 0.025702f
C5036 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND 0.09754f
C5037 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND 0.09754f
C5038 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND 0.025702f
C5039 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND 0.025702f
C5040 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND 0.09754f
C5041 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND 0.025702f
C5042 SUNSAR_SAR8B_CV_0.SARP VGND 70.6156f
C5043 a_21402_29612# VGND 0.395457f $ **FLOATING
C5044 a_17730_29612# VGND 0.396085f $ **FLOATING
C5045 a_16362_29612# VGND 0.395557f $ **FLOATING
C5046 a_12690_29612# VGND 0.396085f $ **FLOATING
C5047 a_11322_29612# VGND 0.395557f $ **FLOATING
C5048 a_7650_29612# VGND 0.394934f $ **FLOATING
C5049 a_6282_29612# VGND 0.393715f $ **FLOATING
C5050 a_2610_29612# VGND 0.39591f $ **FLOATING
C5051 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318943f
C5052 a_22770_29964# VGND 0.400512f $ **FLOATING
C5053 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND 0.103281f
C5054 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N VGND 1.27143f
C5055 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND 0.056913f
C5056 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND 0.100021f
C5057 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N VGND 1.26485f
C5058 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND 0.100021f
C5059 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N VGND 1.26371f
C5060 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND 0.048787f
C5061 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND 0.048787f
C5062 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND 0.100021f
C5063 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N VGND 1.26485f
C5064 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND 0.100021f
C5065 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N VGND 1.26371f
C5066 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND 0.048787f
C5067 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND 0.048787f
C5068 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND 0.100021f
C5069 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N VGND 1.2592f
C5070 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND 0.100021f
C5071 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N VGND 1.25309f
C5072 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND 0.048787f
C5073 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND 0.048787f
C5074 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND 0.100021f
C5075 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N VGND 1.26397f
C5076 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND 0.048787f
C5077 a_21402_30316# VGND 0.401758f $ **FLOATING
C5078 a_17730_30316# VGND 0.401042f $ **FLOATING
C5079 a_16362_30316# VGND 0.401042f $ **FLOATING
C5080 a_12690_30316# VGND 0.401042f $ **FLOATING
C5081 a_11322_30316# VGND 0.401042f $ **FLOATING
C5082 a_7650_30316# VGND 0.399891f $ **FLOATING
C5083 a_6282_30316# VGND 0.399113f $ **FLOATING
C5084 a_2610_30316# VGND 0.40113f $ **FLOATING
C5085 SUNSAR_SAR8B_CV_0.XA20.CPO VGND 15.3105f
C5086 a_22770_30844# VGND 0.421853f $ **FLOATING
C5087 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND 2.24318f
C5088 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND 2.22173f
C5089 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND 2.22173f
C5090 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND 2.22173f
C5091 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND 2.22173f
C5092 SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND 2.20887f
C5093 SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND 2.19727f
C5094 SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND 2.21994f
C5095 a_21402_31196# VGND 0.4255f $ **FLOATING
C5096 a_17730_31196# VGND 0.426037f $ **FLOATING
C5097 a_16362_31196# VGND 0.426037f $ **FLOATING
C5098 a_12690_31196# VGND 0.426037f $ **FLOATING
C5099 a_11322_31196# VGND 0.426037f $ **FLOATING
C5100 a_7650_31196# VGND 0.424886f $ **FLOATING
C5101 a_6282_31196# VGND 0.424108f $ **FLOATING
C5102 a_2610_31196# VGND 0.426125f $ **FLOATING
C5103 SUNSAR_SAR8B_CV_0.XA20.CNO VGND 19.4735f
C5104 a_22770_31724# VGND 0.423601f $ **FLOATING
C5105 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.99934f
C5106 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.97905f
C5107 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.97808f
C5108 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.97905f
C5109 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.97808f
C5110 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.85563f
C5111 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.37219f
C5112 a_21402_32076# VGND 0.426091f $ **FLOATING
C5113 a_17730_32076# VGND 0.42666f $ **FLOATING
C5114 a_16362_32076# VGND 0.42666f $ **FLOATING
C5115 a_12690_32076# VGND 0.42666f $ **FLOATING
C5116 a_11322_32076# VGND 0.42666f $ **FLOATING
C5117 a_7650_32076# VGND 0.42666f $ **FLOATING
C5118 a_6282_32076# VGND 0.42666f $ **FLOATING
C5119 a_2610_32076# VGND 0.426748f $ **FLOATING
C5120 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND 1.5559f
C5121 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C5122 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND 3.1974f
C5123 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND 3.22975f
C5124 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND 3.22837f
C5125 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND 3.22975f
C5126 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND 3.22837f
C5127 SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND 3.22679f
C5128 SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND 3.22546f
C5129 SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND 3.31251f
C5130 SUNSAR_SAR8B_CV_0.XA20.XA3a.A VGND 2.68984f
C5131 a_21402_32956# VGND 0.426069f $ **FLOATING
C5132 a_17730_32956# VGND 0.426069f $ **FLOATING
C5133 a_16362_32956# VGND 0.426069f $ **FLOATING
C5134 a_12690_32956# VGND 0.426069f $ **FLOATING
C5135 a_11322_32956# VGND 0.426069f $ **FLOATING
C5136 a_7650_32956# VGND 0.426069f $ **FLOATING
C5137 a_6282_32956# VGND 0.426069f $ **FLOATING
C5138 a_2610_32956# VGND 0.426316f $ **FLOATING
C5139 SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND 2.84889f
C5140 a_22770_33132# VGND 0.403395f $ **FLOATING
C5141 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 2.99891f
C5142 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.00352f
C5143 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.00364f
C5144 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.00352f
C5145 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.00364f
C5146 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.52399f
C5147 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.7728f
C5148 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 12.070401f
C5149 a_21402_33836# VGND 0.426756f $ **FLOATING
C5150 a_17730_33836# VGND 0.426756f $ **FLOATING
C5151 a_16362_33836# VGND 0.426756f $ **FLOATING
C5152 a_12690_33836# VGND 0.426756f $ **FLOATING
C5153 a_11322_33836# VGND 0.426756f $ **FLOATING
C5154 a_7650_33836# VGND 0.426756f $ **FLOATING
C5155 a_6282_33836# VGND 0.426756f $ **FLOATING
C5156 a_2610_33836# VGND 0.42696f $ **FLOATING
C5157 SUNSAR_SAR8B_CV_0.SARN VGND 71.385f
C5158 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND 0.149691f
C5159 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND 0.515646f
C5160 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C5161 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND 0.149691f
C5162 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.7282f
C5163 a_22770_34540# VGND 0.39377f $ **FLOATING
C5164 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND 0.102f
C5165 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND 0.149691f
C5166 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 4.17485f
C5167 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND 0.149691f
C5168 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.28054f
C5169 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND 0.102f
C5170 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND 0.102f
C5171 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND 0.149691f
C5172 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.31554f
C5173 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND 0.149691f
C5174 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.67606f
C5175 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND 0.102f
C5176 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND 0.102f
C5177 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND 0.149691f
C5178 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 4.24545f
C5179 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND 0.149988f
C5180 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 10.143099f
C5181 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND 0.102f
C5182 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND 0.102f
C5183 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND 0.102353f
C5184 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 8.215441f
C5185 a_21402_34716# VGND 0.39476f $ **FLOATING
C5186 a_17730_34716# VGND 0.39476f $ **FLOATING
C5187 a_16362_34716# VGND 0.39476f $ **FLOATING
C5188 a_12690_34716# VGND 0.39476f $ **FLOATING
C5189 a_11322_34716# VGND 0.39476f $ **FLOATING
C5190 a_7650_34716# VGND 0.39476f $ **FLOATING
C5191 a_6282_34716# VGND 0.39476f $ **FLOATING
C5192 a_2610_34716# VGND 0.394847f $ **FLOATING
C5193 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND 4.75786f
C5194 a_22770_34892# VGND 0.394644f $ **FLOATING
C5195 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.67604f
C5196 SUNSAR_SAR8B_CV_0.XA7.EN VGND 4.51423f
C5197 SUNSAR_SAR8B_CV_0.XA6.EN VGND 4.46115f
C5198 SUNSAR_SAR8B_CV_0.XA5.EN VGND 4.27635f
C5199 SUNSAR_SAR8B_CV_0.XA4.EN VGND 4.50206f
C5200 SUNSAR_SAR8B_CV_0.XA3.EN VGND 4.42499f
C5201 SUNSAR_SAR8B_CV_0.XA2.EN VGND 4.44362f
C5202 SUNSAR_SAR8B_CV_0.XA1.EN VGND 4.39196f
C5203 a_21402_35068# VGND 0.389563f $ **FLOATING
C5204 a_17730_35068# VGND 0.389563f $ **FLOATING
C5205 a_16362_35068# VGND 0.389563f $ **FLOATING
C5206 a_12690_35068# VGND 0.389563f $ **FLOATING
C5207 a_11322_35068# VGND 0.389563f $ **FLOATING
C5208 a_7650_35068# VGND 0.389563f $ **FLOATING
C5209 a_6282_35068# VGND 0.389563f $ **FLOATING
C5210 a_2610_35068# VGND 0.389651f $ **FLOATING
C5211 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND 0.096791f
C5212 SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND 4.54543f
C5213 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C5214 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C5215 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C5216 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C5217 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C5218 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C5219 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557089f
C5220 a_22770_35420# VGND 0.395535f $ **FLOATING
C5221 a_21402_35420# VGND 0.389041f $ **FLOATING
C5222 a_17730_35420# VGND 0.388925f $ **FLOATING
C5223 a_16362_35420# VGND 0.389297f $ **FLOATING
C5224 a_12690_35420# VGND 0.388925f $ **FLOATING
C5225 a_11322_35420# VGND 0.389297f $ **FLOATING
C5226 a_7650_35420# VGND 0.388925f $ **FLOATING
C5227 a_6282_35420# VGND 0.389297f $ **FLOATING
C5228 a_2610_35420# VGND 0.389228f $ **FLOATING
C5229 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND 1.07774f
C5230 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND 0.112889f
C5231 SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND 1.50901f
C5232 SUNSAR_SAR8B_CV_0.XA7.XA9.B VGND 1.53168f
C5233 SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND 1.50964f
C5234 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND 0.112889f
C5235 SUNSAR_SAR8B_CV_0.XA6.XA9.B VGND 1.54335f
C5236 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND 0.112889f
C5237 SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND 1.51005f
C5238 SUNSAR_SAR8B_CV_0.XA5.XA9.B VGND 1.53305f
C5239 SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND 1.50964f
C5240 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND 0.112889f
C5241 SUNSAR_SAR8B_CV_0.XA4.XA9.B VGND 1.54335f
C5242 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND 0.112889f
C5243 SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND 1.51005f
C5244 SUNSAR_SAR8B_CV_0.XA3.XA9.B VGND 1.53305f
C5245 SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND 1.50964f
C5246 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND 0.112889f
C5247 SUNSAR_SAR8B_CV_0.XA2.XA9.B VGND 1.54335f
C5248 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND 0.112889f
C5249 SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND 1.51005f
C5250 SUNSAR_SAR8B_CV_0.XA1.XA9.B VGND 1.53305f
C5251 SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND 1.52043f
C5252 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND 0.112889f
C5253 SUNSAR_SAR8B_CV_0.XA0.XA9.B VGND 1.61547f
C5254 a_22770_35948# VGND 0.414038f $ **FLOATING
C5255 a_21402_35948# VGND 0.390722f $ **FLOATING
C5256 a_17730_35948# VGND 0.391291f $ **FLOATING
C5257 a_16362_35948# VGND 0.391291f $ **FLOATING
C5258 a_12690_35948# VGND 0.391291f $ **FLOATING
C5259 a_11322_35948# VGND 0.391291f $ **FLOATING
C5260 a_7650_35948# VGND 0.391291f $ **FLOATING
C5261 a_6282_35948# VGND 0.391291f $ **FLOATING
C5262 a_2610_35948# VGND 0.391539f $ **FLOATING
C5263 SUNSAR_SAR8B_CV_0.XA20.XA12.Y VGND 0.79133f
C5264 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C5265 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C5266 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C5267 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C5268 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C5269 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C5270 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C5271 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.896463f
C5272 a_22770_36300# VGND 0.472701f $ **FLOATING
C5273 a_21402_36300# VGND 0.393831f $ **FLOATING
C5274 a_17730_36300# VGND 0.394738f $ **FLOATING
C5275 a_16362_36300# VGND 0.3944f $ **FLOATING
C5276 a_12690_36300# VGND 0.394718f $ **FLOATING
C5277 a_11322_36300# VGND 0.3944f $ **FLOATING
C5278 a_7650_36300# VGND 0.394715f $ **FLOATING
C5279 a_6282_36300# VGND 0.3944f $ **FLOATING
C5280 a_2610_36300# VGND 0.394963f $ **FLOATING
C5281 a_23922_36652# VGND 0.092794f $ **FLOATING
C5282 a_22770_36652# VGND 0.542519f $ **FLOATING
C5283 SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND 0.882078f
C5284 SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND 0.885089f
C5285 SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND 0.877233f
C5286 SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND 0.885067f
C5287 SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND 0.877221f
C5288 SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND 0.885066f
C5289 SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND 0.877233f
C5290 SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND 0.894319f
C5291 SUNSAR_SAR8B_CV_0.XB2.TIE_L VGND 30.566f
C5292 a_21402_36828# VGND 0.414394f $ **FLOATING
C5293 a_17730_36828# VGND 0.414304f $ **FLOATING
C5294 a_16362_36828# VGND 0.414011f $ **FLOATING
C5295 a_12690_36828# VGND 0.414294f $ **FLOATING
C5296 a_11322_36828# VGND 0.414011f $ **FLOATING
C5297 a_7650_36828# VGND 0.414296f $ **FLOATING
C5298 a_6282_36828# VGND 0.414011f $ **FLOATING
C5299 a_2610_36828# VGND 0.414386f $ **FLOATING
C5300 SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND 1.08827f
C5301 SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND 2.06522f
C5302 SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND 1.11123f
C5303 SUNSAR_SAR8B_CV_0.XA7.CEIN VGND 1.46079f
C5304 SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND 1.07013f
C5305 SUNSAR_SAR8B_CV_0.XA6.CEIN VGND 1.71822f
C5306 SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND 1.11118f
C5307 SUNSAR_SAR8B_CV_0.XA5.CEIN VGND 1.53183f
C5308 SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND 1.07013f
C5309 SUNSAR_SAR8B_CV_0.XA4.CEIN VGND 1.7182f
C5310 SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND 1.11119f
C5311 SUNSAR_SAR8B_CV_0.XA3.CEIN VGND 1.53184f
C5312 SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND 1.07013f
C5313 SUNSAR_SAR8B_CV_0.XA2.CEIN VGND 1.7182f
C5314 SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND 1.12334f
C5315 SUNSAR_SAR8B_CV_0.XA1.CEIN VGND 1.53659f
C5316 a_21402_37180# VGND 0.475717f $ **FLOATING
C5317 a_17730_37180# VGND 0.475516f $ **FLOATING
C5318 a_16362_37180# VGND 0.477063f $ **FLOATING
C5319 a_12690_37180# VGND 0.475497f $ **FLOATING
C5320 a_11322_37180# VGND 0.477061f $ **FLOATING
C5321 a_7650_37180# VGND 0.475501f $ **FLOATING
C5322 a_6282_37180# VGND 0.477063f $ **FLOATING
C5323 a_2610_37180# VGND 0.475473f $ **FLOATING
C5324 a_21402_37532# VGND 0.547813f $ **FLOATING
C5325 a_20250_37532# VGND 0.09709f $ **FLOATING
C5326 a_18882_37532# VGND 0.097424f $ **FLOATING
C5327 a_17730_37532# VGND 0.55015f $ **FLOATING
C5328 a_16362_37532# VGND 0.548796f $ **FLOATING
C5329 a_15210_37532# VGND 0.097424f $ **FLOATING
C5330 a_13842_37532# VGND 0.097424f $ **FLOATING
C5331 a_12690_37532# VGND 0.549979f $ **FLOATING
C5332 a_11322_37532# VGND 0.548796f $ **FLOATING
C5333 a_10170_37532# VGND 0.097424f $ **FLOATING
C5334 a_8802_37532# VGND 0.097424f $ **FLOATING
C5335 a_7650_37532# VGND 0.550021f $ **FLOATING
C5336 a_6282_37532# VGND 0.548798f $ **FLOATING
C5337 a_5130_37532# VGND 0.097424f $ **FLOATING
C5338 a_3762_37532# VGND 0.097737f $ **FLOATING
C5339 a_2610_37532# VGND 0.548506f $ **FLOATING
C5340 a_28727_39955# VGND 0.090364f $ **FLOATING
C5341 a_27575_39955# VGND 0.440387f $ **FLOATING
C5342 a_27575_40307# VGND 0.408627f $ **FLOATING
C5343 tt_um_TT06_SAR_done_0.x3.MP1.G VGND 1.07773f
C5344 a_27575_40659# VGND 0.389133f $ **FLOATING
C5345 tt_um_TT06_SAR_done_0.x4.MP0.G VGND 0.822801f
C5346 a_23942_40296# VGND 0.09752f $ **FLOATING
C5347 a_22790_40296# VGND 0.546732f $ **FLOATING
C5348 a_21422_40296# VGND 0.54563f $ **FLOATING
C5349 a_20270_40296# VGND 0.096349f $ **FLOATING
C5350 a_18902_40296# VGND 0.096349f $ **FLOATING
C5351 a_17750_40296# VGND 0.546813f $ **FLOATING
C5352 a_16382_40296# VGND 0.547966f $ **FLOATING
C5353 a_15230_40296# VGND 0.096349f $ **FLOATING
C5354 a_13862_40296# VGND 0.096349f $ **FLOATING
C5355 a_12710_40296# VGND 0.546813f $ **FLOATING
C5356 a_11342_40296# VGND 0.547969f $ **FLOATING
C5357 a_10190_40296# VGND 0.096349f $ **FLOATING
C5358 a_8822_40296# VGND 0.096349f $ **FLOATING
C5359 a_7670_40296# VGND 0.54681f $ **FLOATING
C5360 a_6302_40296# VGND 0.547966f $ **FLOATING
C5361 a_5150_40296# VGND 0.096349f $ **FLOATING
C5362 a_3782_40296# VGND 0.096349f $ **FLOATING
C5363 a_2630_40296# VGND 0.54539f $ **FLOATING
C5364 a_22790_40648# VGND 0.492438f $ **FLOATING
C5365 a_21422_40648# VGND 0.49034f $ **FLOATING
C5366 a_17750_40648# VGND 0.492453f $ **FLOATING
C5367 a_16382_40648# VGND 0.490883f $ **FLOATING
C5368 a_12710_40648# VGND 0.492453f $ **FLOATING
C5369 a_11342_40648# VGND 0.490883f $ **FLOATING
C5370 a_7670_40648# VGND 0.492453f $ **FLOATING
C5371 a_6302_40648# VGND 0.490883f $ **FLOATING
C5372 a_2630_40648# VGND 0.492826f $ **FLOATING
C5373 a_27575_41011# VGND 0.472817f $ **FLOATING
C5374 tt_um_TT06_SAR_done_0.DONE VGND 22.5544f
C5375 a_22790_41000# VGND 0.388777f $ **FLOATING
C5376 a_21422_41000# VGND 0.388174f $ **FLOATING
C5377 a_17750_41000# VGND 0.388174f $ **FLOATING
C5378 a_16382_41000# VGND 0.388174f $ **FLOATING
C5379 a_12710_41000# VGND 0.388174f $ **FLOATING
C5380 a_11342_41000# VGND 0.388174f $ **FLOATING
C5381 a_7670_41000# VGND 0.388174f $ **FLOATING
C5382 a_6302_41000# VGND 0.388174f $ **FLOATING
C5383 a_2630_41000# VGND 0.388638f $ **FLOATING
C5384 a_28727_41363# VGND 0.090304f $ **FLOATING
C5385 a_27575_41363# VGND 0.532318f $ **FLOATING
C5386 a_22790_41352# VGND 0.374594f $ **FLOATING
C5387 a_21422_41352# VGND 0.393558f $ **FLOATING
C5388 a_17750_41352# VGND 0.393558f $ **FLOATING
C5389 a_16382_41352# VGND 0.393558f $ **FLOATING
C5390 a_12710_41352# VGND 0.393558f $ **FLOATING
C5391 a_11342_41352# VGND 0.393558f $ **FLOATING
C5392 a_7670_41352# VGND 0.393558f $ **FLOATING
C5393 a_6302_41352# VGND 0.393558f $ **FLOATING
C5394 a_2630_41352# VGND 0.394022f $ **FLOATING
C5395 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND 0.803097f
C5396 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND 0.107737f
C5397 SUNSAR_SAR8B_CV_0.D<0> VGND 5.90005f
C5398 SUNSAR_SAR8B_CV_0.D<1> VGND 13.8814f
C5399 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND 0.107643f
C5400 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND 0.107643f
C5401 SUNSAR_SAR8B_CV_0.D<2> VGND 12.6887f
C5402 SUNSAR_SAR8B_CV_0.D<3> VGND 11.534699f
C5403 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND 0.107643f
C5404 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND 0.107643f
C5405 SUNSAR_SAR8B_CV_0.D<4> VGND 11.933901f
C5406 SUNSAR_SAR8B_CV_0.D<5> VGND 12.816799f
C5407 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND 0.107643f
C5408 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND 0.107643f
C5409 SUNSAR_SAR8B_CV_0.D<6> VGND 12.1313f
C5410 SUNSAR_SAR8B_CV_0.D<7> VGND 17.8451f
C5411 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND 0.107643f
C5412 a_22790_41880# VGND 0.394408f $ **FLOATING
C5413 a_21422_41880# VGND 0.395138f $ **FLOATING
C5414 a_17750_41880# VGND 0.395707f $ **FLOATING
C5415 a_16382_41880# VGND 0.395707f $ **FLOATING
C5416 a_12710_41880# VGND 0.395707f $ **FLOATING
C5417 a_11342_41880# VGND 0.395707f $ **FLOATING
C5418 a_7670_41880# VGND 0.395707f $ **FLOATING
C5419 a_6302_41880# VGND 0.395707f $ **FLOATING
C5420 a_2630_41880# VGND 0.396052f $ **FLOATING
C5421 SUNSAR_CAPT8B_CV_0.XA5.B VGND 1.95346f
C5422 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S VGND 0.097545f
C5423 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S VGND 0.097545f
C5424 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S VGND 0.097545f
C5425 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S VGND 0.097545f
C5426 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S VGND 0.097545f
C5427 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S VGND 0.097545f
C5428 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S VGND 0.097545f
C5429 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S VGND 0.097545f
C5430 a_22790_42408# VGND 0.410698f $ **FLOATING
C5431 a_21422_42408# VGND 0.389697f $ **FLOATING
C5432 a_17750_42408# VGND 0.390266f $ **FLOATING
C5433 a_16382_42408# VGND 0.390266f $ **FLOATING
C5434 a_12710_42408# VGND 0.390266f $ **FLOATING
C5435 a_11342_42408# VGND 0.390266f $ **FLOATING
C5436 a_7670_42408# VGND 0.390266f $ **FLOATING
C5437 a_6302_42408# VGND 0.390266f $ **FLOATING
C5438 a_2630_42408# VGND 0.390612f $ **FLOATING
C5439 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C5440 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND 1.28758f
C5441 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND 1.27933f
C5442 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND 1.27933f
C5443 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND 1.27933f
C5444 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND 1.27933f
C5445 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND 1.27933f
C5446 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND 1.27933f
C5447 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND 1.29578f
C5448 a_22790_42760# VGND 0.378208f $ **FLOATING
C5449 a_21422_42760# VGND 0.393027f $ **FLOATING
C5450 a_17750_42760# VGND 0.393596f $ **FLOATING
C5451 a_16382_42760# VGND 0.393596f $ **FLOATING
C5452 a_12710_42760# VGND 0.393596f $ **FLOATING
C5453 a_11342_42760# VGND 0.393596f $ **FLOATING
C5454 a_7670_42760# VGND 0.393596f $ **FLOATING
C5455 a_6302_42760# VGND 0.393596f $ **FLOATING
C5456 a_2630_42760# VGND 0.393942f $ **FLOATING
C5457 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 23.7501f
C5458 SUNSAR_SAR8B_CV_0.EN VGND 10.7275f
C5459 a_22790_43112# VGND 0.388427f $ **FLOATING
C5460 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S VGND 0.098268f
C5461 SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND 1.29446f
C5462 SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND 1.29655f
C5463 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S VGND 0.098268f
C5464 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S VGND 0.098268f
C5465 SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND 1.29655f
C5466 SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND 1.29655f
C5467 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S VGND 0.098268f
C5468 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S VGND 0.098268f
C5469 SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND 1.29655f
C5470 SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND 1.29655f
C5471 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S VGND 0.098268f
C5472 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S VGND 0.098268f
C5473 SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND 1.29655f
C5474 SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND 1.29893f
C5475 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S VGND 0.098268f
C5476 SUNSAR_CAPT8B_CV_0.XA6.A VGND 2.38038f
C5477 a_21422_43288# VGND 0.394124f $ **FLOATING
C5478 a_17750_43288# VGND 0.394693f $ **FLOATING
C5479 a_16382_43288# VGND 0.394693f $ **FLOATING
C5480 a_12710_43288# VGND 0.394693f $ **FLOATING
C5481 a_11342_43288# VGND 0.394693f $ **FLOATING
C5482 a_7670_43288# VGND 0.394693f $ **FLOATING
C5483 a_6302_43288# VGND 0.394693f $ **FLOATING
C5484 a_2630_43288# VGND 0.395039f $ **FLOATING
C5485 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND 0.103608f
C5486 SUNSAR_CAPT8B_CV_0.XA6.B VGND 1.64884f
C5487 a_22790_43640# VGND 0.387806f $ **FLOATING
C5488 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND 0.112889f
C5489 SUNSAR_CAPT8B_CV_0.XI14.XA7.C VGND 2.58298f
C5490 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN VGND 1.69058f
C5491 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND 0.112889f
C5492 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN VGND 1.69315f
C5493 SUNSAR_CAPT8B_CV_0.XH13.XA7.C VGND 2.56583f
C5494 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND 0.112889f
C5495 SUNSAR_CAPT8B_CV_0.XG12.XA7.C VGND 2.61645f
C5496 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN VGND 1.69315f
C5497 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND 0.112889f
C5498 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN VGND 1.69315f
C5499 SUNSAR_CAPT8B_CV_0.XF11.XA7.C VGND 2.61645f
C5500 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND 0.112889f
C5501 SUNSAR_CAPT8B_CV_0.XE10.XA7.C VGND 2.5725f
C5502 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN VGND 1.69797f
C5503 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND 0.112889f
C5504 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN VGND 1.69797f
C5505 SUNSAR_CAPT8B_CV_0.XD09.XA7.C VGND 2.5725f
C5506 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND 0.112889f
C5507 SUNSAR_CAPT8B_CV_0.XC08.XA7.C VGND 2.61716f
C5508 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN VGND 1.69797f
C5509 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND 0.112889f
C5510 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN VGND 1.69726f
C5511 SUNSAR_CAPT8B_CV_0.XB07.XA7.C VGND 2.68306f
C5512 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.88269f
C5513 a_21422_43816# VGND 0.390629f $ **FLOATING
C5514 a_17750_43816# VGND 0.391198f $ **FLOATING
C5515 a_16382_43816# VGND 0.391198f $ **FLOATING
C5516 a_12710_43816# VGND 0.391198f $ **FLOATING
C5517 a_11342_43816# VGND 0.391198f $ **FLOATING
C5518 a_7670_43816# VGND 0.391198f $ **FLOATING
C5519 a_6302_43816# VGND 0.391198f $ **FLOATING
C5520 a_2630_43816# VGND 0.391544f $ **FLOATING
C5521 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 26.3388f
C5522 a_22790_43992# VGND 0.384235f $ **FLOATING
C5523 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.23582f
C5524 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.23517f
C5525 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.23517f
C5526 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.23517f
C5527 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26123f
C5528 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C5529 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C5530 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C5531 SUNSAR_CAPT8B_CV_0.XA7.MP0.G VGND 0.5774f
C5532 a_21422_44168# VGND 0.425534f $ **FLOATING
C5533 a_20270_44168# VGND 0.088963f $ **FLOATING
C5534 a_18902_44168# VGND 0.088963f $ **FLOATING
C5535 a_17750_44168# VGND 0.425449f $ **FLOATING
C5536 a_16382_44168# VGND 0.425864f $ **FLOATING
C5537 a_15230_44168# VGND 0.088963f $ **FLOATING
C5538 a_13862_44168# VGND 0.088963f $ **FLOATING
C5539 a_12710_44168# VGND 0.425449f $ **FLOATING
C5540 a_11342_44168# VGND 0.425864f $ **FLOATING
C5541 a_10190_44168# VGND 0.088963f $ **FLOATING
C5542 a_8822_44168# VGND 0.088963f $ **FLOATING
C5543 a_7670_44168# VGND 0.425449f $ **FLOATING
C5544 a_6302_44168# VGND 0.425864f $ **FLOATING
C5545 a_5150_44168# VGND 0.088963f $ **FLOATING
C5546 a_3782_44168# VGND 0.088963f $ **FLOATING
C5547 a_2630_44168# VGND 0.426034f $ **FLOATING
C5548 TIE_L VGND 6.36945f
C5549 a_23942_44344# VGND 0.090134f $ **FLOATING
C5550 a_22790_44344# VGND 0.423601f $ **FLOATING
.ends

