* NGSPICE file created from tt_um_TT06_SAR_wulffern.ext - technology: sky130A

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt tt_um_TT06_SAR_wulffern VPWR VGND ui_in[7] ui_in[6] ui_in[5] ui_in[4] ui_in[3] ui_in[2] ui_in[1] ui_in[0]
+ uo_out[7] uo_out[6] uo_out[5] uo_out[4] uo_out[3] uo_out[2] uo_out[1] uo_out[0] uio_in[7] uio_in[6] uio_in[5] uio_in[4] uio_in[3] uio_in[2] uio_in[1] uio_in[0]
+ uio_out[7] uio_out[6] uio_out[5] uio_out[4] uio_out[3] uio_out[2] uio_out[1] uio_out[0] uio_oe[7] uio_oe[6] uio_oe[5] uio_oe[4] uio_oe[3] uio_oe[2] uio_oe[1] uio_oe[0] ua[7] ua[6] ua[5] ua[4] ua[3] ua[2] ua[1] ua[0]
+ ena clk rst_n
*.subckt tt_um_TT06_SAR_wulffern ena rst_n ua[2] ua[3] ua[4] ua[5] ua[6] ua[7]
*+ ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1]
*+ uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[1] uio_oe[2]
*+ uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[1] uio_out[2] uio_out[3]
*+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[7] uio_oe[0] ui_in[0]
*+ uo_out[6] uo_out[4] ua[0] uo_out[5] clk uo_out[1] ua[1] uo_out[0] uo_out[3] uio_out[0]
*+ VPWR VGND
X0 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA0.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X3 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X4 VGND SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X5 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.359999 w=1.08 l=0.18
X6 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R0 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X8 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X11 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X12 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X14 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X15 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R1 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X16 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=243.93959 ps=1.2855k w=1.08 l=0.18
X17 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X18 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=247.698 ps=1.29678k w=1.08 l=0.18
X19 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X20 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X21 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 VGND clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X24 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X25 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X26 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X28 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X29 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X30 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X31 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X32 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X34 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X35 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X36 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S SUNSAR_CAPT8B_CV_0.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X37 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X38 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X39 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X40 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X41 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R2 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X42 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X43 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X44 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X45 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X46 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X47 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R3 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X48 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R4 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X49 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X50 VPWR tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X51 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X52 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X53 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X54 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X55 SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X56 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X57 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=4.536 ps=21.359999 w=1.08 l=0.18
X58 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X59 SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X60 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X61 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R5 uio_out[3] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X62 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X63 SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X64 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X65 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R6 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X66 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X67 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X68 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X69 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X70 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X71 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X72 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X73 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X74 SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X75 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X76 VGND SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X77 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X78 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X79 SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X80 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X81 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S uo_out[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X82 SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X83 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X84 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X85 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X86 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R7 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X87 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X88 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X89 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X90 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X91 SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X92 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X93 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X94 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X95 VGND SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X96 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X97 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X98 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X99 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R8 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_4848# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X100 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X101 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA3.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X102 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X103 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X104 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X105 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X106 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X107 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X108 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R9 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X109 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X110 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X111 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X112 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X113 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X114 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CNO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X115 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X116 SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA1.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X117 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X118 VGND SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X119 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X120 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X121 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X122 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X123 SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X124 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R10 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X125 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X126 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X127 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X128 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X129 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X130 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X131 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X132 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X133 SUNSAR_SAR8B_CV_0.XA0.XA10.A SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X134 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X135 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X136 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X137 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CNO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X138 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X139 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R11 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X140 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X141 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X142 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X143 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X144 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X145 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X146 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X147 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X148 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X149 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X150 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X151 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X152 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X153 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X154 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X155 SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X156 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X157 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X158 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X159 SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X160 SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X161 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X162 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X163 VGND SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X164 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X165 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X166 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X167 SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X168 VPWR SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R12 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B SUNSAR_SAR8B_CV_0.D<3> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X169 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X170 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X171 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X172 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X173 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X174 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X175 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X176 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X177 VGND SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R13 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R14 uio_oe[2] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X178 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X179 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X180 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X181 SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X182 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X183 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X184 VPWR SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X185 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X186 ua[1] SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X187 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X188 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X189 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA1.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X190 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X191 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X192 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R15 uio_oe[4] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X193 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X194 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X195 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X196 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X197 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X198 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X199 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X200 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R16 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X201 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X202 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X203 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X204 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X205 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X206 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X207 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X208 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X209 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X210 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X211 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X212 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X213 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X214 VGND SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X215 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X216 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X217 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X218 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X219 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X220 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X221 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R17 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_2768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X222 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X223 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R18 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X224 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X225 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X226 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X227 SUNSAR_SAR8B_CV_0.XA3.XA12.A SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X228 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X229 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X230 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X231 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X232 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X233 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X234 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X235 SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X236 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X237 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X238 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X239 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X240 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X241 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X242 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X243 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X244 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X245 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X246 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X247 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X248 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X249 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X250 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X251 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X252 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R19 uio_out[5] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X253 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X254 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X255 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X256 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X257 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X258 SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X259 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X260 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X261 SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XE10.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X262 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X263 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X264 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S uo_out[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X265 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X266 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<2> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X267 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X268 SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X269 VPWR SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X270 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X271 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X272 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X273 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X274 SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X275 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X276 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X277 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X278 uio_oe[0] tt_um_TT06_SAR_done_0.x4.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X279 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R20 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X280 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X281 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X282 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X283 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X284 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X285 SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R21 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X286 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X287 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X289 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X290 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X291 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X292 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X293 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R22 m3_2358_6608# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X294 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X295 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X296 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X297 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X298 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X299 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X300 uio_out[0] tt_um_TT06_SAR_done_0.x3.MP1.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X301 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA2.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X302 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X303 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X304 VPWR SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X305 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X306 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X307 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X308 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X309 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X310 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X311 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X312 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X313 VPWR SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA2.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X314 VGND SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X315 SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA6.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X316 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X317 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X318 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X319 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X320 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R23 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X321 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X322 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X323 SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<1> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R24 uio_out[4] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X324 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X325 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X326 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X327 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X328 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X329 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X330 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X331 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X332 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R25 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R26 uio_out[6] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X333 SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X334 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X335 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X336 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X337 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X338 VGND SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R27 uio_out[7] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X339 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X340 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X341 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R28 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R29 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_2928# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X342 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X343 SUNSAR_SAR8B_CV_0.XA5.CEIN SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X344 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X345 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X346 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X347 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X348 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R30 uio_oe[1] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X349 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X350 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X351 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X352 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X353 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X354 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X355 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<4> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X356 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X357 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X358 SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X359 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X360 SUNSAR_CAPT8B_CV_0.XI14.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X361 VGND SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X362 SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X363 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X364 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X365 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X366 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X367 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA6.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X368 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X369 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X370 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X371 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<1> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X372 VGND SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X373 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R31 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X374 SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X375 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X376 VPWR SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X377 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X378 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X379 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X380 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X381 SUNSAR_SAR8B_CV_0.XA6.XA11.A SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X382 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X383 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X384 SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S uo_out[5] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X385 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X386 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
R32 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X387 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X388 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X389 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X390 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X391 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X392 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X393 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R33 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.D<4> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X394 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X395 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X396 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X397 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X398 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X399 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X400 VPWR SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X401 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R34 uio_oe[5] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X402 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X403 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X404 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X405 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X406 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X407 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X408 SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA4.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X409 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X410 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X411 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X412 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R35 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X413 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X414 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X415 VGND SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X416 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X417 SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<3> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X418 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X419 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X420 SUNSAR_SAR8B_CV_0.XA20.XA11.Y tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X421 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X422 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R36 uio_out[1] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X423 uo_out[6] SUNSAR_CAPT8B_CV_0.XC08.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X424 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X425 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X426 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X427 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X428 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X429 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X430 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X431 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X432 VGND SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X433 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X434 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X435 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R37 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_5648# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X436 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X437 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X438 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X439 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R38 uio_oe[3] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X440 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R39 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X441 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X442 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X443 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X444 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X445 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X446 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.D<7> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R40 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X447 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X448 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X449 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X450 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X451 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X452 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X453 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X454 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X455 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X456 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X457 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA4.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X458 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X459 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X460 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X461 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X462 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X463 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<3> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X464 VPWR SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X465 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X466 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X467 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X468 SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S uo_out[7] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X469 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X470 SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X471 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X472 uo_out[0] SUNSAR_CAPT8B_CV_0.XI14.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X473 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X474 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X475 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X476 VGND SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R41 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X477 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X478 SUNSAR_CAPT8B_CV_0.XD09.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X479 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X480 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X481 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R42 m3_2358_4688# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X482 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X483 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X484 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X485 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X486 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X487 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X488 VGND SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X489 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X490 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X491 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X492 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X493 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X494 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X495 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X496 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X497 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X498 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X499 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X500 VPWR SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X501 VGND SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R43 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X502 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X503 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X504 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X505 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R44 uio_out[2] TIE_L1 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X506 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X507 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X508 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X509 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X510 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R45 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X511 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X512 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X513 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X514 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X515 SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA5.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X516 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X517 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X518 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X519 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X520 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X521 VGND SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X522 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X523 SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<2> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X524 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X525 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X526 SUNSAR_SAR8B_CV_0.XA20.CK_CMP SUNSAR_SAR8B_CV_0.XA7.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X527 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X528 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X529 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X530 SUNSAR_SAR8B_CV_0.XA4.XA10.A SUNSAR_SAR8B_CV_0.XA4.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X531 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XA5.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R46 uio_oe[6] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X532 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X533 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X534 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X535 SUNSAR_CAPT8B_CV_0.XB07.QN SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X536 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X537 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X538 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X539 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X540 SUNSAR_CAPT8B_CV_0.XI14.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X541 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X542 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X543 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R47 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X544 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R48 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_5808# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X545 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X546 SUNSAR_SAR8B_CV_0.XA20.XA10.MN1.S SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X547 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X548 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X549 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X550 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X551 SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X552 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X553 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X554 SUNSAR_SAR8B_CV_0.XA4.XA9.A SUNSAR_SAR8B_CV_0.XA5.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X555 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X556 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X557 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X558 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X559 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X560 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X561 VGND SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X562 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X563 SUNSAR_CAPT8B_CV_0.XB07.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X564 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X565 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X566 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X567 VPWR SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X568 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X569 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S uo_out[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X570 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X571 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X572 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X573 SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S uo_out[6] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X574 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X575 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X576 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X577 SUNSAR_CAPT8B_CV_0.XA2.MP0.G SUNSAR_CAPT8B_CV_0.XA2.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X578 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X579 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X580 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X581 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
R49 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X582 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X583 ua[1] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X584 SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S SUNSAR_CAPT8B_CV_0.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X585 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X586 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA5.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X587 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X588 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X589 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X590 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X591 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X592 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X593 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X594 SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA3.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X595 VGND SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R50 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X596 VGND SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X597 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X598 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X599 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.D<0> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X600 VGND SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X601 SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X602 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X603 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X604 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X605 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X606 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X607 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X608 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R51 TIE_L2 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X609 VGND SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X610 VGND SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X611 SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XA3.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X612 VGND SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X613 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X614 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X615 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X616 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X617 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X618 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X619 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X620 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X621 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X622 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X623 SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X624 SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S uo_out[0] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X625 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X626 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X627 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X628 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X629 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X630 SUNSAR_SAR8B_CV_0.XA5.XA10.A SUNSAR_SAR8B_CV_0.XA5.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X631 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X632 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<0> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X633 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X634 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X635 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X636 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X637 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X638 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X639 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X640 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X641 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X642 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X643 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X644 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R52 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X645 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X646 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X647 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X648 SUNSAR_SAR8B_CV_0.XA7.XA6.MP1.S SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X649 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X650 SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XD09.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X651 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X652 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X653 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R53 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X654 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X655 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X656 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X657 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X658 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X659 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X660 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X661 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X662 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X663 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X664 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X665 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X666 SUNSAR_CAPT8B_CV_0.XC08.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R54 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R55 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X667 SUNSAR_CAPT8B_CV_0.XC08.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R56 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_3728# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X668 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X669 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X670 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X671 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X672 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X673 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X674 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X675 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X676 VPWR clk SUNSAR_CAPT8B_CV_0.XA4.MP1.G VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X677 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X678 VGND SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X679 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X680 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X681 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X682 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X683 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X684 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X685 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X686 VPWR SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X687 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X688 VPWR VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X689 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X690 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X691 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X692 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X693 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X694 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X695 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.B VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R57 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X696 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X697 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X698 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X699 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X700 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X701 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X702 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X703 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X704 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X705 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X706 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R58 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X707 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X708 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X709 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X710 VGND tt_um_TT06_SAR_done_0.DONE tt_um_TT06_SAR_done_0.x3.MP1.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X711 SUNSAR_CAPT8B_CV_0.XI14.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X712 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X713 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X714 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X715 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X716 SUNSAR_CAPT8B_CV_0.XA6.XA2.A SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X717 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R59 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X718 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X719 SUNSAR_CAPT8B_CV_0.XG12.QN SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X720 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R60 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_3888# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X721 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X722 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X723 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X724 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X725 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X726 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R61 VGND SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X727 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X728 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X729 VGND SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X730 VGND SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X731 SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X732 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA6.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X733 VPWR SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X734 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X735 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X736 SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X737 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X738 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X739 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X740 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X741 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X742 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X743 SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X744 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X745 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X746 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X747 ua[0] SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X748 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X749 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X750 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R62 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X751 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X752 SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X753 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R63 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X754 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X755 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X756 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S uo_out[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X757 SUNSAR_SAR8B_CV_0.XA2.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X758 VGND SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X759 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R64 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X760 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X761 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X762 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X763 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X764 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X765 SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S uo_out[1] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X766 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X767 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X768 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X769 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CNO VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R65 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.D<1> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X770 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X771 VGND SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X772 VGND SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X773 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X774 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X775 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA4.EN VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X776 VPWR SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X777 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X778 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X779 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X780 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X781 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X782 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CNO VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X783 VGND SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X784 SUNSAR_SAR8B_CV_0.XA1.XA12.A SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X785 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X786 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X787 SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R66 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X788 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X789 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X790 VPWR SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X791 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X792 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X793 VGND SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X794 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X795 uo_out[2] SUNSAR_CAPT8B_CV_0.XG12.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X796 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X797 SUNSAR_SAR8B_CV_0.XA7.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X798 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X799 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X800 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.D<1> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X801 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X802 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X803 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X804 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X805 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X806 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X807 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X808 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X809 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X810 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X811 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X812 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XA4.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X813 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X814 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X815 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X816 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MN1.S SUNSAR_SAR8B_CV_0.XA20.CPO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X817 SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X818 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X819 SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<7> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X820 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X821 VGND SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X822 SUNSAR_CAPT8B_CV_0.XC08.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X823 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X824 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X825 SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XC08.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X826 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X827 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X828 SUNSAR_SAR8B_CV_0.XA2.XA9.A SUNSAR_SAR8B_CV_0.XA3.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X829 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X830 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X831 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X832 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X833 SUNSAR_SAR8B_CV_0.XA0.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X834 VPWR SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X835 ua[1] SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X836 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X837 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X838 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X839 VGND SUNSAR_SAR8B_CV_0.XA3.XA2.A SUNSAR_SAR8B_CV_0.XA3.CN1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X840 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X841 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X842 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X843 SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S uo_out[3] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
R67 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.D<2> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X844 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X845 SUNSAR_CAPT8B_CV_0.XB07.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X846 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X847 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X848 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R68 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.CP<9> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X849 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X850 SUNSAR_CAPT8B_CV_0.XH13.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X851 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X852 VGND SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X853 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X854 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X855 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R69 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_6608# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X856 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X857 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X858 SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA7.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X859 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X860 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X861 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X862 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X863 SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X864 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X865 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X866 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X867 SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X868 uo_out[5] SUNSAR_CAPT8B_CV_0.XD09.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X869 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X870 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X871 VGND SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X872 VPWR SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R70 uio_oe[7] TIE_L2 sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X873 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X874 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X875 SUNSAR_CAPT8B_CV_0.XH13.XA6.A SUNSAR_CAPT8B_CV_0.XH13.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X876 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X877 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X878 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X879 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X880 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X881 VGND SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X882 SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XI14.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X883 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X884 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X885 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X886 VGND SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X887 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X888 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X889 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
X890 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X891 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.QN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X892 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> SUNSAR_SAR8B_CV_0.XA5.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X893 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.D<3> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X894 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X895 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X896 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X897 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X898 VGND SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X899 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.D<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X900 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X901 uo_out[1] SUNSAR_CAPT8B_CV_0.XH13.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R71 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.CP<8> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X902 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X903 VGND SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X904 SUNSAR_SAR8B_CV_0.XA1.XA10.A SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X905 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R72 m3_2358_5648# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X906 SUNSAR_CAPT8B_CV_0.XF11.QN SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X907 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X908 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X909 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X910 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R73 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R74 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_9126_6768# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X911 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X912 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X913 VGND SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X914 tt_um_TT06_SAR_done_0.x4.MP0.G tt_um_TT06_SAR_done_0.x4.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X915 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X916 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X917 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
R75 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B SUNSAR_SAR8B_CV_0.D<5> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X918 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X919 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X920 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X921 SUNSAR_SAR8B_CV_0.XA20.CPO SUNSAR_SAR8B_CV_0.XA20.XA3.CO VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X922 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X923 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S SUNSAR_SAR8B_CV_0.D<6> VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X924 SUNSAR_CAPT8B_CV_0.XI14.QN SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X925 SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<6> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X926 VPWR SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X927 VPWR VGND sky130_fd_pr__cap_mim_m3_1 l=18 w=18
X928 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X929 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X930 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X931 SUNSAR_CAPT8B_CV_0.XG12.XA5.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X932 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X933 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN2.S SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X934 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X935 SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X936 uio_out[0] tt_um_TT06_SAR_done_0.x3.MP1.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X937 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X938 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X939 SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X940 SUNSAR_CAPT8B_CV_0.XF11.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XF11.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X941 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X942 SUNSAR_SAR8B_CV_0.XA1.XA6.MP1.S SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XA1.XA9.B VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X943 VGND SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X944 SUNSAR_SAR8B_CV_0.XA4.CN1 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X945 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X946 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S uo_out[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X947 SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S uo_out[2] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X948 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R76 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
R77 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X949 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X950 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X951 SUNSAR_SAR8B_CV_0.XA0.DONE SUNSAR_SAR8B_CV_0.XA0.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X952 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X953 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X954 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X955 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X956 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X957 VPWR SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X958 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B SUNSAR_SAR8B_CV_0.XB1.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X959 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA5.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X960 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X961 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X962 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A SUNSAR_SAR8B_CV_0.D<7> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R78 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X963 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X964 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X965 VGND SUNSAR_SAR8B_CV_0.XB2.TIE_L SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X966 SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S SUNSAR_SAR8B_CV_0.XA2.XA11.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X967 VGND SUNSAR_SAR8B_CV_0.XA6.XA4.A SUNSAR_SAR8B_CV_0.XA6.CP0 VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X968 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X969 TIE_L SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X970 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.XA6.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X971 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X972 SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S SUNSAR_SAR8B_CV_0.D<0> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X973 SUNSAR_SAR8B_CV_0.XA6.XA12.A SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X974 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X975 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X976 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X977 SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S SUNSAR_SAR8B_CV_0.D<5> VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X978 ua[0] SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X979 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X980 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_CAPT8B_CV_0.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X981 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X982 uo_out[3] SUNSAR_CAPT8B_CV_0.XF11.QN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X983 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X984 VGND SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X985 SUNSAR_SAR8B_CV_0.XA7.CN0 SUNSAR_SAR8B_CV_0.XA7.CP0 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X986 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XA2.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X987 VGND SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X988 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X989 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X990 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X991 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X992 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X993 VGND SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<5> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R79 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B SUNSAR_SAR8B_CV_0.D<6> sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X994 SUNSAR_SAR8B_CV_0.XA2.XA2.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X995 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN SUNSAR_CAPT8B_CV_0.XI14.XA7.C VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X996 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP2.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X997 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X998 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X999 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1000 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1001 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1002 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1003 ua[0] SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1004 VPWR SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1005 VGND SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1006 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GN VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1007 VGND SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R80 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1008 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S uo_out[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1009 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1010 SUNSAR_CAPT8B_CV_0.XB07.XA4.MN1.S SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1011 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1012 SUNSAR_SAR8B_CV_0.XA3.XA10.A SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1013 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1014 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1015 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R81 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B sky130_fd_pr__res_generic_l1 w=0.34 l=0.34
X1016 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.CKN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1017 SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1018 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA4.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1019 SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S SUNSAR_CAPT8B_CV_0.XH13.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1020 VGND SUNSAR_SAR8B_CV_0.XA3.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1021 VGND SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1022 SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP2.S SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1023 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1024 VPWR SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
R82 TIE_L1 TIE_L sky130_fd_pr__res_generic_m4 w=0.3 l=0.3
X1025 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S SUNSAR_SAR8B_CV_0.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1026 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1027 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S uo_out[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1028 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1029 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1030 SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S uo_out[4] VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1031 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S SUNSAR_SAR8B_CV_0.XA20.CNO VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1032 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1033 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.ENO VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
R83 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A m3_24750_4688# sky130_fd_pr__res_generic_m3 w=0.4 l=0.36
X1034 SUNSAR_CAPT8B_CV_0.XD09.QN SUNSAR_CAPT8B_CV_0.XD09.XA7.CN SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1035 SUNSAR_CAPT8B_CV_0.XG12.XA6.MN1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1036 VGND VGND VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1037 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1038 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA9.Y VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1039 SUNSAR_CAPT8B_CV_0.XG12.XA6.MP1.S SUNSAR_CAPT8B_CV_0.XG12.XA6.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1040 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X1041 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S uo_out[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1042 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1043 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1044 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1045 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1046 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1047 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1048 SUNSAR_SAR8B_CV_0.XA1.DONE SUNSAR_SAR8B_CV_0.XA1.XA9.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1049 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1050 VGND tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.378 ps=1.78 w=1.08 l=0.18
X1051 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XA0.XA4.A VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1052 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN2.S SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.378 ps=1.78 w=1.08 l=0.18
X1053 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND VGND sky130_fd_pr__nfet_01v8 ad=0.378 pd=1.78 as=0.6156 ps=3.3 w=1.08 l=0.18
X1054 VPWR VPWR VPWR VPWR sky130_fd_pr__pfet_01v8 ad=0.378 pd=1.78 as=0 ps=0 w=1.08 l=0.18
C0 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA4.CEIN 0.432008f
C1 SUNSAR_CAPT8B_CV_0.XI14.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C2 SUNSAR_CAPT8B_CV_0.XF11.XA5.A a_12710_42408# 0.111909f
C3 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.EN 0.13041f
C4 VPWR a_8802_28556# 0.406628f
C5 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S ua[0] 0.100365f
C6 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.11641f
C7 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CP0 0.722427f
C8 a_6302_42408# SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.113479f
C9 VPWR a_20250_28204# 0.361706f
C10 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.MP1.S 0.106927f
C11 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB2.CKN 0.669708f
C12 VPWR a_23922_27148# 0.483246f
C13 VPWR SUNSAR_SAR8B_CV_0.XA2.XA6.MP3.S 0.112858f
C14 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 4.25569f
C15 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.201839f
C16 VPWR a_23942_42408# 0.3915f
C17 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN a_17750_42408# 0.100131f
C18 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 13.6519f
C19 VPWR a_5130_36300# 0.398846f
C20 VPWR a_9990_5270# 0.490626f
C21 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.924613f
C22 a_13842_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C23 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C24 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.40569f
C25 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.649845f
C26 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.MP1.S 0.119314f
C27 VPWR SUNSAR_SAR8B_CV_0.XA7.CN0 1.70987f
C28 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XA5.EN 0.11536f
C29 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.432466f
C30 VPWR a_18882_27500# 0.382189f
C31 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S ua[1] 0.100365f
C32 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C33 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.16236f
C34 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.126085f
C35 VPWR a_16542_5974# 0.449888f
C36 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.449584f
C37 VPWR a_20250_31196# 0.437f
C38 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.107427f
C39 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_7670_41000# 0.114097f
C40 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.301485f
C41 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.145483f
C42 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 3.23197f
C43 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C44 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.151329f
C45 VPWR a_15210_28908# 0.395394f
C46 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.D<1> 0.327152f
C47 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN 0.152052f
C48 VPWR a_18882_37532# 0.458364f
C49 VPWR SUNSAR_SAR8B_CV_0.D<5> 5.39172f
C50 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.CO 1.43919f
C51 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.303978f
C52 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.178114f
C53 VPWR a_15210_26796# 0.441753f
C54 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.40569f
C55 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.D<3> 0.433299f
C56 VPWR a_3762_30316# 0.404384f
C57 VPWR SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.720096f
C58 SUNSAR_CAPT8B_CV_0.XA6.A clk 0.206733f
C59 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA6.A 1.63909f
C60 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_SAR8B_CV_0.D<0> 0.393578f
C61 SUNSAR_SAR8B_CV_0.XA5.CN1 a_16362_31196# 0.109137f
C62 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.559553f
C63 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 3.86364f
C64 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA4.CEIN 0.220689f
C65 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.379175p
C66 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARP 0.187721f
C67 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.57155f
C68 VPWR a_18882_35068# 0.394528f
C69 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.112859f
C70 VPWR SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G 0.808658f
C71 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.SARN 1.62434f
C72 VPWR a_23942_43640# 0.412992f
C73 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN 0.152052f
C74 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA1.EN 0.11341f
C75 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.12241f
C76 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.D<0> 0.409858f
C77 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 0.432466f
C78 SUNSAR_SAR8B_CV_0.SARP ua[1] 1.01369f
C79 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_SAR8B_CV_0.D<3> 0.241356f
C80 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA7.CEIN 0.324105f
C81 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.204048f
C82 SUNSAR_SAR8B_CV_0.XA20.CK_CMP tt_um_TT06_SAR_done_0.DONE 0.301665f
C83 VPWR a_13842_32076# 0.436368f
C84 SUNSAR_SAR8B_CV_0.XA2.XA11.A SUNSAR_SAR8B_CV_0.XA2.CEIN 0.303978f
C85 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142977f
C86 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA4.A 0.638386f
C87 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP2.S 0.150467f
C88 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.176792f
C89 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.136678f
C90 SUNSAR_SAR8B_CV_0.XA1.XA2.A SUNSAR_SAR8B_CV_0.EN 0.166192f
C91 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.40569f
C92 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.166192f
C93 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.11884f
C94 uo_out[1] uo_out[0] 0.355472f
C95 VPWR a_10170_28204# 0.361706f
C96 a_15230_41000# SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.156079f
C97 SUNSAR_SAR8B_CV_0.XA3.XA11.A a_11322_36300# 0.13402f
C98 VPWR a_15210_27852# 0.358413f
C99 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.145048f
C100 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.158152f
C101 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.449584f
C102 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.339883f
C103 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.142061f
C104 VPWR a_18902_44168# 0.3405f
C105 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.787331f
C106 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA6.A 0.545186f
C107 VPWR a_15210_34716# 0.399819f
C108 VPWR a_23922_34892# 0.395601f
C109 a_2610_35948# SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.132671f
C110 VPWR a_18882_28556# 0.406628f
C111 VPWR a_5130_27852# 0.358413f
C112 VPWR SUNSAR_SAR8B_CV_0.XA2.XA2.A 2.45309f
C113 VPWR SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.725614f
C114 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.207877f
C115 SUNSAR_CAPT8B_CV_0.XE10.QN SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.318734f
C116 VPWR SUNSAR_SAR8B_CV_0.XA7.EN 5.54203f
C117 VPWR SUNSAR_CAPT8B_CV_0.XG12.QN 0.901622f
C118 VPWR a_15230_42408# 0.391292f
C119 VPWR a_3762_26796# 0.442908f
C120 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.29297f
C121 VPWR a_8802_36300# 0.399161f
C122 SUNSAR_SAR8B_CV_0.XA6.CN1 a_17730_31196# 0.107567f
C123 VPWR tt_um_TT06_SAR_done_0.x3.MP1.G 0.695784f
C124 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.D<4> 3.07223f
C125 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.CO 4.93712f
C126 VPWR a_15210_28556# 0.406628f
C127 VPWR SUNSAR_SAR8B_CV_0.CK_SAMPLE 9.97874f
C128 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.665179f
C129 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.CN1 0.625035f
C130 VPWR a_3762_34716# 0.399819f
C131 VPWR a_3762_27500# 0.382189f
C132 a_21402_32956# SUNSAR_SAR8B_CV_0.XA7.CP0 0.102695f
C133 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.CNO 0.108751f
C134 VPWR SUNSAR_SAR8B_CV_0.XA0.XA2.A 2.45309f
C135 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA0.DONE 0.143554f
C136 VPWR a_9990_2630# 0.447601f
C137 VPWR a_5130_35068# 0.394528f
C138 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.224309f
C139 VPWR a_5130_36828# 0.395767f
C140 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.145483f
C141 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.527529f
C142 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.CN1 0.702226f
C143 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.EN 0.849501f
C144 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.244517f
C145 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MP1.S 0.104609f
C146 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 1.7759f
C147 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.180903f
C148 VPWR a_5150_41000# 0.38821f
C149 a_16542_3334# SUNSAR_SAR8B_CV_0.XB2.CKN 0.120042f
C150 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.147435f
C151 SUNSAR_SAR8B_CV_0.XA5.EN a_12690_28556# 0.132757f
C152 VPWR SUNSAR_SAR8B_CV_0.XA20.XA10.Y 2.1352f
C153 a_7650_35068# SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.127528f
C154 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.527529f
C155 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 54.2165f
C156 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.145483f
C157 a_16362_32956# SUNSAR_SAR8B_CV_0.XA5.CP0 0.102695f
C158 VPWR a_18902_40296# 0.458821f
C159 a_23942_42760# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.101843f
C160 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_SAR8B_CV_0.D<1> 0.241356f
C161 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN a_5150_41880# 0.100592f
C162 uo_out[6] uo_out[5] 0.327382f
C163 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.79343f
C164 SUNSAR_SAR8B_CV_0.XA0.XA11.A a_2610_36300# 0.13253f
C165 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.426291f
C166 VPWR a_8802_37180# 0.473729f
C167 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> a_10170_33836# 0.101833f
C168 a_22770_34540# SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.103065f
C169 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA5.A 0.898003f
C170 VPWR a_15230_44168# 0.340085f
C171 TIE_L2 uo_out[7] 0.100011f
C172 VPWR SUNSAR_CAPT8B_CV_0.XD09.QN 0.901622f
C173 TIE_L uio_oe[0] 1.21913f
C174 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 6.86675f
C175 a_11322_35068# SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.129098f
C176 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA3.EN 0.434116f
C177 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.209352f
C178 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.432466f
C179 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.EN 0.166272f
C180 VPWR a_23942_43112# 0.393308f
C181 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 0.635098f
C182 VPWR SUNSAR_SAR8B_CV_0.XA6.XA2.A 2.44986f
C183 a_8802_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C184 VPWR a_5130_32956# 0.436368f
C185 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.250503f
C186 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XA2.XA4.A 0.227341f
C187 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.342913f
C188 VPWR SUNSAR_SAR8B_CV_0.XA7.XA2.A 2.45124f
C189 VPWR a_28727_41363# 0.440399f
C190 a_7650_35948# SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.132671f
C191 SUNSAR_CAPT8B_CV_0.XD09.XA7.C uo_out[5] 0.245678f
C192 SUNSAR_CAPT8B_CV_0.XC08.XA6.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.649845f
C193 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 1.7759f
C194 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142956f
C195 VPWR a_3762_35948# 0.417826f
C196 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.383512f
C197 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.138f
C198 SUNSAR_SAR8B_CV_0.EN SUNSAR_CAPT8B_CV_0.XA6.B 0.176398f
C199 VPWR SUNSAR_SAR8B_CV_0.XA6.CP0 2.64055f
C200 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA6.A 0.744161f
C201 VPWR a_8802_37532# 0.45854f
C202 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.ENO 0.15234f
C203 SUNSAR_SAR8B_CV_0.XA5.XA2.A a_15210_30316# 0.127528f
C204 VPWR a_18882_37180# 0.473682f
C205 VPWR SUNSAR_SAR8B_CV_0.D<3> 5.44842f
C206 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C207 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA3.MP1.S 0.106927f
C208 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.744161f
C209 VPWR a_23922_33132# 0.415713f
C210 uo_out[7] uo_out[5] 1.57818f
C211 VPWR a_13842_37532# 0.458421f
C212 SUNSAR_SAR8B_CV_0.D<6> tt_um_TT06_SAR_done_0.DONE 0.2961f
C213 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.39306f
C214 VPWR a_8822_40648# 0.491776f
C215 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.253395f
C216 VPWR a_23942_40648# 0.490244f
C217 VPWR a_13842_37180# 0.473697f
C218 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 0.419738f
C219 VPWR SUNSAR_SAR8B_CV_0.XA7.XA9.A 1.20972f
C220 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B 0.40569f
C221 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_SAR8B_CV_0.D<6> 0.241356f
C222 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 54.2165f
C223 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.199516f
C224 a_6282_35420# SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.160931f
C225 a_17750_41000# SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.114097f
C226 TIE_L1 TIE_L 0.257793f
C227 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.201839f
C228 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.649845f
C229 a_20250_30316# SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.127528f
C230 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.A 1.22023f
C231 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.12241f
C232 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.D<3> 0.228326f
C233 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA7.EN 0.144331f
C234 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.174845f
C235 VPWR a_13842_33836# 0.409601f
C236 VPWR a_23922_35420# 0.416528f
C237 VPWR a_20270_43816# 0.391817f
C238 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.MP1.S 0.106927f
C239 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.227352f
C240 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.393055f
C241 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.280191f
C242 VPWR a_3762_28204# 0.36179f
C243 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA2.CEIN 0.13078f
C244 SUNSAR_CAPT8B_CV_0.XF11.QN uo_out[3] 0.267395f
C245 VPWR a_3762_27148# 0.471462f
C246 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.118226f
C247 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA20.CPO 0.255261f
C248 SUNSAR_CAPT8B_CV_0.XB07.XA6.A a_3782_42760# 0.113305f
C249 VPWR a_13842_32956# 0.436368f
C250 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.746324f
C251 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.105541f
C252 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_SAR8B_CV_0.XA3.CP0 0.327909f
C253 SUNSAR_SAR8B_CV_0.XA20.XA11.Y tt_um_TT06_SAR_done_0.DONE 0.111867f
C254 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CP0 0.722417f
C255 VPWR a_5130_28908# 0.395394f
C256 VPWR a_20270_43288# 0.394205f
C257 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 0.635098f
C258 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA3.MP1.S 0.106927f
C259 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.133602f
C260 SUNSAR_SAR8B_CV_0.XA7.XA12.A a_21402_36828# 0.104051f
C261 VPWR SUNSAR_SAR8B_CV_0.XA5.XA2.A 2.45309f
C262 VPWR a_23922_35948# 0.390687f
C263 VPWR a_18882_35420# 0.39968f
C264 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.324243f
C265 VPWR a_15210_31196# 0.44007f
C266 a_11342_41000# SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.115667f
C267 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 3.55251f
C268 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111173f
C269 a_7670_42408# SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.100131f
C270 TIE_L1 uio_oe[0] 0.902557f
C271 VPWR SUNSAR_CAPT8B_CV_0.XH13.QN 0.901622f
C272 a_23922_29964# SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.151031f
C273 SUNSAR_SAR8B_CV_0.SARP ua[0] 0.694484f
C274 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.SARP 27.1615f
C275 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.1501f
C276 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.A 0.722887f
C277 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111173f
C278 a_2630_42408# SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.100131f
C279 VPWR a_20250_26796# 0.441753f
C280 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.276413f
C281 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C282 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_2982# 0.158066f
C283 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_21422_41000# 0.115667f
C284 a_15210_35420# SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.133834f
C285 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_SAR8B_CV_0.D<2> 0.241356f
C286 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3334# 0.163985f
C287 a_11322_35948# SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.134161f
C288 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.EN 0.3401f
C289 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.649845f
C290 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA4.MP1.S 0.104609f
C291 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.QN 0.318734f
C292 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142977f
C293 VPWR a_20250_36300# 0.395776f
C294 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B 0.419738f
C295 a_9990_3334# SUNSAR_SAR8B_CV_0.XB1.CKN 0.118471f
C296 VPWR SUNSAR_SAR8B_CV_0.XA7.XA4.A 2.30036f
C297 a_10190_41880# SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.100592f
C298 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 0.40569f
C299 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.898003f
C300 VPWR SUNSAR_SAR8B_CV_0.XA6.CN1 2.62329f
C301 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<3> 2.98135f
C302 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.CKN 0.41624f
C303 a_16362_36828# SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.104051f
C304 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA5.A 0.898003f
C305 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 3.3576f
C306 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA6.A 1.63909f
C307 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.686731f
C308 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.271482f
C309 VPWR a_28727_41011# 0.468616f
C310 SUNSAR_CAPT8B_CV_0.XE10.QN a_11342_43816# 0.129239f
C311 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.744161f
C312 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.748719f
C313 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> a_6282_31196# 0.11263f
C314 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.SARP 6.86675f
C315 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.143148f
C316 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B 3.55251f
C317 SUNSAR_CAPT8B_CV_0.XH13.XA6.A a_18902_42760# 0.113305f
C318 VPWR a_15210_27148# 0.470364f
C319 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C320 VPWR SUNSAR_SAR8B_CV_0.XA1.XA11.MP1.S 0.101979f
C321 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.A 0.725614f
C322 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.363295f
C323 SUNSAR_CAPT8B_CV_0.XI14.XA7.C uo_out[0] 0.245678f
C324 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.224309f
C325 VPWR a_10190_43288# 0.394205f
C326 VPWR a_5130_29612# 0.397362f
C327 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.CN 1.7759f
C328 SUNSAR_SAR8B_CV_0.XA6.XA10.A a_17730_35948# 0.132671f
C329 VPWR a_20250_34716# 0.396749f
C330 VPWR SUNSAR_CAPT8B_CV_0.XE10.QN 0.901622f
C331 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.C 2.97224f
C332 VPWR a_3782_40296# 0.458821f
C333 VPWR a_23922_28556# 0.499441f
C334 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.144331f
C335 VPWR a_20250_33836# 0.407174f
C336 SUNSAR_SAR8B_CV_0.CK_SAMPLE SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.106828f
C337 a_20250_29612# SUNSAR_SAR8B_CV_0.EN 0.142592f
C338 VPWR SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.784656f
C339 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA6.A 0.301485f
C340 VPWR a_20270_41000# 0.388204f
C341 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C342 VPWR SUNSAR_SAR8B_CV_0.XA3.CP0 2.64054f
C343 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA6.A 1.63909f
C344 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 6.34383f
C345 VPWR TIE_L 0.387688f
C346 VPWR SUNSAR_SAR8B_CV_0.XA2.EN 4.84607f
C347 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.EN 0.11263f
C348 a_16382_43816# SUNSAR_CAPT8B_CV_0.XG12.QN 0.129239f
C349 VPWR a_20250_36828# 0.392512f
C350 VPWR a_9990_2982# 0.491909f
C351 a_21422_43816# SUNSAR_CAPT8B_CV_0.XI14.QN 0.129239f
C352 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.EN 0.13041f
C353 VPWR SUNSAR_SAR8B_CV_0.XA5.CP0 2.64054f
C354 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.SARN 5.22744f
C355 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.SARP 54.2165f
C356 VPWR a_9990_3334# 0.380282f
C357 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 13.6519f
C358 VPWR a_20250_32956# 0.433941f
C359 VPWR a_3762_36828# 0.395857f
C360 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.204048f
C361 VPWR a_8802_27148# 0.471462f
C362 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.D<3> 0.438277f
C363 VPWR a_8802_27500# 0.382189f
C364 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.15651f
C365 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.D<4> 0.297363f
C366 VPWR a_23942_43992# 0.388156f
C367 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.GN 0.665179f
C368 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.MP1.S 0.119314f
C369 VPWR SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.779986f
C370 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.379175p
C371 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.SARP 0.524159f
C372 a_12582_4742# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.156331f
C373 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 0.63636f
C374 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.144331f
C375 VPWR a_10190_44168# 0.340085f
C376 VPWR a_8822_41000# 0.388305f
C377 SUNSAR_SAR8B_CV_0.XA7.XA9.B tt_um_TT06_SAR_done_0.DONE 0.291229f
C378 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.CPO 0.131536f
C379 VPWR a_10170_36828# 0.396003f
C380 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA20.CPO 1.15994f
C381 SUNSAR_SAR8B_CV_0.XA7.XA12.A SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.182595f
C382 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.D<4> 0.228332f
C383 VPWR a_15210_29612# 0.397362f
C384 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S 0.104122f
C385 VPWR SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 2.50679f
C386 m3_18054_6768# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.105547f
C387 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA6.A 0.301485f
C388 a_18882_35420# SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.133834f
C389 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_21402_35068# 0.129098f
C390 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_5648# 0.172147f
C391 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.30776f
C392 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.386137f
C393 VPWR a_5150_42408# 0.391292f
C394 VPWR uio_oe[0] 1.67769f
C395 SUNSAR_SAR8B_CV_0.XA4.XA2.A a_13842_30316# 0.129098f
C396 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.466806f
C397 SUNSAR_CAPT8B_CV_0.XE10.QN uo_out[4] 0.248612f
C398 VPWR SUNSAR_SAR8B_CV_0.D<1> 5.470241f
C399 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.246063f
C400 VPWR a_10170_35420# 0.39968f
C401 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.101993f
C402 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MP1.S 0.104609f
C403 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.93081f
C404 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.449584f
C405 VPWR a_18882_32076# 0.436368f
C406 VPWR a_5150_42760# 0.391454f
C407 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142956f
C408 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.179089f
C409 uo_out[4] TIE_L 0.31941f
C410 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> a_18882_33836# 0.103403f
C411 SUNSAR_SAR8B_CV_0.D<5> tt_um_TT06_SAR_done_0.DONE 0.295822f
C412 VPWR SUNSAR_SAR8B_CV_0.XA4.DONE 0.246222f
C413 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 27.1615f
C414 VPWR a_8822_43816# 0.391817f
C415 VPWR SUNSAR_SAR8B_CV_0.XA20.XA12.Y 1.13456f
C416 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.A 0.722887f
C417 a_7650_35420# SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.160931f
C418 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.D<1> 0.232115f
C419 a_3762_35420# SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.133834f
C420 SUNSAR_SAR8B_CV_0.XA6.XA10.A VPWR 0.780003f
C421 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 0.432466f
C422 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.898003f
C423 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 1.08082f
C424 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.284482f
C425 VPWR a_5130_32076# 0.436368f
C426 m3_18054_2928# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.105547f
C427 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.649845f
C428 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.CN 1.7759f
C429 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP2.S 0.155821f
C430 VPWR a_8802_35948# 0.417826f
C431 VPWR a_28727_39955# 0.355584f
C432 a_12690_32956# SUNSAR_SAR8B_CV_0.XA4.CP0 0.101124f
C433 VPWR a_18882_27852# 0.358599f
C434 VPWR a_23922_26796# 0.442318f
C435 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.437693f
C436 a_7650_36300# SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.13253f
C437 VPWR a_13862_40648# 0.491776f
C438 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XF11.QN 0.318734f
C439 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.386305f
C440 a_2630_41000# SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.114097f
C441 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B 27.1615f
C442 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.284482f
C443 VPWR TIE_L1 0.114647f
C444 VPWR a_8802_33836# 0.409601f
C445 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C446 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XA5.CP0 0.327909f
C447 VPWR a_18902_40648# 0.491776f
C448 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP2.S 0.150467f
C449 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CNO 0.504801f
C450 SUNSAR_SAR8B_CV_0.XA6.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.178114f
C451 uo_out[4] uio_oe[0] 0.550054f
C452 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.152052f
C453 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.271482f
C454 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN0 0.52234f
C455 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.CKN 0.200119f
C456 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.474658f
C457 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 2.72889f
C458 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.435464f
C459 SUNSAR_SAR8B_CV_0.XB2.XA4.GN ua[0] 0.765539f
C460 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N 0.204048f
C461 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.276413f
C462 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.41624f
C463 VPWR a_15230_42760# 0.391454f
C464 VPWR SUNSAR_SAR8B_CV_0.XA7.XA6.MP3.S 0.112098f
C465 VPWR SUNSAR_SAR8B_CV_0.XA3.XA11.MP1.S 0.101979f
C466 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.EN 1.04628f
C467 SUNSAR_CAPT8B_CV_0.XH13.QN SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.318734f
C468 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N 0.271482f
C469 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.375196f
C470 VPWR SUNSAR_SAR8B_CV_0.XB2.TIE_L 11.0126f
C471 VPWR SUNSAR_SAR8B_CV_0.D<4> 5.44389f
C472 VPWR SUNSAR_SAR8B_CV_0.XA3.XA4.A 2.31184f
C473 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.449584f
C474 a_10170_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C475 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.VMR 4.6743f
C476 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 4.25689f
C477 VPWR SUNSAR_SAR8B_CV_0.XA2.XA9.B 0.930839f
C478 VPWR a_20270_42760# 0.391454f
C479 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B SUNSAR_SAR8B_CV_0.XB1.CKN 0.26479f
C480 VPWR SUNSAR_SAR8B_CV_0.XA5.CEIN 2.30385f
C481 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.726497f
C482 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<1> 3.87301f
C483 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.EN 0.242472f
C484 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142977f
C485 VPWR a_18882_32956# 0.436368f
C486 uo_out[0] uio_out[0] 0.201579f
C487 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.201839f
C488 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N 0.271482f
C489 VPWR a_3762_37180# 0.473713f
C490 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.74594f
C491 tt_um_TT06_SAR_done_0.x3.MP1.G tt_um_TT06_SAR_done_0.DONE 0.186749f
C492 VPWR SUNSAR_SAR8B_CV_0.XB1.CKN 2.34497f
C493 VPWR a_15230_40296# 0.457171f
C494 SUNSAR_SAR8B_CV_0.XA7.XA10.A a_21402_35948# 0.134161f
C495 tt_um_TT06_SAR_done_0.DONE SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.403015f
C496 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 3.63372f
C497 SUNSAR_SAR8B_CV_0.XB1.XA4.GN ua[1] 0.762388f
C498 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.QN 0.318734f
C499 VPWR a_13842_36300# 0.399161f
C500 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA2.EN 0.129613f
C501 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.12241f
C502 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.301485f
C503 SUNSAR_CAPT8B_CV_0.XI14.QN uo_out[0] 0.24816f
C504 VPWR a_20270_40296# 0.456842f
C505 VPWR a_3782_42760# 0.391454f
C506 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.101001f
C507 SUNSAR_SAR8B_CV_0.D<7> a_2610_31196# 0.11099f
C508 VPWR a_15210_30316# 0.404384f
C509 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.437693f
C510 VPWR SUNSAR_SAR8B_CV_0.XA6.XA6.MP3.S 0.112858f
C511 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S 0.101001f
C512 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B 3.55549f
C513 VPWR a_5130_31196# 0.44007f
C514 VPWR a_18902_41880# 0.395781f
C515 a_22790_42408# SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.10248f
C516 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.300065f
C517 TIE_L clk 0.146712f
C518 VPWR SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H 0.452478f
C519 VPWR SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G 0.519052f
C520 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.297144f
C521 uio_out[0] uo_out[5] 0.109219f
C522 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.MP1.S 0.119314f
C523 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142977f
C524 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_5150_41000# 0.156079f
C525 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.63636f
C526 VPWR a_5130_33836# 0.409601f
C527 VPWR SUNSAR_SAR8B_CV_0.XA5.DONE 0.245452f
C528 VPWR SUNSAR_SAR8B_CV_0.XA2.CEIN 1.06023f
C529 VPWR SUNSAR_SAR8B_CV_0.XA20.CNO 6.94539f
C530 VPWR a_13842_28204# 0.36179f
C531 a_7650_32956# SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.101124f
C532 a_13950_3686# SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.16579f
C533 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111217f
C534 a_7670_42408# SUNSAR_CAPT8B_CV_0.XD09.XA5.A 0.111909f
C535 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.108405f
C536 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.201839f
C537 SUNSAR_SAR8B_CV_0.XB2.XA4.GN SUNSAR_SAR8B_CV_0.SARN 0.36754f
C538 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.22339f
C539 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.80606f
C540 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA4.MP1.S 0.104609f
C541 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.220689f
C542 VPWR a_3762_37532# 0.458479f
C543 m3_9126_3888# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.105547f
C544 VPWR SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 1.50269f
C545 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.380687f
C546 VPWR a_20250_27148# 0.470364f
C547 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR a_23922_30844# 0.100515f
C548 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C549 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA5.A 0.898003f
C550 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 13.6519f
C551 VPWR a_3782_41880# 0.395781f
C552 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.D<4> 0.233744f
C553 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.CN0 0.671839f
C554 clk uio_oe[0] 0.260056f
C555 SUNSAR_SAR8B_CV_0.XA4.DONE SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.143554f
C556 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18344f
C557 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 1.7759f
C558 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.189112f
C559 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C560 VPWR a_10170_31196# 0.44007f
C561 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 1.77591f
C562 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA6.A 0.301485f
C563 VPWR a_15230_43288# 0.394205f
C564 SUNSAR_SAR8B_CV_0.XA2.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.377598f
C565 VPWR a_3782_41352# 0.394053f
C566 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.393076f
C567 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.252966f
C568 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.SARN 0.591428f
C569 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MP1.S 0.104609f
C570 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.D<4> 0.625175f
C571 VPWR SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H 0.452478f
C572 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.CN1 0.466806f
C573 VPWR SUNSAR_SAR8B_CV_0.XA4.XA4.A 2.31184f
C574 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 4.25322f
C575 SUNSAR_SAR8B_CV_0.D<3> tt_um_TT06_SAR_done_0.DONE 0.295397f
C576 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.449584f
C577 SUNSAR_SAR8B_CV_0.XA4.XA11.A SUNSAR_SAR8B_CV_0.XA4.CEIN 0.303978f
C578 VPWR SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.720133f
C579 VPWR a_20250_35948# 0.414756f
C580 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 1.20727f
C581 VPWR SUNSAR_CAPT8B_CV_0.XB07.QN 0.901622f
C582 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA10.Y 1.59176f
C583 VPWR a_18902_41352# 0.394053f
C584 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 0.419738f
C585 VPWR a_13842_35948# 0.417826f
C586 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<3> 0.105016f
C587 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_SAR8B_CV_0.D<1> 0.393049f
C588 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA3.EN 0.3401f
C589 SUNSAR_SAR8B_CV_0.XA7.XA9.A tt_um_TT06_SAR_done_0.DONE 0.182408f
C590 VPWR a_18882_29612# 0.397362f
C591 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.142956f
C592 SUNSAR_CAPT8B_CV_0.XD09.XA6.A a_8822_42760# 0.113305f
C593 VPWR a_20250_30316# 0.403745f
C594 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA20.CPO 0.328435f
C595 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111217f
C596 SUNSAR_SAR8B_CV_0.XB2.TIE_L ua[1] 0.837206f
C597 VPWR SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.720114f
C598 VPWR a_23942_42760# 0.388156f
C599 VPWR a_3782_43816# 0.391817f
C600 a_11322_36828# SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.104051f
C601 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.152045f
C602 m3_18054_3888# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.105547f
C603 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 0.164325f
C604 VPWR a_10170_35068# 0.394528f
C605 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.267238f
C606 a_11322_32956# SUNSAR_SAR8B_CV_0.XA3.CP0 0.102695f
C607 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 3.55251f
C608 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2165f
C609 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G SUNSAR_SAR8B_CV_0.XA20.CPO 0.143023f
C610 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.EN 0.13041f
C611 SUNSAR_SAR8B_CV_0.XA2.DONE SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.143554f
C612 a_16362_35948# SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.134161f
C613 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 0.363295f
C614 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.MP1.S 0.106927f
C615 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_4688# 0.172147f
C616 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.166272f
C617 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN 0.3401f
C618 VPWR uo_out[4] 1.03021f
C619 m3_18054_5808# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.105547f
C620 VPWR SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.725614f
C621 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.201839f
C622 SUNSAR_SAR8B_CV_0.XB1.CKN ua[1] 0.175642f
C623 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.EN 0.893904f
C624 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B m3_2358_6608# 0.172147f
C625 VPWR a_8802_27852# 0.358599f
C626 SUNSAR_SAR8B_CV_0.XA0.XA9.A SUNSAR_SAR8B_CV_0.XA1.EN 0.144331f
C627 a_7650_36828# SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.10248f
C628 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.CEIN 0.352238f
C629 VPWR a_23922_34540# 0.502044f
C630 a_5130_35420# VPWR 0.39968f
C631 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.290432f
C632 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B 0.419738f
C633 SUNSAR_CAPT8B_CV_0.XC08.XA7.C a_6302_41000# 0.115667f
C634 VPWR a_8802_34716# 0.399819f
C635 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.845515f
C636 VPWR a_23922_30844# 0.425847f
C637 VPWR a_10190_42760# 0.391454f
C638 VPWR a_15210_27500# 0.382397f
C639 VPWR a_5150_44168# 0.340085f
C640 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.276252f
C641 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA20.CNO 0.180455f
C642 VPWR a_5130_28556# 0.406628f
C643 VPWR SUNSAR_SAR8B_CV_0.D<2> 5.45951f
C644 VPWR SUNSAR_SAR8B_CV_0.XA6.DONE 0.246222f
C645 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.432466f
C646 VPWR SUNSAR_CAPT8B_CV_0.XA2.MP0.G 0.667429f
C647 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA6.A 1.63909f
C648 VPWR a_20270_42408# 0.391292f
C649 uo_out[3] TIE_L 0.185333f
C650 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.206912f
C651 VPWR a_16542_4038# 0.379979f
C652 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 0.449584f
C653 VPWR a_23922_36652# 0.449853f
C654 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B 3.55251f
C655 a_12690_35420# SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.160931f
C656 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B 13.6519f
C657 SUNSAR_CAPT8B_CV_0.XG12.QN uo_out[2] 0.249322f
C658 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B 0.419738f
C659 SUNSAR_SAR8B_CV_0.XA5.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.791351f
C660 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA6.B 0.504864f
C661 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 6.86675f
C662 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N 0.271482f
C663 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 5.19722f
C664 VPWR SUNSAR_SAR8B_CV_0.D<7> 3.79388f
C665 VPWR SUNSAR_SAR8B_CV_0.XA3.CN1 2.62342f
C666 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.241356f
C667 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03123f
C668 SUNSAR_CAPT8B_CV_0.XA5.B a_22790_41000# 0.11811f
C669 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA4.CEIN 0.13078f
C670 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.CN1 0.702226f
C671 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.EN 0.340491f
C672 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.146492f
C673 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.A 1.22023f
C674 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B ua[1] 0.241597f
C675 SUNSAR_SAR8B_CV_0.XA7.XA10.A SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.205884f
C676 VPWR a_13862_41000# 0.388305f
C677 VPWR a_13862_43816# 0.391817f
C678 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA2.EN 0.154232f
C679 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C680 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03123f
C681 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CN1 0.625035f
C682 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S 0.104122f
C683 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.126806f
C684 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.63636f
C685 VPWR ua[1] 0.349347f
C686 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA3.MP1.S 0.106927f
C687 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 1.38576f
C688 uo_out[3] uio_oe[0] 0.212351f
C689 VPWR a_13842_36828# 0.395703f
C690 a_12690_36828# SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.10248f
C691 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.238862f
C692 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.178114f
C693 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_SAR8B_CV_0.D<3> 0.393049f
C694 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.170578f
C695 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.649845f
C696 SUNSAR_SAR8B_CV_0.XA0.XA9.A a_2610_35068# 0.127528f
C697 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA7.XA2.A 0.118152f
C698 VPWR SUNSAR_SAR8B_CV_0.XA3.EN 5.52623f
C699 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.A 1.22023f
C700 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 13.6519f
C701 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.206292f
C702 SUNSAR_CAPT8B_CV_0.XE10.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C703 VPWR a_23922_29964# 0.429137f
C704 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.178114f
C705 VPWR a_15210_35068# 0.394528f
C706 VPWR SUNSAR_SAR8B_CV_0.XA2.XA4.A 2.31184f
C707 VPWR SUNSAR_SAR8B_CV_0.XA5.EN 5.52623f
C708 VPWR a_8802_32956# 0.436368f
C709 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XD09.QN 0.318734f
C710 VPWR a_16542_5622# 0.472384f
C711 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA2.EN 0.144331f
C712 VPWR a_13862_41880# 0.395781f
C713 VPWR SUNSAR_SAR8B_CV_0.XA1.XA6.MP3.S 0.112858f
C714 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.215251f
C715 SUNSAR_CAPT8B_CV_0.XE10.XA6.A a_10190_42760# 0.111734f
C716 VPWR clk 0.644902f
C717 VPWR a_10170_32076# 0.436368f
C718 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN uo_out[3] 0.309657f
C719 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.34399f
C720 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP2.S 0.155821f
C721 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.437693f
C722 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.118161f
C723 a_10170_35420# SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.133834f
C724 SUNSAR_CAPT8B_CV_0.XH13.QN uo_out[1] 0.248827f
C725 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA7.C 2.9722f
C726 a_13950_5446# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.102604f
C727 a_12582_5094# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.160184f
C728 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.149144f
C729 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 6.19724f
C730 VPWR a_10170_30316# 0.404384f
C731 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN uo_out[2] 0.305131f
C732 VPWR a_18882_28908# 0.395394f
C733 SUNSAR_SAR8B_CV_0.XA6.XA10.A SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.205884f
C734 SUNSAR_SAR8B_CV_0.XA0.XA11.A SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.300886f
C735 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA2.EN 0.118226f
C736 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.118161f
C737 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA7.C 2.97208f
C738 SUNSAR_SAR8B_CV_0.XA2.XA10.A SUNSAR_SAR8B_CV_0.XA2.XA11.A 0.201839f
C739 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 0.635098f
C740 VPWR a_18882_28204# 0.36179f
C741 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.898003f
C742 VPWR a_15230_41352# 0.394053f
C743 SUNSAR_SAR8B_CV_0.XA6.DONE SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.143554f
C744 SUNSAR_SAR8B_CV_0.D<1> tt_um_TT06_SAR_done_0.DONE 0.295407f
C745 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.EN 0.166192f
C746 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.179089f
C747 VPWR a_3762_36300# 0.399161f
C748 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 1.06875f
C749 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 3.09787f
C750 VPWR SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.780003f
C751 VPWR SUNSAR_CAPT8B_CV_0.XA5.B 1.20915f
C752 VPWR a_10170_26796# 0.441753f
C753 SUNSAR_SAR8B_CV_0.XA7.CN1 SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.466806f
C754 m3_9126_2928# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.105547f
C755 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARN 0.175967f
C756 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> a_5130_33836# 0.101833f
C757 VPWR a_8822_41880# 0.395781f
C758 VPWR a_10190_42408# 0.391292f
C759 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.109021f
C760 SUNSAR_SAR8B_CV_0.XB2.TIE_L ua[0] 1.50732f
C761 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 0.107427f
C762 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.475004f
C763 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN uo_out[1] 0.305131f
C764 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.101993f
C765 SUNSAR_SAR8B_CV_0.XA6.XA12.A a_17730_36828# 0.10248f
C766 SUNSAR_CAPT8B_CV_0.XD09.QN a_7670_43816# 0.127669f
C767 VPWR a_13842_28908# 0.395394f
C768 VPWR a_8822_41352# 0.394053f
C769 VPWR a_23942_41352# 0.376408f
C770 SUNSAR_SAR8B_CV_0.XA7.XA9.A a_20250_35420# 0.133834f
C771 VPWR a_13842_26796# 0.442908f
C772 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.XA5.XA2.A 0.702226f
C773 TIE_L uo_out[1] 0.50141f
C774 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 4.24508f
C775 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.S 0.137646f
C776 VPWR SUNSAR_SAR8B_CV_0.XA4.CEIN 1.06023f
C777 VPWR a_5130_37180# 0.474051f
C778 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_SAR8B_CV_0.D<2> 0.393063f
C779 VPWR SUNSAR_SAR8B_CV_0.XA5.XA6.MP3.S 0.112858f
C780 VPWR SUNSAR_SAR8B_CV_0.XA1.DONE 0.245452f
C781 SUNSAR_SAR8B_CV_0.XA6.XA2.A SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.133602f
C782 a_12710_41000# SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.114097f
C783 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.724217f
C784 a_12710_43816# SUNSAR_CAPT8B_CV_0.XF11.QN 0.127669f
C785 VPWR a_10190_40296# 0.457269f
C786 SUNSAR_CAPT8B_CV_0.XF11.XA6.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.649845f
C787 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP2.S 0.150467f
C788 a_8802_35420# SUNSAR_SAR8B_CV_0.XA2.XA9.A 0.133834f
C789 a_7650_31196# SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.110962f
C790 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.144778f
C791 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 3.0515f
C792 a_5130_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C793 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.722427f
C794 VPWR SUNSAR_SAR8B_CV_0.XA0.XA11.A 0.728421f
C795 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.B 0.93081f
C796 SUNSAR_SAR8B_CV_0.D<4> tt_um_TT06_SAR_done_0.DONE 0.295493f
C797 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.EN 0.793076f
C798 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA4.MP1.S 0.106927f
C799 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XA3.CP0 0.791351f
C800 SUNSAR_SAR8B_CV_0.XA4.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.377598f
C801 VPWR SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G 0.808658f
C802 m3_18054_4848# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 0.105547f
C803 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.16676f
C804 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XA3.EN 0.118161f
C805 VPWR SUNSAR_SAR8B_CV_0.XA0.XA6.MP3.S 0.112858f
C806 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.116058f
C807 VPWR a_5130_37532# 0.459635f
C808 TIE_L uo_out[6] 0.204625f
C809 VPWR a_5150_43288# 0.394205f
C810 uo_out[1] uio_oe[0] 0.432144f
C811 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.144331f
C812 VPWR a_8802_28204# 0.36179f
C813 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.204048f
C814 VPWR a_13842_27852# 0.358599f
C815 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 0.128204f
C816 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.EN 0.952619f
C817 VPWR a_28727_40307# 0.410063f
C818 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.284482f
C819 VPWR uo_out[3] 1.25759f
C820 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.250503f
C821 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 4.24834f
C822 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA4.MP1.S 0.104609f
C823 VPWR a_13842_34716# 0.399819f
C824 SUNSAR_CAPT8B_CV_0.XE10.XA5.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.432466f
C825 VPWR a_5150_40648# 0.493192f
C826 VPWR SUNSAR_SAR8B_CV_0.XA4.XA6.MP3.S 0.112858f
C827 SUNSAR_CAPT8B_CV_0.XD09.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.233892f
C828 a_12690_35068# SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.127528f
C829 SUNSAR_SAR8B_CV_0.XA1.XA11.A SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.201839f
C830 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA4.MP1.S 0.106927f
C831 VPWR a_10170_37180# 0.474068f
C832 VPWR a_3762_27852# 0.358599f
C833 SUNSAR_CAPT8B_CV_0.XI14.XA6.A a_20270_42760# 0.111734f
C834 VPWR a_10170_28556# 0.406628f
C835 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.201839f
C836 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN 0.154232f
C837 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP2.S 0.152518f
C838 VPWR a_13862_42408# 0.391292f
C839 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B 0.635098f
C840 a_8802_33836# SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.103403f
C841 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.538639f
C842 SUNSAR_CAPT8B_CV_0.XI14.XA5.A SUNSAR_CAPT8B_CV_0.XI14.XA7.C 0.12241f
C843 VPWR SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.930839f
C844 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA2.CEIN 0.432008f
C845 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.41635f
C846 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B 0.441867f
C847 VPWR a_28727_40659# 0.39147f
C848 VPWR ua[0] 0.629451f
C849 VPWR SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 1.05322f
C850 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.182744f
C851 SUNSAR_SAR8B_CV_0.XA0.XA12.A SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.222689f
C852 VPWR a_13842_28556# 0.406628f
C853 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N 0.271482f
C854 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.SARN 0.205975f
C855 VPWR SUNSAR_SAR8B_CV_0.XB2.CKN 2.34497f
C856 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA4.MP1.S 0.106927f
C857 a_15210_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C858 SUNSAR_SAR8B_CV_0.XA6.CP0 a_17730_32956# 0.101124f
C859 VPWR a_16542_4566# 0.413433f
C860 uo_out[2] TIE_L 0.156661f
C861 SUNSAR_SAR8B_CV_0.XA2.XA12.A SUNSAR_SAR8B_CV_0.XA2.CEIN 0.220689f
C862 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.EN 0.339883f
C863 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.A 1.2202f
C864 VPWR a_20250_27500# 0.382397f
C865 uo_out[7] TIE_L 0.471918f
C866 SUNSAR_SAR8B_CV_0.XA3.EN a_7650_28556# 0.132757f
C867 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA9.Y 0.530644f
C868 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN uo_out[5] 0.30523f
C869 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.199693f
C870 a_6282_35948# SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.134161f
C871 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1625f
C872 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.437693f
C873 SUNSAR_CAPT8B_CV_0.XD09.XA7.C a_8822_41000# 0.15757f
C874 SUNSAR_CAPT8B_CV_0.XE10.XA7.C SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.63636f
C875 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB2.CKN 0.200119f
C876 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA4.MP1.S 0.106927f
C877 VPWR SUNSAR_SAR8B_CV_0.XA1.CEIN 2.30575f
C878 VPWR a_3762_35068# 0.394528f
C879 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XA20.CNO 0.189429f
C880 VPWR a_15210_35420# 0.39968f
C881 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.6934f
C882 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.63636f
C883 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA6.CEIN 0.13078f
C884 a_13950_2982# SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.158066f
C885 VPWR a_3782_41000# 0.388305f
C886 VPWR a_20250_37532# 0.454489f
C887 VPWR SUNSAR_SAR8B_CV_0.XA1.XA9.A 1.2202f
C888 uo_out[4] uo_out[3] 0.854997f
C889 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 3.55251f
C890 VPWR SUNSAR_SAR8B_CV_0.XA2.XA12.A 0.723762f
C891 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.MP1.S 0.106927f
C892 SUNSAR_SAR8B_CV_0.XA0.XA9.B SUNSAR_SAR8B_CV_0.XA0.XA10.A 0.205884f
C893 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N 0.154232f
C894 a_15390_3334# SUNSAR_SAR8B_CV_0.XB2.CKN 0.113134f
C895 a_13950_3334# SUNSAR_SAR8B_CV_0.XB2.XA4.GN 0.163985f
C896 SUNSAR_CAPT8B_CV_0.XD09.QN uo_out[5] 0.248535f
C897 VPWR a_5130_30316# 0.404384f
C898 VPWR tt_um_TT06_SAR_done_0.DONE 8.70939f
C899 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C900 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA7.C 2.97221f
C901 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.466806f
C902 a_22790_42760# SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.13379f
C903 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.S 0.138148f
C904 uo_out[2] uio_oe[0] 0.267754f
C905 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN VPWR 1.7759f
C906 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.62393f
C907 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C908 VPWR a_13862_44168# 0.3405f
C909 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.D<4> 0.503825f
C910 VPWR SUNSAR_SAR8B_CV_0.XA2.DONE 0.246222f
C911 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 3.55251f
C912 uo_out[7] uio_oe[0] 0.43252f
C913 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA4.A 0.118226f
C914 VPWR a_9990_4918# 0.468783f
C915 a_17730_35068# SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.127528f
C916 SUNSAR_CAPT8B_CV_0.XA5.B clk 0.210661f
C917 SUNSAR_SAR8B_CV_0.XA7.ENO a_21402_28556# 0.134248f
C918 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.394834f
C919 SUNSAR_SAR8B_CV_0.D<2> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 2.4271f
C920 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.ENO 0.144331f
C921 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.293159f
C922 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.C 2.97213f
C923 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA6.A 1.63909f
C924 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA7.C 0.12241f
C925 VPWR a_3762_32956# 0.436368f
C926 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 1.88588f
C927 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.63636f
C928 a_16362_35068# SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.129098f
C929 VPWR SUNSAR_SAR8B_CV_0.XA1.XA4.A 2.31184f
C930 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.SARN 3.55251f
C931 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.431984f
C932 VPWR SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 1.50177f
C933 SUNSAR_CAPT8B_CV_0.XI14.XA6.A SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.744161f
C934 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.D<4> 2.42393f
C935 VPWR SUNSAR_SAR8B_CV_0.XA6.EN 4.84607f
C936 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.D<4> 0.17528f
C937 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.718455f
C938 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<6> 1.62595f
C939 a_16382_41000# SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.115667f
C940 VPWR SUNSAR_SAR8B_CV_0.SARN 0.133035f
C941 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.123668f
C942 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 0.437693f
C943 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 1.06875f
C944 VPWR SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.728492f
C945 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.EN 0.11263f
C946 tt_um_TT06_SAR_done_0.x3.MP1.G uio_out[0] 0.165429f
C947 VPWR a_20270_44168# 0.340085f
C948 a_16542_4038# SUNSAR_SAR8B_CV_0.XB2.CKN 0.135393f
C949 VPWR SUNSAR_SAR8B_CV_0.XA20.XA9.Y 3.91346f
C950 SUNSAR_CAPT8B_CV_0.XB07.XA7.C SUNSAR_CAPT8B_CV_0.XB07.QN 0.318734f
C951 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.310451f
C952 VPWR a_20250_28556# 0.406628f
C953 TIE_L1 uo_out[7] 0.206895f
C954 a_5130_35420# SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.133834f
C955 VPWR SUNSAR_SAR8B_CV_0.D<0> 5.69433f
C956 VPWR a_5130_26796# 0.441753f
C957 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.SARN 0.259325f
C958 SUNSAR_CAPT8B_CV_0.XD09.XA6.A SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.744161f
C959 VPWR a_10170_36300# 0.398846f
C960 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 4.27988f
C961 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S 0.104122f
C962 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.441867f
C963 SUNSAR_SAR8B_CV_0.XA6.XA9.A SUNSAR_SAR8B_CV_0.XA6.XA9.B 0.527529f
C964 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.241356f
C965 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.18612f
C966 VPWR a_18902_43816# 0.391817f
C967 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.898003f
C968 VPWR SUNSAR_CAPT8B_CV_0.XC08.QN 0.901622f
C969 VPWR a_5130_34716# 0.399819f
C970 SUNSAR_CAPT8B_CV_0.XF11.XA6.A a_13862_42760# 0.113305f
C971 VPWR a_5130_27500# 0.382397f
C972 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA1.EN 0.118161f
C973 SUNSAR_SAR8B_CV_0.XA3.XA9.B SUNSAR_SAR8B_CV_0.XA3.XA10.A 0.205884f
C974 VPWR ui_in[0] 2.01351f
C975 SUNSAR_SAR8B_CV_0.D<2> tt_um_TT06_SAR_done_0.DONE 0.295646f
C976 ua[1] ua[0] 3.85017f
C977 VPWR SUNSAR_SAR8B_CV_0.XA7.XA11.MP1.S 0.101562f
C978 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.MP1.S 0.106927f
C979 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MP1.S 0.108436f
C980 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.118161f
C981 SUNSAR_CAPT8B_CV_0.XH13.XA5.A SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.301485f
C982 VPWR a_3762_28908# 0.395394f
C983 VPWR a_18902_43288# 0.394205f
C984 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 0.167f
C985 VPWR uo_out[1] 1.02322f
C986 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.D<2> 0.137975f
C987 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.S 0.137646f
C988 SUNSAR_SAR8B_CV_0.XA4.XA11.A a_12690_36300# 0.13253f
C989 VPWR SUNSAR_SAR8B_CV_0.XA4.CN1 2.62342f
C990 VPWR SUNSAR_SAR8B_CV_0.XA4.EN 4.84607f
C991 VPWR a_13842_31196# 0.44007f
C992 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.228326f
C993 a_10190_41000# SUNSAR_CAPT8B_CV_0.XE10.XA7.C 0.156079f
C994 a_22770_29964# SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.134249f
C995 m3_24750_4688# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.172147f
C996 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.126806f
C997 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA3.MP1.S 0.106927f
C998 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.CNO 0.159359f
C999 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA20.CNO 2.96993f
C1000 SUNSAR_SAR8B_CV_0.D<7> tt_um_TT06_SAR_done_0.DONE 0.292137f
C1001 SUNSAR_CAPT8B_CV_0.XF11.XA5.A SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.12241f
C1002 SUNSAR_SAR8B_CV_0.D<4> SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.241356f
C1003 VPWR a_18882_26796# 0.442908f
C1004 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP2.S 0.155821f
C1005 VPWR SUNSAR_SAR8B_CV_0.XA7.CN1 2.62711f
C1006 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA7.C 2.97211f
C1007 m3_24750_6608# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.172147f
C1008 SUNSAR_CAPT8B_CV_0.XI14.XA7.C a_20270_41000# 0.156079f
C1009 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.178111f
C1010 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.744161f
C1011 VPWR SUNSAR_SAR8B_CV_0.XA7.CEIN 2.28789f
C1012 VPWR a_15210_32076# 0.436368f
C1013 VPWR SUNSAR_SAR8B_CV_0.XA3.XA6.MP3.S 0.112858f
C1014 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.XA4.CN1 0.466806f
C1015 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.D<2> 0.503825f
C1016 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.129613f
C1017 VPWR a_18882_36300# 0.399161f
C1018 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.107674f
C1019 TIE_L uo_out[0] 0.280844f
C1020 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.18141f
C1021 a_8802_30316# SUNSAR_SAR8B_CV_0.XA2.XA2.A 0.129098f
C1022 VPWR SUNSAR_SAR8B_CV_0.XA3.DONE 0.245452f
C1023 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 4.2492f
C1024 VPWR SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.765792f
C1025 SUNSAR_SAR8B_CV_0.XA4.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.791379f
C1026 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 2.72582f
C1027 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.393125f
C1028 VPWR uo_out[6] 1.34623f
C1029 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B 0.449584f
C1030 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.618979f
C1031 VPWR SUNSAR_SAR8B_CV_0.EN 41.914997f
C1032 a_6282_36828# SUNSAR_SAR8B_CV_0.XA1.XA12.A 0.104051f
C1033 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.693521f
C1034 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B 0.441867f
C1035 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.SARP 0.102632f
C1036 VPWR a_10190_41352# 0.394053f
C1037 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 0.316693f
C1038 VPWR a_5130_35948# 0.417826f
C1039 SUNSAR_SAR8B_CV_0.XA20.XA3.CO SUNSAR_SAR8B_CV_0.XA20.CPO 0.464697f
C1040 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.162703f
C1041 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.SARN 0.161316f
C1042 VPWR a_10190_40648# 0.493224f
C1043 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.10132f
C1044 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.398331f
C1045 VPWR a_13842_27148# 0.471462f
C1046 SUNSAR_CAPT8B_CV_0.XA6.B SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.134182f
C1047 VPWR a_10170_37532# 0.459696f
C1048 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA3.MP1.S 0.106927f
C1049 VPWR a_20250_37180# 0.469114f
C1050 m3_24750_2768# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.172147f
C1051 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.535136f
C1052 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.193518f
C1053 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B 27.1615f
C1054 SUNSAR_SAR8B_CV_0.XA4.XA4.A SUNSAR_SAR8B_CV_0.EN 0.112859f
C1055 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.C 2.97208f
C1056 VPWR a_8822_43288# 0.394205f
C1057 VPWR a_3762_29612# 0.397362f
C1058 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA4.MP1.S 0.106927f
C1059 SUNSAR_SAR8B_CV_0.XA20.XA11.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.106002f
C1060 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.294852f
C1061 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 1.05322f
C1062 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.105906f
C1063 VPWR a_15210_37532# 0.459576f
C1064 TIE_L uo_out[5] 1.3092f
C1065 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> a_6282_32956# 0.102695f
C1066 uo_out[0] uio_oe[0] 0.670799f
C1067 VPWR a_18882_34716# 0.399819f
C1068 a_9990_4038# SUNSAR_SAR8B_CV_0.XB1.CKN 0.135393f
C1069 VPWR SUNSAR_SAR8B_CV_0.XA7.CP0 2.66621f
C1070 VPWR a_15210_37180# 0.474036f
C1071 SUNSAR_SAR8B_CV_0.SARN ua[1] 0.806872f
C1072 VPWR a_18882_33836# 0.409601f
C1073 VPWR uo_out[2] 1.02322f
C1074 a_18882_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C1075 VPWR a_18902_41000# 0.388305f
C1076 SUNSAR_CAPT8B_CV_0.XG12.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1077 VPWR SUNSAR_SAR8B_CV_0.XA5.CN1 2.62342f
C1078 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C1079 VPWR uo_out[7] 1.27659f
C1080 VPWR SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.324111f
C1081 VPWR a_8802_28908# 0.395394f
C1082 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.308722f
C1083 VPWR a_15210_33836# 0.409601f
C1084 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.XA12.A 0.377598f
C1085 VPWR a_18882_36828# 0.395703f
C1086 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.CPO 0.372599f
C1087 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.EN 1.2771f
C1088 VPWR SUNSAR_SAR8B_CV_0.XA0.DONE 0.247527f
C1089 VPWR SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.723713f
C1090 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.204048f
C1091 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N 0.279205f
C1092 SUNSAR_SAR8B_CV_0.XA2.XA9.B SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.205884f
C1093 uo_out[4] uo_out[6] 0.843602f
C1094 VPWR a_5130_28204# 0.361706f
C1095 SUNSAR_CAPT8B_CV_0.XH13.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1096 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CNO 0.276413f
C1097 VPWR a_5130_27148# 0.470364f
C1098 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.363295f
C1099 VPWR SUNSAR_SAR8B_CV_0.XA4.XA9.B 0.930839f
C1100 VPWR SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 1.7759f
C1101 SUNSAR_SAR8B_CV_0.XA3.XA4.A SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.133602f
C1102 VPWR a_15210_32956# 0.436368f
C1103 a_18882_30316# SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.129098f
C1104 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.321724f
C1105 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B 0.449584f
C1106 SUNSAR_CAPT8B_CV_0.XC08.XA5.A SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.12241f
C1107 SUNSAR_SAR8B_CV_0.XA1.EN a_2610_28556# 0.132757f
C1108 uio_oe[0] uo_out[5] 1.55329f
C1109 VPWR a_8822_44168# 0.3405f
C1110 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA4.MP1.S 0.106927f
C1111 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.B 0.94014f
C1112 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B 0.437693f
C1113 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA5.A 0.432466f
C1114 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.S 0.138148f
C1115 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.QN 0.263255f
C1116 VPWR a_8802_36828# 0.396052f
C1117 VPWR a_20250_35420# 0.39661f
C1118 VPWR a_13842_29612# 0.397362f
C1119 SUNSAR_CAPT8B_CV_0.XI14.XA5.A a_21422_42408# 0.113479f
C1120 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.S 0.138148f
C1121 a_17730_35420# SUNSAR_SAR8B_CV_0.XA6.XA9.A 0.160931f
C1122 VPWR SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.779986f
C1123 SUNSAR_SAR8B_CV_0.XA6.CP0 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 0.791379f
C1124 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 1.26537f
C1125 VPWR a_3782_42408# 0.391292f
C1126 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW SUNSAR_SAR8B_CV_0.XB2.TIE_L 6.83332f
C1127 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.122781f
C1128 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N 0.271482f
C1129 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2173f
C1130 a_12690_31196# SUNSAR_SAR8B_CV_0.XA4.CN1 0.107567f
C1131 a_16362_35420# SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.160931f
C1132 VPWR a_8802_35420# 0.39968f
C1133 m3_2358_2768# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.172147f
C1134 VPWR a_9990_4038# 0.379979f
C1135 a_13862_41000# SUNSAR_CAPT8B_CV_0.XF11.XA7.C 0.15757f
C1136 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111173f
C1137 SUNSAR_CAPT8B_CV_0.XC08.QN a_6302_43816# 0.129239f
C1138 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.231927f
C1139 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 1.06875f
C1140 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> SUNSAR_SAR8B_CV_0.D<4> 2.09966f
C1141 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B 6.86675f
C1142 uo_out[7] uo_out[4] 0.121648f
C1143 a_11142_3334# SUNSAR_SAR8B_CV_0.XB1.CKN 0.114704f
C1144 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.EN 1.2771f
C1145 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.EN 0.37807f
C1146 SUNSAR_SAR8B_CV_0.XB1.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.169642f
C1147 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.EN 0.343905f
C1148 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.204048f
C1149 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA7.MP1.S 0.106927f
C1150 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 0.635098f
C1151 clk ui_in[0] 0.169609f
C1152 SUNSAR_CAPT8B_CV_0.XG12.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.12241f
C1153 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B 0.419738f
C1154 a_2610_35420# SUNSAR_SAR8B_CV_0.XA0.XA9.A 0.160931f
C1155 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA7.MP1.S 0.106927f
C1156 VPWR SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S 0.429492f
C1157 TIE_L1 uo_out[5] 0.275794f
C1158 SUNSAR_SAR8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.133602f
C1159 VPWR tt_um_TT06_SAR_done_0.x4.MP0.G 0.511762f
C1160 SUNSAR_SAR8B_CV_0.XA1.XA9.A SUNSAR_SAR8B_CV_0.XA1.DONE 0.145738f
C1161 VPWR a_3762_32076# 0.436368f
C1162 uo_out[4] SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.305131f
C1163 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 0.139471f
C1164 SUNSAR_SAR8B_CV_0.XA5.CN1 SUNSAR_SAR8B_CV_0.D<2> 0.625175f
C1165 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 2.59087f
C1166 VPWR SUNSAR_SAR8B_CV_0.XA6.XA4.A 2.31184f
C1167 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XA20.XA10.Y 0.506551f
C1168 a_2630_42408# SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.111909f
C1169 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.133602f
C1170 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA9.A 0.527529f
C1171 VPWR SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.93081f
C1172 VPWR SUNSAR_SAR8B_CV_0.XA2.XA10.A 0.780003f
C1173 TIE_L uio_out[0] 0.44106f
C1174 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B 0.437693f
C1175 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.EN 1.02916f
C1176 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.CK_CMP 0.127551f
C1177 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_4848# 0.105547f
C1178 VPWR a_5150_40296# 0.457199f
C1179 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 54.2165f
C1180 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.S 0.137646f
C1181 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G 1.06875f
C1182 VPWR SUNSAR_SAR8B_CV_0.XA1.XA2.A 2.45309f
C1183 SUNSAR_SAR8B_CV_0.XB2.CKN ua[0] 0.175642f
C1184 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.EN 0.112859f
C1185 SUNSAR_SAR8B_CV_0.XA7.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.183415f
C1186 VPWR SUNSAR_SAR8B_CV_0.XA3.XA2.A 2.45309f
C1187 SUNSAR_SAR8B_CV_0.XA5.EN SUNSAR_SAR8B_CV_0.EN 1.02916f
C1188 SUNSAR_CAPT8B_CV_0.XH13.XA7.C uo_out[1] 0.245678f
C1189 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MP1.S 0.104609f
C1190 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B 6.86675f
C1191 SUNSAR_CAPT8B_CV_0.XE10.XA6.A SUNSAR_CAPT8B_CV_0.XE10.XA7.CN 0.744161f
C1192 SUNSAR_CAPT8B_CV_0.XF11.XA7.C SUNSAR_CAPT8B_CV_0.XG12.XA7.C 0.233892f
C1193 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_6768# 0.105547f
C1194 VPWR a_13862_42760# 0.391454f
C1195 VPWR SUNSAR_SAR8B_CV_0.XA0.XA9.A 1.22398f
C1196 SUNSAR_CAPT8B_CV_0.XB07.XA6.A SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.301485f
C1197 VPWR SUNSAR_SAR8B_CV_0.XA7.XA12.A 0.714341f
C1198 SUNSAR_SAR8B_CV_0.XA7.XA10.A VPWR 0.774301f
C1199 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.S 0.137646f
C1200 SUNSAR_CAPT8B_CV_0.XA5.B ui_in[0] 0.17256f
C1201 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN a_15230_41880# 0.100592f
C1202 SUNSAR_SAR8B_CV_0.XA3.XA11.A SUNSAR_SAR8B_CV_0.XA3.CEIN 0.352238f
C1203 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.126806f
C1204 VPWR a_10170_35948# 0.417826f
C1205 VPWR a_10170_27148# 0.470364f
C1206 VPWR a_10170_27500# 0.382397f
C1207 VPWR a_18902_42760# 0.391454f
C1208 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B 3.55251f
C1209 SUNSAR_SAR8B_CV_0.XA4.EN a_11322_28556# 0.135353f
C1210 VPWR SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 16.830301f
C1211 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B 0.419738f
C1212 VPWR SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MP1.S 0.104609f
C1213 uio_oe[0] uio_out[0] 1.55761f
C1214 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1215 a_13950_4742# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.156331f
C1216 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B 0.419738f
C1217 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.14516f
C1218 VPWR a_10190_41000# 0.388224f
C1219 VPWR a_13862_40296# 0.458821f
C1220 VPWR a_16542_2630# 0.448756f
C1221 SUNSAR_SAR8B_CV_0.XA7.ENO SUNSAR_SAR8B_CV_0.XA20.CNO 0.252047f
C1222 VPWR SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 2.7271f
C1223 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 3.55251f
C1224 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.375196f
C1225 VPWR a_18882_31196# 0.44007f
C1226 SUNSAR_CAPT8B_CV_0.XD09.XA5.A SUNSAR_CAPT8B_CV_0.XD09.XA6.A 0.301485f
C1227 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B SUNSAR_SAR8B_CV_0.SARN 27.1615f
C1228 VPWR SUNSAR_CAPT8B_CV_0.XI14.XA7.C 2.97223f
C1229 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B 0.386137f
C1230 VPWR uo_out[0] 1.02382f
C1231 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 54.2165f
C1232 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B 0.441867f
C1233 m3_24750_3728# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.172147f
C1234 VPWR a_13842_30316# 0.404384f
C1235 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XA4.CP0 0.327152f
C1236 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XA20.CNO 0.191868f
C1237 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 0.40569f
C1238 a_12582_4390# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.15559f
C1239 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.174995f
C1240 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.63636f
C1241 VPWR a_3762_31196# 0.44007f
C1242 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.527529f
C1243 a_3762_30316# SUNSAR_SAR8B_CV_0.XA0.XA2.A 0.129098f
C1244 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA4.MP1.S 0.104609f
C1245 VPWR SUNSAR_CAPT8B_CV_0.XH13.XA6.A 1.63909f
C1246 VPWR SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MP1.S 0.104609f
C1247 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN uo_out[0] 0.305166f
C1248 SUNSAR_CAPT8B_CV_0.XA6.A SUNSAR_CAPT8B_CV_0.XA5.XA2.A 0.107823f
C1249 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G 0.145483f
C1250 SUNSAR_CAPT8B_CV_0.XG12.XA7.C uo_out[2] 0.246146f
C1251 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_CAPT8B_CV_0.XD09.XA7.CN 0.241356f
C1252 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XA2.EN 0.491653f
C1253 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 1.2199f
C1254 VPWR a_20250_32076# 0.433941f
C1255 m3_24750_5648# SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B 0.172147f
C1256 VPWR a_23922_36300# 0.472384f
C1257 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA5.CP0 0.722417f
C1258 VPWR SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G 1.05322f
C1259 VPWR a_16542_4918# 0.470354f
C1260 VPWR SUNSAR_SAR8B_CV_0.XA7.ENO 4.77251f
C1261 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA1.XA4.A 0.204048f
C1262 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B ua[0] 0.241597f
C1263 VPWR SUNSAR_SAR8B_CV_0.XA4.XA1.XA4.MP1.S 0.104609f
C1264 VPWR a_3762_33836# 0.409601f
C1265 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B SUNSAR_SAR8B_CV_0.XB2.CKN 0.26479f
C1266 VPWR SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A 2.50679f
C1267 VPWR a_23922_31724# 0.412398f
C1268 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 2.31666f
C1269 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.316693f
C1270 VPWR a_10190_43816# 0.391817f
C1271 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.62403f
C1272 SUNSAR_SAR8B_CV_0.SARN ua[0] 1.02466f
C1273 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G 1.06002f
C1274 SUNSAR_CAPT8B_CV_0.XH13.XA7.C a_18902_41000# 0.15757f
C1275 SUNSAR_CAPT8B_CV_0.XC08.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1276 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B SUNSAR_SAR8B_CV_0.SARN 6.86675f
C1277 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B 3.55251f
C1278 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA20.CPO 0.820808f
C1279 VPWR uo_out[5] 1.02721f
C1280 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.EN 0.152052f
C1281 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.63636f
C1282 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B 3.55251f
C1283 VPWR SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S 0.183853f
C1284 VPWR a_20250_27852# 0.358413f
C1285 VPWR a_9990_5974# 0.451043f
C1286 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G 0.363295f
C1287 VPWR a_15230_40648# 0.493179f
C1288 VPWR a_18882_27148# 0.471462f
C1289 SUNSAR_SAR8B_CV_0.XA2.EN a_6282_28556# 0.135353f
C1290 a_3782_41000# SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.15757f
C1291 SUNSAR_SAR8B_CV_0.XA7.XA9.A SUNSAR_SAR8B_CV_0.XA7.XA9.B 0.527529f
C1292 SUNSAR_CAPT8B_CV_0.XC08.XA6.A a_5150_42760# 0.111734f
C1293 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B 0.437693f
C1294 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 4.0111f
C1295 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> a_3762_33836# 0.103403f
C1296 VPWR a_10170_33836# 0.409601f
C1297 a_13842_33836# SUNSAR_SAR8B_CV_0.XDAC2.CP<2> 0.103403f
C1298 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 3.07164f
C1299 VPWR SUNSAR_SAR8B_CV_0.XA4.XA2.A 2.45309f
C1300 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111173f
C1301 VPWR a_20270_40648# 0.493179f
C1302 SUNSAR_CAPT8B_CV_0.XB07.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1303 VPWR a_13862_43288# 0.394205f
C1304 VPWR a_8802_29612# 0.397362f
C1305 SUNSAR_CAPT8B_CV_0.XC08.XA7.C SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.233892f
C1306 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.22339f
C1307 a_22790_43640# SUNSAR_CAPT8B_CV_0.XA6.XA2.A 0.127669f
C1308 SUNSAR_SAR8B_CV_0.XA3.CN1 SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.702226f
C1309 SUNSAR_SAR8B_CV_0.XA1.CEIN SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.158152f
C1310 VPWR a_8802_31196# 0.44007f
C1311 SUNSAR_CAPT8B_CV_0.XG12.XA6.A SUNSAR_CAPT8B_CV_0.XG12.XA7.CN 0.744161f
C1312 VPWR a_23942_41000# 0.390915f
C1313 VPWR SUNSAR_CAPT8B_CV_0.XA6.B 0.868246f
C1314 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B 0.441867f
C1315 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B 0.40569f
C1316 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.D<1> 3.10225f
C1317 SUNSAR_SAR8B_CV_0.XA4.XA2.A SUNSAR_SAR8B_CV_0.XA4.XA4.A 0.133602f
C1318 SUNSAR_SAR8B_CV_0.XA4.XA9.B SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.205884f
C1319 SUNSAR_CAPT8B_CV_0.XF11.XA7.C uo_out[3] 0.249907f
C1320 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.S 0.138148f
C1321 VPWR a_18882_35948# 0.417826f
C1322 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B SUNSAR_SAR8B_CV_0.SARN 54.2165f
C1323 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA3.MP1.S 0.106927f
C1324 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B 13.6519f
C1325 VPWR SUNSAR_SAR8B_CV_0.XA20.CK_CMP 1.1111f
C1326 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.SARN 0.103734f
C1327 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B 13.6519f
C1328 VPWR SUNSAR_CAPT8B_CV_0.XG12.XA4.MP1.S 0.106927f
C1329 SUNSAR_SAR8B_CV_0.XA4.XA12.A SUNSAR_SAR8B_CV_0.XA5.CEIN 0.158152f
C1330 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.327208f
C1331 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA7.EN 0.291697f
C1332 VPWR a_10190_41880# 0.395781f
C1333 SUNSAR_SAR8B_CV_0.D<0> tt_um_TT06_SAR_done_0.DONE 0.490252f
C1334 VPWR SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G 0.519052f
C1335 SUNSAR_SAR8B_CV_0.XA1.XA11.A a_6282_36300# 0.13402f
C1336 uo_out[4] uo_out[5] 1.16093f
C1337 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.144331f
C1338 VPWR a_8802_35068# 0.394528f
C1339 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA20.XA3.CO 0.137745f
C1340 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.268016f
C1341 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[1] 0.238239f
C1342 VPWR SUNSAR_SAR8B_CV_0.XA3.CEIN 2.30393f
C1343 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 2.18614f
C1344 VPWR a_15210_36300# 0.398846f
C1345 VPWR SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.635621f
C1346 SUNSAR_CAPT8B_CV_0.XC08.QN SUNSAR_CAPT8B_CV_0.XC08.XA7.C 0.318734f
C1347 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 3.39041f
C1348 tt_um_TT06_SAR_done_0.DONE ui_in[0] 0.201929f
C1349 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.412143f
C1350 SUNSAR_SAR8B_CV_0.XA1.XA9.A a_6282_35068# 0.129098f
C1351 VPWR a_20270_41880# 0.395781f
C1352 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.XA1.EN 1.2771f
C1353 SUNSAR_SAR8B_CV_0.XA7.CN1 a_21402_31196# 0.109137f
C1354 VPWR a_13842_35420# 0.39968f
C1355 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA5.XA4.A 0.204048f
C1356 SUNSAR_SAR8B_CV_0.XA3.DONE SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.145738f
C1357 a_3762_35420# VPWR 0.39968f
C1358 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP2.S 0.150467f
C1359 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G 0.145483f
C1360 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.SARN 0.64474f
C1361 a_2630_43816# SUNSAR_CAPT8B_CV_0.XB07.QN 0.127669f
C1362 SUNSAR_SAR8B_CV_0.XB1.XA4.GN SUNSAR_SAR8B_CV_0.SARP 0.263588f
C1363 VPWR a_8822_42760# 0.391454f
C1364 VPWR SUNSAR_CAPT8B_CV_0.XD09.XA6.A 1.63909f
C1365 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<4> 0.180772f
C1366 VPWR a_13842_27500# 0.382189f
C1367 VPWR a_3782_44168# 0.3405f
C1368 SUNSAR_SAR8B_CV_0.XA3.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.109613f
C1369 a_11342_42408# SUNSAR_CAPT8B_CV_0.XE10.XA5.A 0.113479f
C1370 SUNSAR_SAR8B_CV_0.XA3.CEIN SUNSAR_SAR8B_CV_0.XA3.XA12.A 0.293159f
C1371 a_20270_41880# SUNSAR_CAPT8B_CV_0.XI14.XA7.CN 0.100592f
C1372 a_10170_30316# SUNSAR_SAR8B_CV_0.XA3.XA2.A 0.127528f
C1373 VPWR SUNSAR_CAPT8B_CV_0.XF11.XA4.MP1.S 0.106927f
C1374 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.383512f
C1375 uo_out[3] uo_out[2] 0.109993f
C1376 VPWR a_3762_28556# 0.406628f
C1377 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B 27.1615f
C1378 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<7> 2.50324f
C1379 SUNSAR_SAR8B_CV_0.XA2.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<4> 0.738812f
C1380 VPWR a_15210_28204# 0.361706f
C1381 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A 1.62434f
C1382 SUNSAR_SAR8B_CV_0.XA6.EN a_16362_28556# 0.135353f
C1383 VPWR a_18902_42408# 0.391292f
C1384 SUNSAR_SAR8B_CV_0.XA5.XA9.A SUNSAR_SAR8B_CV_0.XA5.XA9.B 0.527529f
C1385 SUNSAR_SAR8B_CV_0.XA5.XA11.A SUNSAR_SAR8B_CV_0.XA5.CEIN 0.352238f
C1386 SUNSAR_CAPT8B_CV_0.XF11.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1387 VPWR uio_out[0] 0.408488f
C1388 a_15210_33836# SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.101833f
C1389 SUNSAR_SAR8B_CV_0.D<3> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1390 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.383512f
C1391 VPWR SUNSAR_SAR8B_CV_0.XA20.XA11.MP1.S 0.106794f
C1392 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.205884f
C1393 VPWR a_9990_5622# 0.470814f
C1394 SUNSAR_SAR8B_CV_0.XA1.XA9.B SUNSAR_SAR8B_CV_0.XA1.XA10.A 0.205884f
C1395 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.CPO 0.11826f
C1396 a_21402_35420# SUNSAR_SAR8B_CV_0.XA7.XA9.A 0.160931f
C1397 VPWR a_5150_41880# 0.395781f
C1398 SUNSAR_CAPT8B_CV_0.XC08.XA7.C uo_out[6] 0.251051f
C1399 VPWR SUNSAR_CAPT8B_CV_0.XI14.QN 0.901631f
C1400 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.303428f
C1401 SUNSAR_SAR8B_CV_0.XA7.EN a_17730_28556# 0.132757f
C1402 SUNSAR_SAR8B_CV_0.EN tt_um_TT06_SAR_done_0.DONE 0.131506f
C1403 VPWR SUNSAR_SAR8B_CV_0.XA4.XA12.A 0.723728f
C1404 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.375196f
C1405 a_20250_33836# SUNSAR_SAR8B_CV_0.XA7.CN0 0.101833f
C1406 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B 0.441867f
C1407 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> SUNSAR_SAR8B_CV_0.XDAC2.CP<5> 0.143675f
C1408 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA7.MP1.S 0.106927f
C1409 a_16382_42408# SUNSAR_CAPT8B_CV_0.XG12.XA5.A 0.113479f
C1410 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN uo_out[6] 0.306905f
C1411 VPWR SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S 0.405511f
C1412 VPWR a_10170_28908# 0.395394f
C1413 VPWR a_5150_41352# 0.394053f
C1414 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A m3_9126_5808# 0.105547f
C1415 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.30589f
C1416 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<6> 0.738798f
C1417 SUNSAR_CAPT8B_CV_0.XI14.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA7.C 0.233892f
C1418 SUNSAR_CAPT8B_CV_0.XD09.XA7.C tt_um_TT06_SAR_done_0.DONE 0.227625f
C1419 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S SUNSAR_SAR8B_CV_0.XB1.CKN 0.669708f
C1420 SUNSAR_SAR8B_CV_0.XA7.XA11.A SUNSAR_SAR8B_CV_0.XA7.CEIN 0.381914f
C1421 VPWR a_16542_2982# 0.490338f
C1422 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.EN 0.11263f
C1423 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA6.A 1.63909f
C1424 VPWR a_20270_41352# 0.394053f
C1425 VPWR a_15210_35948# 0.417826f
C1426 VPWR a_16542_3334# 0.380282f
C1427 VPWR a_13842_35068# 0.394528f
C1428 SUNSAR_CAPT8B_CV_0.XH13.XA7.C SUNSAR_CAPT8B_CV_0.XH13.XA6.A 0.649845f
C1429 VPWR a_20250_29612# 0.398044f
C1430 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.EN 0.952619f
C1431 SUNSAR_SAR8B_CV_0.D<0> SUNSAR_SAR8B_CV_0.XA7.CN1 0.595738f
C1432 VPWR a_23942_41880# 0.398828f
C1433 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.SARN 0.473354f
C1434 VPWR a_5150_43816# 0.391817f
C1435 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA5.A 0.898003f
C1436 SUNSAR_CAPT8B_CV_0.XH13.QN a_17750_43816# 0.127669f
C1437 SUNSAR_CAPT8B_CV_0.XB07.XA5.A SUNSAR_CAPT8B_CV_0.XB07.XA7.CN 0.432466f
C1438 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B 3.55251f
C1439 VPWR a_20250_35068# 0.391458f
C1440 VPWR SUNSAR_SAR8B_CV_0.XA5.XA4.A 2.31184f
C1441 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.257526f
C1442 SUNSAR_SAR8B_CV_0.XA20.CNO SUNSAR_SAR8B_CV_0.XA20.CPO 7.93512f
C1443 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G 0.145483f
C1444 VPWR SUNSAR_SAR8B_CV_0.D<6> 5.43027f
C1445 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.13041f
C1446 SUNSAR_SAR8B_CV_0.XA20.XA9.Y SUNSAR_SAR8B_CV_0.XA20.XA3.N1 0.331207f
C1447 VPWR a_8802_32076# 0.436368f
C1448 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.A 0.722887f
C1449 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B 0.441867f
C1450 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.109613f
C1451 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> SUNSAR_SAR8B_CV_0.XDAC2.CP<4> 3.45828f
C1452 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B SUNSAR_SAR8B_CV_0.SARN 3.57448f
C1453 VPWR a_23942_40296# 0.455498f
C1454 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.596437f
C1455 VPWR SUNSAR_SAR8B_CV_0.XA7.XA1.XA4.MP1.S 0.104609f
C1456 a_12582_5446# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.101033f
C1457 VPWR a_18882_30316# 0.403802f
C1458 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.D<0> 0.315968f
C1459 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.126354f
C1460 VPWR a_10170_27852# 0.358413f
C1461 uo_out[7] SUNSAR_CAPT8B_CV_0.XB07.XA7.C 0.248979f
C1462 VPWR a_8802_30316# 0.404384f
C1463 VPWR SUNSAR_SAR8B_CV_0.XDAC2.CP<0> 4.36162f
C1464 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B 0.441867f
C1465 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN a_12710_42408# 0.100131f
C1466 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.740872f
C1467 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC1.CP<9> 0.268769f
C1468 VPWR a_10170_34716# 0.399819f
C1469 VPWR SUNSAR_SAR8B_CV_0.XA20.CPO 6.88568f
C1470 SUNSAR_CAPT8B_CV_0.XC08.QN uo_out[6] 0.258218f
C1471 SUNSAR_CAPT8B_CV_0.XA5.XA2.A SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.239611f
C1472 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<1> 0.202832f
C1473 SUNSAR_SAR8B_CV_0.EN ui_in[0] 0.968121f
C1474 VPWR a_9990_4566# 0.413433f
C1475 SUNSAR_SAR8B_CV_0.XA20.XA9.Y a_22770_28556# 0.140127f
C1476 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.145339f
C1477 VPWR SUNSAR_SAR8B_CV_0.XA20.XA11.Y 0.658328f
C1478 VPWR a_13862_41352# 0.394053f
C1479 VPWR SUNSAR_CAPT8B_CV_0.XA6.A 1.18734f
C1480 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XDAC2.CP<3> 0.174995f
C1481 VPWR SUNSAR_CAPT8B_CV_0.XC08.XA3.MP1.S 0.106927f
C1482 VPWR SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S 0.183853f
C1483 SUNSAR_SAR8B_CV_0.XA7.CP0 SUNSAR_SAR8B_CV_0.D<0> 0.331282f
C1484 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.XDAC2.CP<8> 0.165965f
C1485 SUNSAR_SAR8B_CV_0.XB1.XA4.GN a_12582_3686# 0.16579f
C1486 a_13842_35420# SUNSAR_SAR8B_CV_0.XA4.XA9.A 0.133834f
C1487 SUNSAR_SAR8B_CV_0.XA3.XA9.A SUNSAR_SAR8B_CV_0.XA3.XA9.B 0.527529f
C1488 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.EN 0.952619f
C1489 VPWR SUNSAR_SAR8B_CV_0.XA5.XA11.MP1.S 0.101979f
C1490 SUNSAR_SAR8B_CV_0.XA20.XA10.Y SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.11382f
C1491 VPWR a_8802_26796# 0.442908f
C1492 SUNSAR_SAR8B_CV_0.XA5.DONE SUNSAR_SAR8B_CV_0.XA5.XA9.A 0.145738f
C1493 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B SUNSAR_SAR8B_CV_0.SARN 13.6523f
C1494 SUNSAR_SAR8B_CV_0.XA6.CEIN SUNSAR_SAR8B_CV_0.XA5.CEIN 0.432008f
C1495 a_2610_36828# SUNSAR_SAR8B_CV_0.XA0.XA12.A 0.10248f
C1496 SUNSAR_CAPT8B_CV_0.XA4.MP1.G clk 0.438597f
C1497 SUNSAR_SAR8B_CV_0.XA5.XA11.A a_16362_36300# 0.13402f
C1498 VPWR a_8822_42408# 0.391292f
C1499 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA6.B 0.254583f
C1500 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<6> 2.2622f
C1501 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MP1.S 0.104609f
C1502 VPWR SUNSAR_CAPT8B_CV_0.XA5.XA1.MP1.S 0.118162f
C1503 a_17730_36300# SUNSAR_SAR8B_CV_0.XA6.XA11.A 0.13253f
C1504 a_11322_31196# SUNSAR_SAR8B_CV_0.XA3.CN1 0.109137f
C1505 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B SUNSAR_SAR8B_CV_0.SARP 27.1615f
C1506 VPWR a_15230_41000# 0.388204f
C1507 VPWR a_15230_43816# 0.391817f
C1508 SUNSAR_SAR8B_CV_0.XA2.EN SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.111217f
C1509 SUNSAR_SAR8B_CV_0.XA4.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.316693f
C1510 SUNSAR_SAR8B_CV_0.XA6.CN1 SUNSAR_SAR8B_CV_0.XA6.XA2.A 0.702226f
C1511 SUNSAR_SAR8B_CV_0.XA7.XA2.A SUNSAR_SAR8B_CV_0.XA7.XA4.A 0.133602f
C1512 a_12690_35948# SUNSAR_SAR8B_CV_0.XA4.XA10.A 0.132671f
C1513 a_22790_41880# SUNSAR_CAPT8B_CV_0.XA6.A 0.111538f
C1514 SUNSAR_SAR8B_CV_0.XA5.XA4.A SUNSAR_SAR8B_CV_0.D<2> 0.228332f
C1515 VPWR SUNSAR_SAR8B_CV_0.XA5.XA9.A 1.2202f
C1516 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW ua[0] 0.453892f
C1517 VPWR a_15210_36828# 0.395582f
C1518 SUNSAR_SAR8B_CV_0.XA1.EN SUNSAR_SAR8B_CV_0.XA20.CNO 1.03107f
C1519 SUNSAR_SAR8B_CV_0.D<6> SUNSAR_SAR8B_CV_0.D<2> 0.200315f
C1520 VPWR a_23942_44344# 0.342053f
C1521 SUNSAR_SAR8B_CV_0.XB2.CKN SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW 0.169642f
C1522 VPWR SUNSAR_CAPT8B_CV_0.XB07.XA3.MP1.S 0.106927f
C1523 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.665724f
C1524 a_21402_36300# SUNSAR_SAR8B_CV_0.XA7.XA11.A 0.13402f
C1525 VPWR SUNSAR_SAR8B_CV_0.XA5.XA10.A 0.779986f
C1526 VPWR SUNSAR_SAR8B_CV_0.XA2.XA1.XA4.MP1.S 0.104609f
C1527 a_5130_30316# SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.127528f
C1528 clk uio_out[0] 0.120689f
C1529 VPWR SUNSAR_SAR8B_CV_0.XA20.XA2.N2 0.337652f
C1530 VPWR SUNSAR_SAR8B_CV_0.XA4.XA11.MP1.S 0.119314f
C1531 SUNSAR_SAR8B_CV_0.XA0.XA4.A SUNSAR_SAR8B_CV_0.XA20.CNO 0.231927f
C1532 VPWR SUNSAR_SAR8B_CV_0.SARP 0.1398f
C1533 VPWR SUNSAR_CAPT8B_CV_0.XF11.QN 0.901622f
C1534 VPWR a_10170_32956# 0.436368f
C1535 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B 0.635098f
C1536 VPWR SUNSAR_SAR8B_CV_0.XA6.XA1.XA4.MP1.S 0.104609f
C1537 VPWR a_16542_5270# 0.489055f
C1538 m3_2358_3728# SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B 0.172147f
C1539 SUNSAR_SAR8B_CV_0.XA7.EN SUNSAR_SAR8B_CV_0.D<1> 0.438277f
C1540 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> SUNSAR_SAR8B_CV_0.D<2> 0.155424f
C1541 VPWR a_15230_41880# 0.395781f
C1542 SUNSAR_SAR8B_CV_0.D<5> SUNSAR_SAR8B_CV_0.D<4> 0.587991f
C1543 SUNSAR_SAR8B_CV_0.SARP SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B 3.55251f
C1544 VPWR a_8822_40296# 0.458821f
C1545 SUNSAR_CAPT8B_CV_0.XA5.B SUNSAR_CAPT8B_CV_0.XA4.MP1.G 0.138433f
C1546 SUNSAR_CAPT8B_CV_0.XG12.XA6.A a_15230_42760# 0.111734f
C1547 VPWR SUNSAR_SAR8B_CV_0.XA1.EN 5.52718f
C1548 a_3762_29612# SUNSAR_SAR8B_CV_0.EN 0.143959f
C1549 SUNSAR_SAR8B_CV_0.SARN SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B 3.55251f
C1550 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> SUNSAR_SAR8B_CV_0.XDAC2.CP<1> 0.26609f
C1551 SUNSAR_SAR8B_CV_0.EN SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G 0.145483f
C1552 SUNSAR_SAR8B_CV_0.D<1> SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.180769f
C1553 SUNSAR_SAR8B_CV_0.XA6.EN SUNSAR_SAR8B_CV_0.XA6.XA4.A 0.129613f
C1554 VPWR a_10170_29612# 0.397362f
C1555 a_13950_4390# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.15559f
C1556 SUNSAR_SAR8B_CV_0.XA5.XA9.B SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.179089f
C1557 SUNSAR_SAR8B_CV_0.XA7.CEIN SUNSAR_SAR8B_CV_0.XA6.XA12.A 0.158152f
C1558 a_2610_32956# SUNSAR_SAR8B_CV_0.XDAC1.CP<8> 0.101124f
C1559 a_11322_35420# SUNSAR_SAR8B_CV_0.XA3.XA9.A 0.160931f
C1560 SUNSAR_SAR8B_CV_0.XA5.XA12.A SUNSAR_SAR8B_CV_0.XA5.CEIN 0.293159f
C1561 VPWR SUNSAR_SAR8B_CV_0.XA0.XA4.A 2.31184f
C1562 a_13950_5094# SUNSAR_SAR8B_CV_0.XB2.TIE_L 0.160184f
C1563 SUNSAR_SAR8B_CV_0.XA1.XA4.A SUNSAR_SAR8B_CV_0.XA1.XA2.A 0.133602f
C1564 uo_out[7] uo_out[6] 2.38922f
C1565 SUNSAR_CAPT8B_CV_0.XH13.XA5.A a_17750_42408# 0.111909f
C1566 VPWR SUNSAR_SAR8B_CV_0.XA4.CP0 2.64055f
C1567 VPWR a_3782_43288# 0.394205f
C1568 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B 0.40569f
C1569 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 0.440586f
C1570 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA20.CPO 0.375025f
C1571 VPWR a_20250_28908# 0.395394f
C1572 SUNSAR_SAR8B_CV_0.D<7> SUNSAR_SAR8B_CV_0.XA20.CPO 0.240612f
C1573 VPWR SUNSAR_SAR8B_CV_0.XA6.CEIN 1.06023f
C1574 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A SUNSAR_SAR8B_CV_0.XB2.CKN 0.143148f
C1575 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N SUNSAR_SAR8B_CV_0.XA4.EN 0.339883f
C1576 SUNSAR_SAR8B_CV_0.XA20.XA12.Y SUNSAR_SAR8B_CV_0.CK_SAMPLE 0.151003f
C1577 VPWR a_3782_40648# 0.491776f
C1578 ua[2] VGND 0.117454f
C1579 ua[3] VGND 0.117454f
C1580 ua[4] VGND 0.118698f
C1581 ua[5] VGND 0.120088f
C1582 ua[6] VGND 0.120088f
C1583 ua[7] VGND 0.111009f
C1584 ua[0] VGND 7.63113f
C1585 ua[1] VGND 7.01035f
C1586 uio_out[0] VGND 8.52142f
C1587 uio_oe[0] VGND 7.87718f
C1588 ui_in[0] VGND 5.4069f
C1589 clk VGND 6.22723f
C1590 uo_out[0] VGND 2.40292f
C1591 uo_out[1] VGND 1.50319f
C1592 uo_out[2] VGND 1.42895f
C1593 uo_out[3] VGND 1.68048f
C1594 uo_out[4] VGND 1.55276f
C1595 uo_out[5] VGND 1.75883f
C1596 uo_out[6] VGND 2.73387f
C1597 uo_out[7] VGND 3.23518f
C1598 VPWR VGND 0.949219p
C1599 TIE_L1 VGND 1.33691f
C1600 TIE_L2 VGND 1.67804f
C1601 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1A.B VGND 6.93682f
C1602 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1A.B VGND 6.93682f
C1603 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES16.B VGND 14.555001f
C1604 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES16.B VGND 14.555001f
C1605 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES2.B VGND 7.335569f
C1606 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES2.B VGND 7.335569f
C1607 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES8.B VGND 10.4697f
C1608 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES8.B VGND 10.4697f
C1609 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES4.B VGND 8.43607f
C1610 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES4.B VGND 8.43607f
C1611 SUNSAR_SAR8B_CV_0.XDAC2.XC1.XRES1B.B VGND 6.67818f
C1612 SUNSAR_SAR8B_CV_0.XDAC1.XC1.XRES1B.B VGND 6.67818f
C1613 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1A.B VGND 6.66914f
C1614 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1A.B VGND 6.66914f
C1615 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES16.B VGND 14.5762f
C1616 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES16.B VGND 14.5762f
C1617 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES2.B VGND 7.33485f
C1618 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES2.B VGND 7.33485f
C1619 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES8.B VGND 10.4697f
C1620 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES8.B VGND 10.4697f
C1621 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES4.B VGND 8.43607f
C1622 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES4.B VGND 8.43607f
C1623 SUNSAR_SAR8B_CV_0.XDAC2.XC32a<0>.XRES1B.B VGND 6.67818f
C1624 SUNSAR_SAR8B_CV_0.XDAC1.XC32a<0>.XRES1B.B VGND 6.67818f
C1625 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1A.B VGND 6.66914f
C1626 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1A.B VGND 6.66914f
C1627 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES16.B VGND 14.5768f
C1628 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES16.B VGND 14.5768f
C1629 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES2.B VGND 7.33485f
C1630 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES2.B VGND 7.33485f
C1631 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES8.B VGND 10.4697f
C1632 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES8.B VGND 10.4697f
C1633 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES4.B VGND 8.43607f
C1634 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES4.B VGND 8.43607f
C1635 SUNSAR_SAR8B_CV_0.XDAC2.X16ab.XRES1B.B VGND 6.67818f
C1636 SUNSAR_SAR8B_CV_0.XDAC1.X16ab.XRES1B.B VGND 6.67818f
C1637 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1A.B VGND 6.66914f
C1638 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1A.B VGND 6.66914f
C1639 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES16.B VGND 14.5735f
C1640 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES16.B VGND 14.5735f
C1641 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES2.B VGND 7.33485f
C1642 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES2.B VGND 7.33485f
C1643 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES8.B VGND 10.472599f
C1644 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES8.B VGND 10.472599f
C1645 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES4.B VGND 8.44055f
C1646 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES4.B VGND 8.44327f
C1647 SUNSAR_SAR8B_CV_0.XDAC2.XC0.XRES1B.B VGND 7.38664f
C1648 SUNSAR_SAR8B_CV_0.XDAC1.XC0.XRES1B.B VGND 7.3834f
C1649 a_15390_2630# VGND 0.543325f $ **FLOATING
C1650 a_13950_2630# VGND 0.428911f $ **FLOATING
C1651 a_12582_2630# VGND 0.428496f $ **FLOATING
C1652 a_11142_2630# VGND 0.544481f $ **FLOATING
C1653 a_15390_2982# VGND 0.492315f $ **FLOATING
C1654 a_13950_2982# VGND 0.352955f $ **FLOATING
C1655 a_12582_2982# VGND 0.352955f $ **FLOATING
C1656 a_11142_2982# VGND 0.490744f $ **FLOATING
C1657 a_15390_3334# VGND 0.375184f $ **FLOATING
C1658 a_13950_3334# VGND 0.352694f $ **FLOATING
C1659 a_12582_3334# VGND 0.352694f $ **FLOATING
C1660 a_11142_3334# VGND 0.375184f $ **FLOATING
C1661 a_13950_3686# VGND 0.352463f $ **FLOATING
C1662 a_12582_3686# VGND 0.352463f $ **FLOATING
C1663 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.B VGND 41.754498f
C1664 SUNSAR_SAR8B_CV_0.XB2.XA3.MP0.S VGND 0.702101f
C1665 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.B VGND 41.754498f
C1666 SUNSAR_SAR8B_CV_0.XB1.XA3.MP0.S VGND 0.702101f
C1667 a_15390_4038# VGND 0.397033f $ **FLOATING
C1668 a_13950_4038# VGND 0.354407f $ **FLOATING
C1669 a_12582_4038# VGND 0.354407f $ **FLOATING
C1670 a_11142_4038# VGND 0.397033f $ **FLOATING
C1671 SUNSAR_SAR8B_CV_0.XB2.XCAPB1.A VGND 37.790997f
C1672 SUNSAR_SAR8B_CV_0.XB2.CKN VGND 2.38663f
C1673 SUNSAR_SAR8B_CV_0.XB2.XA4.MN1.S VGND 0.103625f
C1674 a_13950_4390# VGND 0.352432f $ **FLOATING
C1675 a_12582_4390# VGND 0.352432f $ **FLOATING
C1676 SUNSAR_SAR8B_CV_0.XB1.XA4.MN1.S VGND 0.103625f
C1677 SUNSAR_SAR8B_CV_0.XB1.CKN VGND 2.38663f
C1678 SUNSAR_SAR8B_CV_0.XB1.XCAPB1.A VGND 37.790997f
C1679 SUNSAR_SAR8B_CV_0.XB2.XA4.GN VGND 3.12067f
C1680 a_15390_4566# VGND 0.389036f $ **FLOATING
C1681 SUNSAR_SAR8B_CV_0.XB1.XA4.GN VGND 3.08351f
C1682 a_11142_4566# VGND 0.389036f $ **FLOATING
C1683 SUNSAR_SAR8B_CV_0.XB2.XA4.TIE_H VGND 0.970036f
C1684 a_13950_4742# VGND 0.352456f $ **FLOATING
C1685 a_12582_4742# VGND 0.352456f $ **FLOATING
C1686 SUNSAR_SAR8B_CV_0.XB2.XA1.MP0.G VGND 0.7964f
C1687 a_15390_4918# VGND 0.470144f $ **FLOATING
C1688 SUNSAR_SAR8B_CV_0.XB1.XA1.MP0.G VGND 0.7964f
C1689 SUNSAR_SAR8B_CV_0.XB1.XA4.TIE_H VGND 0.970036f
C1690 a_11142_4918# VGND 0.471715f $ **FLOATING
C1691 a_13950_5094# VGND 0.353103f $ **FLOATING
C1692 a_12582_5094# VGND 0.353103f $ **FLOATING
C1693 a_15390_5270# VGND 0.492927f $ **FLOATING
C1694 a_11142_5270# VGND 0.491356f $ **FLOATING
C1695 SUNSAR_SAR8B_CV_0.XB2.XA2.MP0.G VGND 0.596866f
C1696 a_13950_5446# VGND 0.433341f $ **FLOATING
C1697 a_12582_5446# VGND 0.433756f $ **FLOATING
C1698 a_15390_5622# VGND 0.47219f $ **FLOATING
C1699 a_15390_5974# VGND 0.541341f $ **FLOATING
C1700 SUNSAR_SAR8B_CV_0.XB1.XA2.MP0.G VGND 0.596866f
C1701 a_11142_5622# VGND 0.47376f $ **FLOATING
C1702 a_11142_5974# VGND 0.540186f $ **FLOATING
C1703 a_22770_26796# VGND 0.529341f $ **FLOATING
C1704 a_21402_26796# VGND 0.531659f $ **FLOATING
C1705 a_17730_26796# VGND 0.530834f $ **FLOATING
C1706 a_16362_26796# VGND 0.531989f $ **FLOATING
C1707 a_12690_26796# VGND 0.530834f $ **FLOATING
C1708 a_11322_26796# VGND 0.531989f $ **FLOATING
C1709 a_7650_26796# VGND 0.530213f $ **FLOATING
C1710 a_6282_26796# VGND 0.530979f $ **FLOATING
C1711 a_2610_26796# VGND 0.531666f $ **FLOATING
C1712 a_22770_27148# VGND 0.499848f $ **FLOATING
C1713 a_21402_27148# VGND 0.467094f $ **FLOATING
C1714 a_17730_27148# VGND 0.471508f $ **FLOATING
C1715 a_16362_27148# VGND 0.467722f $ **FLOATING
C1716 a_12690_27148# VGND 0.471508f $ **FLOATING
C1717 a_11322_27148# VGND 0.467722f $ **FLOATING
C1718 a_7650_27148# VGND 0.470266f $ **FLOATING
C1719 a_6282_27148# VGND 0.465734f $ **FLOATING
C1720 a_2610_27148# VGND 0.471719f $ **FLOATING
C1721 a_21402_27500# VGND 0.385968f $ **FLOATING
C1722 a_17730_27500# VGND 0.387712f $ **FLOATING
C1723 a_16362_27500# VGND 0.386249f $ **FLOATING
C1724 a_12690_27500# VGND 0.387712f $ **FLOATING
C1725 a_11322_27500# VGND 0.386249f $ **FLOATING
C1726 a_7650_27500# VGND 0.38671f $ **FLOATING
C1727 a_6282_27500# VGND 0.384229f $ **FLOATING
C1728 a_2610_27500# VGND 0.387692f $ **FLOATING
C1729 a_21402_27852# VGND 0.370125f $ **FLOATING
C1730 a_17730_27852# VGND 0.370785f $ **FLOATING
C1731 a_16362_27852# VGND 0.368771f $ **FLOATING
C1732 a_12690_27852# VGND 0.370785f $ **FLOATING
C1733 a_11322_27852# VGND 0.368771f $ **FLOATING
C1734 a_7650_27852# VGND 0.369543f $ **FLOATING
C1735 a_6282_27852# VGND 0.366751f $ **FLOATING
C1736 a_2610_27852# VGND 0.370525f $ **FLOATING
C1737 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MN2.S VGND 0.506947f
C1738 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MN2.S VGND 0.502211f
C1739 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MN2.S VGND 0.477244f
C1740 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MN2.S VGND 0.502211f
C1741 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MN2.S VGND 0.477244f
C1742 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MN2.S VGND 0.502211f
C1743 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MN2.S VGND 0.477244f
C1744 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MN2.S VGND 0.502211f
C1745 a_21402_28204# VGND 0.405715f $ **FLOATING
C1746 a_17730_28204# VGND 0.406284f $ **FLOATING
C1747 a_16362_28204# VGND 0.406284f $ **FLOATING
C1748 a_12690_28204# VGND 0.406284f $ **FLOATING
C1749 a_11322_28204# VGND 0.406284f $ **FLOATING
C1750 a_7650_28204# VGND 0.405133f $ **FLOATING
C1751 a_6282_28204# VGND 0.404355f $ **FLOATING
C1752 a_2610_28204# VGND 0.406115f $ **FLOATING
C1753 SUNSAR_SAR8B_CV_0.XA20.XA1.MP0.S VGND 0.609217f
C1754 SUNSAR_SAR8B_CV_0.XA7.XA1.XA1.MP3.G VGND 0.741242f
C1755 SUNSAR_SAR8B_CV_0.XA6.XA1.XA1.MP3.G VGND 0.749251f
C1756 SUNSAR_SAR8B_CV_0.XA5.XA1.XA1.MP3.G VGND 0.735502f
C1757 SUNSAR_SAR8B_CV_0.XA4.XA1.XA1.MP3.G VGND 0.749251f
C1758 SUNSAR_SAR8B_CV_0.XA3.XA1.XA1.MP3.G VGND 0.735502f
C1759 SUNSAR_SAR8B_CV_0.XA2.XA1.XA1.MP3.G VGND 0.746591f
C1760 SUNSAR_SAR8B_CV_0.XA1.XA1.XA1.MP3.G VGND 0.73057f
C1761 SUNSAR_SAR8B_CV_0.XA0.XA1.XA1.MP3.G VGND 0.749198f
C1762 a_22770_28556# VGND 0.401649f $ **FLOATING
C1763 a_21402_28556# VGND 0.387558f $ **FLOATING
C1764 a_17730_28556# VGND 0.388127f $ **FLOATING
C1765 a_16362_28556# VGND 0.388127f $ **FLOATING
C1766 a_12690_28556# VGND 0.388127f $ **FLOATING
C1767 a_11322_28556# VGND 0.388127f $ **FLOATING
C1768 a_7650_28556# VGND 0.386976f $ **FLOATING
C1769 a_6282_28556# VGND 0.386198f $ **FLOATING
C1770 a_2610_28556# VGND 0.387958f $ **FLOATING
C1771 a_21402_28908# VGND 0.394283f $ **FLOATING
C1772 a_17730_28908# VGND 0.394852f $ **FLOATING
C1773 a_16362_28908# VGND 0.394852f $ **FLOATING
C1774 a_12690_28908# VGND 0.394852f $ **FLOATING
C1775 a_11322_28908# VGND 0.394852f $ **FLOATING
C1776 a_7650_28908# VGND 0.393701f $ **FLOATING
C1777 a_6282_28908# VGND 0.392923f $ **FLOATING
C1778 a_2610_28908# VGND 0.394683f $ **FLOATING
C1779 SUNSAR_SAR8B_CV_0.SARP VGND 70.1062f
C1780 a_21402_29612# VGND 0.395457f $ **FLOATING
C1781 a_17730_29612# VGND 0.396116f $ **FLOATING
C1782 a_16362_29612# VGND 0.395588f $ **FLOATING
C1783 a_12690_29612# VGND 0.396116f $ **FLOATING
C1784 a_11322_29612# VGND 0.395588f $ **FLOATING
C1785 a_7650_29612# VGND 0.394965f $ **FLOATING
C1786 a_6282_29612# VGND 0.393746f $ **FLOATING
C1787 a_2610_29612# VGND 0.395941f $ **FLOATING
C1788 SUNSAR_SAR8B_CV_0.XA20.XA2.N2 VGND 0.318943f
C1789 a_22770_29964# VGND 0.400512f $ **FLOATING
C1790 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.MN1.S VGND 0.103281f
C1791 SUNSAR_SAR8B_CV_0.XA7.XA1.XA5.LCK_N VGND 1.27143f
C1792 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.MN1.S VGND 0.100021f
C1793 SUNSAR_SAR8B_CV_0.XA6.XA1.XA5.LCK_N VGND 1.26503f
C1794 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.MN1.S VGND 0.100021f
C1795 SUNSAR_SAR8B_CV_0.XA5.XA1.XA5.LCK_N VGND 1.26391f
C1796 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.MN1.S VGND 0.100021f
C1797 SUNSAR_SAR8B_CV_0.XA4.XA1.XA5.LCK_N VGND 1.26503f
C1798 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.MN1.S VGND 0.100021f
C1799 SUNSAR_SAR8B_CV_0.XA3.XA1.XA5.LCK_N VGND 1.26391f
C1800 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.MN1.S VGND 0.100021f
C1801 SUNSAR_SAR8B_CV_0.XA2.XA1.XA5.LCK_N VGND 1.25938f
C1802 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.MN1.S VGND 0.100021f
C1803 SUNSAR_SAR8B_CV_0.XA1.XA1.XA5.LCK_N VGND 1.25329f
C1804 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.MN1.S VGND 0.100021f
C1805 SUNSAR_SAR8B_CV_0.XA0.XA1.XA5.LCK_N VGND 1.26416f
C1806 a_21402_30316# VGND 0.401758f $ **FLOATING
C1807 a_17730_30316# VGND 0.401074f $ **FLOATING
C1808 a_16362_30316# VGND 0.401074f $ **FLOATING
C1809 a_12690_30316# VGND 0.401074f $ **FLOATING
C1810 a_11322_30316# VGND 0.401074f $ **FLOATING
C1811 a_7650_30316# VGND 0.399923f $ **FLOATING
C1812 a_6282_30316# VGND 0.399145f $ **FLOATING
C1813 a_2610_30316# VGND 0.401161f $ **FLOATING
C1814 SUNSAR_SAR8B_CV_0.XA20.CPO VGND 15.3143f
C1815 a_22770_30844# VGND 0.421853f $ **FLOATING
C1816 SUNSAR_SAR8B_CV_0.XA7.XA2.A VGND 2.24318f
C1817 SUNSAR_SAR8B_CV_0.XA6.XA2.A VGND 2.22194f
C1818 SUNSAR_SAR8B_CV_0.XA5.XA2.A VGND 2.22198f
C1819 SUNSAR_SAR8B_CV_0.XA4.XA2.A VGND 2.22194f
C1820 SUNSAR_SAR8B_CV_0.XA3.XA2.A VGND 2.22198f
C1821 SUNSAR_SAR8B_CV_0.XA2.XA2.A VGND 2.20909f
C1822 SUNSAR_SAR8B_CV_0.XA1.XA2.A VGND 2.19751f
C1823 SUNSAR_SAR8B_CV_0.XA0.XA2.A VGND 2.22015f
C1824 a_21402_31196# VGND 0.4255f $ **FLOATING
C1825 a_17730_31196# VGND 0.426069f $ **FLOATING
C1826 a_16362_31196# VGND 0.426069f $ **FLOATING
C1827 a_12690_31196# VGND 0.426069f $ **FLOATING
C1828 a_11322_31196# VGND 0.426069f $ **FLOATING
C1829 a_7650_31196# VGND 0.424917f $ **FLOATING
C1830 a_6282_31196# VGND 0.42414f $ **FLOATING
C1831 a_2610_31196# VGND 0.426156f $ **FLOATING
C1832 SUNSAR_SAR8B_CV_0.XA20.CNO VGND 19.477f
C1833 a_22770_31724# VGND 0.423601f $ **FLOATING
C1834 SUNSAR_SAR8B_CV_0.XA7.CN1 VGND 2.99939f
C1835 SUNSAR_SAR8B_CV_0.XA6.CN1 VGND 2.97987f
C1836 SUNSAR_SAR8B_CV_0.XA5.CN1 VGND 2.97901f
C1837 SUNSAR_SAR8B_CV_0.XA4.CN1 VGND 2.97987f
C1838 SUNSAR_SAR8B_CV_0.XA3.CN1 VGND 2.97901f
C1839 SUNSAR_SAR8B_CV_0.XDAC2.CP<5> VGND 8.85828f
C1840 SUNSAR_SAR8B_CV_0.XDAC2.CP<7> VGND 8.37577f
C1841 a_21402_32076# VGND 0.426091f $ **FLOATING
C1842 a_17730_32076# VGND 0.42666f $ **FLOATING
C1843 a_16362_32076# VGND 0.42666f $ **FLOATING
C1844 a_12690_32076# VGND 0.42666f $ **FLOATING
C1845 a_11322_32076# VGND 0.42666f $ **FLOATING
C1846 a_7650_32076# VGND 0.42666f $ **FLOATING
C1847 a_6282_32076# VGND 0.42666f $ **FLOATING
C1848 a_2610_32076# VGND 0.426748f $ **FLOATING
C1849 SUNSAR_SAR8B_CV_0.XA20.XA3.N1 VGND 1.5559f
C1850 SUNSAR_SAR8B_CV_0.XA20.XA3.N2 VGND 0.328276f
C1851 SUNSAR_SAR8B_CV_0.XA7.XA4.A VGND 3.19736f
C1852 SUNSAR_SAR8B_CV_0.XA6.XA4.A VGND 3.22974f
C1853 SUNSAR_SAR8B_CV_0.XA5.XA4.A VGND 3.22835f
C1854 SUNSAR_SAR8B_CV_0.XA4.XA4.A VGND 3.22974f
C1855 SUNSAR_SAR8B_CV_0.XA3.XA4.A VGND 3.22835f
C1856 SUNSAR_SAR8B_CV_0.XA2.XA4.A VGND 3.22678f
C1857 SUNSAR_SAR8B_CV_0.XA1.XA4.A VGND 3.22545f
C1858 SUNSAR_SAR8B_CV_0.XA0.XA4.A VGND 3.31226f
C1859 SUNSAR_SAR8B_CV_0.XA20.XA3.VMR VGND 2.68984f
C1860 a_21402_32956# VGND 0.426069f $ **FLOATING
C1861 a_17730_32956# VGND 0.426069f $ **FLOATING
C1862 a_16362_32956# VGND 0.426069f $ **FLOATING
C1863 a_12690_32956# VGND 0.426069f $ **FLOATING
C1864 a_11322_32956# VGND 0.426069f $ **FLOATING
C1865 a_7650_32956# VGND 0.426069f $ **FLOATING
C1866 a_6282_32956# VGND 0.426069f $ **FLOATING
C1867 a_2610_32956# VGND 0.426316f $ **FLOATING
C1868 SUNSAR_SAR8B_CV_0.XA20.XA3.CO VGND 2.84889f
C1869 a_22770_33132# VGND 0.403395f $ **FLOATING
C1870 SUNSAR_SAR8B_CV_0.XA7.CP0 VGND 3.01164f
C1871 SUNSAR_SAR8B_CV_0.XA6.CP0 VGND 3.01628f
C1872 SUNSAR_SAR8B_CV_0.XA5.CP0 VGND 3.01641f
C1873 SUNSAR_SAR8B_CV_0.XA4.CP0 VGND 3.01628f
C1874 SUNSAR_SAR8B_CV_0.XA3.CP0 VGND 3.01641f
C1875 SUNSAR_SAR8B_CV_0.XDAC1.CP<4> VGND 5.54669f
C1876 SUNSAR_SAR8B_CV_0.XDAC1.CP<6> VGND 5.78758f
C1877 SUNSAR_SAR8B_CV_0.XDAC1.CP<8> VGND 12.1081f
C1878 a_21402_33836# VGND 0.426756f $ **FLOATING
C1879 a_17730_33836# VGND 0.426756f $ **FLOATING
C1880 a_16362_33836# VGND 0.426756f $ **FLOATING
C1881 a_12690_33836# VGND 0.426756f $ **FLOATING
C1882 a_11322_33836# VGND 0.426756f $ **FLOATING
C1883 a_7650_33836# VGND 0.426756f $ **FLOATING
C1884 a_6282_33836# VGND 0.426756f $ **FLOATING
C1885 a_2610_33836# VGND 0.42696f $ **FLOATING
C1886 SUNSAR_SAR8B_CV_0.SARN VGND 71.1677f
C1887 SUNSAR_SAR8B_CV_0.XA7.XA6.MN1.S VGND 0.149691f
C1888 SUNSAR_SAR8B_CV_0.XA20.XA4.MP0.S VGND 0.515646f
C1889 SUNSAR_SAR8B_CV_0.XA7.CN0 VGND 0.650909f
C1890 SUNSAR_SAR8B_CV_0.XA6.XA6.MN1.S VGND 0.149691f
C1891 SUNSAR_SAR8B_CV_0.XDAC2.CP<0> VGND 5.72791f
C1892 a_22770_34540# VGND 0.39377f $ **FLOATING
C1893 SUNSAR_SAR8B_CV_0.XA7.XA6.MN3.S VGND 0.102f
C1894 SUNSAR_SAR8B_CV_0.XA5.XA6.MN1.S VGND 0.149691f
C1895 SUNSAR_SAR8B_CV_0.XDAC2.CP<1> VGND 4.1719f
C1896 SUNSAR_SAR8B_CV_0.XA4.XA6.MN1.S VGND 0.149691f
C1897 SUNSAR_SAR8B_CV_0.XDAC2.CP<2> VGND 3.27991f
C1898 SUNSAR_SAR8B_CV_0.XA6.XA6.MN3.S VGND 0.102f
C1899 SUNSAR_SAR8B_CV_0.XA5.XA6.MN3.S VGND 0.102f
C1900 SUNSAR_SAR8B_CV_0.XA3.XA6.MN1.S VGND 0.149691f
C1901 SUNSAR_SAR8B_CV_0.XDAC2.CP<3> VGND 4.31299f
C1902 SUNSAR_SAR8B_CV_0.XA2.XA6.MN1.S VGND 0.149691f
C1903 SUNSAR_SAR8B_CV_0.XDAC2.CP<4> VGND 3.68294f
C1904 SUNSAR_SAR8B_CV_0.XA4.XA6.MN3.S VGND 0.102f
C1905 SUNSAR_SAR8B_CV_0.XA3.XA6.MN3.S VGND 0.102f
C1906 SUNSAR_SAR8B_CV_0.XA1.XA6.MN1.S VGND 0.149691f
C1907 SUNSAR_SAR8B_CV_0.XDAC2.CP<6> VGND 4.25175f
C1908 SUNSAR_SAR8B_CV_0.XA0.XA6.MN1.S VGND 0.149988f
C1909 SUNSAR_SAR8B_CV_0.XDAC2.CP<8> VGND 10.151099f
C1910 SUNSAR_SAR8B_CV_0.XA2.XA6.MN3.S VGND 0.102f
C1911 SUNSAR_SAR8B_CV_0.XA1.XA6.MN3.S VGND 0.102f
C1912 SUNSAR_SAR8B_CV_0.XA0.XA6.MN3.S VGND 0.102353f
C1913 SUNSAR_SAR8B_CV_0.XDAC1.CP<9> VGND 8.127279f
C1914 a_21402_34716# VGND 0.39476f $ **FLOATING
C1915 a_17730_34716# VGND 0.39476f $ **FLOATING
C1916 a_16362_34716# VGND 0.39476f $ **FLOATING
C1917 a_12690_34716# VGND 0.39476f $ **FLOATING
C1918 a_11322_34716# VGND 0.39476f $ **FLOATING
C1919 a_7650_34716# VGND 0.39476f $ **FLOATING
C1920 a_6282_34716# VGND 0.39476f $ **FLOATING
C1921 a_2610_34716# VGND 0.394847f $ **FLOATING
C1922 SUNSAR_SAR8B_CV_0.XA20.XA9.Y VGND 4.75786f
C1923 a_22770_34892# VGND 0.394644f $ **FLOATING
C1924 SUNSAR_SAR8B_CV_0.XA7.ENO VGND 1.67603f
C1925 SUNSAR_SAR8B_CV_0.XA7.EN VGND 4.51439f
C1926 SUNSAR_SAR8B_CV_0.XA6.EN VGND 4.46191f
C1927 SUNSAR_SAR8B_CV_0.XA5.EN VGND 4.27708f
C1928 SUNSAR_SAR8B_CV_0.XA4.EN VGND 4.50282f
C1929 SUNSAR_SAR8B_CV_0.XA3.EN VGND 4.42572f
C1930 SUNSAR_SAR8B_CV_0.XA2.EN VGND 4.44437f
C1931 SUNSAR_SAR8B_CV_0.XA1.EN VGND 4.39269f
C1932 a_21402_35068# VGND 0.389563f $ **FLOATING
C1933 a_17730_35068# VGND 0.389563f $ **FLOATING
C1934 a_16362_35068# VGND 0.389563f $ **FLOATING
C1935 a_12690_35068# VGND 0.389563f $ **FLOATING
C1936 a_11322_35068# VGND 0.389563f $ **FLOATING
C1937 a_7650_35068# VGND 0.389563f $ **FLOATING
C1938 a_6282_35068# VGND 0.389563f $ **FLOATING
C1939 a_2610_35068# VGND 0.389651f $ **FLOATING
C1940 SUNSAR_SAR8B_CV_0.XA20.XA10.Y VGND 4.5454f
C1941 SUNSAR_SAR8B_CV_0.XA6.DONE VGND 0.544956f
C1942 SUNSAR_SAR8B_CV_0.XA5.DONE VGND 0.534184f
C1943 SUNSAR_SAR8B_CV_0.XA4.DONE VGND 0.544956f
C1944 SUNSAR_SAR8B_CV_0.XA3.DONE VGND 0.534184f
C1945 SUNSAR_SAR8B_CV_0.XA2.DONE VGND 0.544956f
C1946 SUNSAR_SAR8B_CV_0.XA1.DONE VGND 0.534184f
C1947 SUNSAR_SAR8B_CV_0.XA0.DONE VGND 0.557089f
C1948 a_22770_35420# VGND 0.395535f $ **FLOATING
C1949 a_21402_35420# VGND 0.389041f $ **FLOATING
C1950 a_17730_35420# VGND 0.388925f $ **FLOATING
C1951 a_16362_35420# VGND 0.389297f $ **FLOATING
C1952 a_12690_35420# VGND 0.388925f $ **FLOATING
C1953 a_11322_35420# VGND 0.389297f $ **FLOATING
C1954 a_7650_35420# VGND 0.388925f $ **FLOATING
C1955 a_6282_35420# VGND 0.389297f $ **FLOATING
C1956 a_2610_35420# VGND 0.389228f $ **FLOATING
C1957 SUNSAR_SAR8B_CV_0.XA20.XA11.Y VGND 1.07774f
C1958 SUNSAR_SAR8B_CV_0.XA7.XA9.MN1.S VGND 0.112889f
C1959 SUNSAR_SAR8B_CV_0.XA7.XA9.A VGND 1.50901f
C1960 SUNSAR_SAR8B_CV_0.XA7.XA9.B VGND 1.53168f
C1961 SUNSAR_SAR8B_CV_0.XA6.XA9.A VGND 1.50964f
C1962 SUNSAR_SAR8B_CV_0.XA6.XA9.MN1.S VGND 0.112889f
C1963 SUNSAR_SAR8B_CV_0.XA6.XA9.B VGND 1.54335f
C1964 SUNSAR_SAR8B_CV_0.XA5.XA9.MN1.S VGND 0.112889f
C1965 SUNSAR_SAR8B_CV_0.XA5.XA9.A VGND 1.51005f
C1966 SUNSAR_SAR8B_CV_0.XA5.XA9.B VGND 1.53305f
C1967 SUNSAR_SAR8B_CV_0.XA4.XA9.A VGND 1.50964f
C1968 SUNSAR_SAR8B_CV_0.XA4.XA9.MN1.S VGND 0.112889f
C1969 SUNSAR_SAR8B_CV_0.XA4.XA9.B VGND 1.54335f
C1970 SUNSAR_SAR8B_CV_0.XA3.XA9.MN1.S VGND 0.112889f
C1971 SUNSAR_SAR8B_CV_0.XA3.XA9.A VGND 1.51005f
C1972 SUNSAR_SAR8B_CV_0.XA3.XA9.B VGND 1.53305f
C1973 SUNSAR_SAR8B_CV_0.XA2.XA9.A VGND 1.50964f
C1974 SUNSAR_SAR8B_CV_0.XA2.XA9.MN1.S VGND 0.112889f
C1975 SUNSAR_SAR8B_CV_0.XA2.XA9.B VGND 1.54335f
C1976 SUNSAR_SAR8B_CV_0.XA1.XA9.MN1.S VGND 0.112889f
C1977 SUNSAR_SAR8B_CV_0.XA1.XA9.A VGND 1.51005f
C1978 SUNSAR_SAR8B_CV_0.XA1.XA9.B VGND 1.53305f
C1979 SUNSAR_SAR8B_CV_0.XA0.XA9.A VGND 1.52043f
C1980 SUNSAR_SAR8B_CV_0.XA0.XA9.MN1.S VGND 0.112889f
C1981 SUNSAR_SAR8B_CV_0.XA0.XA9.B VGND 1.61547f
C1982 a_22770_35948# VGND 0.414038f $ **FLOATING
C1983 a_21402_35948# VGND 0.390722f $ **FLOATING
C1984 a_17730_35948# VGND 0.391291f $ **FLOATING
C1985 a_16362_35948# VGND 0.391291f $ **FLOATING
C1986 a_12690_35948# VGND 0.391291f $ **FLOATING
C1987 a_11322_35948# VGND 0.391291f $ **FLOATING
C1988 a_7650_35948# VGND 0.391291f $ **FLOATING
C1989 a_6282_35948# VGND 0.391291f $ **FLOATING
C1990 a_2610_35948# VGND 0.391539f $ **FLOATING
C1991 SUNSAR_SAR8B_CV_0.XA20.XA12.Y VGND 0.79133f
C1992 SUNSAR_SAR8B_CV_0.XA7.XA10.A VGND 0.882731f
C1993 SUNSAR_SAR8B_CV_0.XA6.XA10.A VGND 0.884425f
C1994 SUNSAR_SAR8B_CV_0.XA5.XA10.A VGND 0.884504f
C1995 SUNSAR_SAR8B_CV_0.XA4.XA10.A VGND 0.884425f
C1996 SUNSAR_SAR8B_CV_0.XA3.XA10.A VGND 0.884504f
C1997 SUNSAR_SAR8B_CV_0.XA2.XA10.A VGND 0.884425f
C1998 SUNSAR_SAR8B_CV_0.XA1.XA10.A VGND 0.884504f
C1999 SUNSAR_SAR8B_CV_0.XA0.XA10.A VGND 0.896463f
C2000 a_22770_36300# VGND 0.472701f $ **FLOATING
C2001 a_21402_36300# VGND 0.393831f $ **FLOATING
C2002 a_17730_36300# VGND 0.394738f $ **FLOATING
C2003 a_16362_36300# VGND 0.3944f $ **FLOATING
C2004 a_12690_36300# VGND 0.394718f $ **FLOATING
C2005 a_11322_36300# VGND 0.3944f $ **FLOATING
C2006 a_7650_36300# VGND 0.394715f $ **FLOATING
C2007 a_6282_36300# VGND 0.3944f $ **FLOATING
C2008 a_2610_36300# VGND 0.394963f $ **FLOATING
C2009 a_22770_36652# VGND 0.542519f $ **FLOATING
C2010 SUNSAR_SAR8B_CV_0.XA7.XA11.A VGND 0.882078f
C2011 SUNSAR_SAR8B_CV_0.XA6.XA11.A VGND 0.885089f
C2012 SUNSAR_SAR8B_CV_0.XA5.XA11.A VGND 0.877233f
C2013 SUNSAR_SAR8B_CV_0.XA4.XA11.A VGND 0.885067f
C2014 SUNSAR_SAR8B_CV_0.XA3.XA11.A VGND 0.877221f
C2015 SUNSAR_SAR8B_CV_0.XA2.XA11.A VGND 0.885066f
C2016 SUNSAR_SAR8B_CV_0.XA1.XA11.A VGND 0.877233f
C2017 SUNSAR_SAR8B_CV_0.XA0.XA11.A VGND 0.894319f
C2018 SUNSAR_SAR8B_CV_0.XB2.TIE_L VGND 30.4079f
C2019 a_21402_36828# VGND 0.414394f $ **FLOATING
C2020 a_17730_36828# VGND 0.414304f $ **FLOATING
C2021 a_16362_36828# VGND 0.414011f $ **FLOATING
C2022 a_12690_36828# VGND 0.414294f $ **FLOATING
C2023 a_11322_36828# VGND 0.414011f $ **FLOATING
C2024 a_7650_36828# VGND 0.414296f $ **FLOATING
C2025 a_6282_36828# VGND 0.414011f $ **FLOATING
C2026 a_2610_36828# VGND 0.414386f $ **FLOATING
C2027 SUNSAR_SAR8B_CV_0.XA7.XA12.A VGND 1.08827f
C2028 SUNSAR_SAR8B_CV_0.XA20.CK_CMP VGND 2.06522f
C2029 SUNSAR_SAR8B_CV_0.XA6.XA12.A VGND 1.11123f
C2030 SUNSAR_SAR8B_CV_0.XA7.CEIN VGND 1.46079f
C2031 SUNSAR_SAR8B_CV_0.XA5.XA12.A VGND 1.07013f
C2032 SUNSAR_SAR8B_CV_0.XA6.CEIN VGND 1.71822f
C2033 SUNSAR_SAR8B_CV_0.XA4.XA12.A VGND 1.11118f
C2034 SUNSAR_SAR8B_CV_0.XA5.CEIN VGND 1.53183f
C2035 SUNSAR_SAR8B_CV_0.XA3.XA12.A VGND 1.07013f
C2036 SUNSAR_SAR8B_CV_0.XA4.CEIN VGND 1.7182f
C2037 SUNSAR_SAR8B_CV_0.XA2.XA12.A VGND 1.11119f
C2038 SUNSAR_SAR8B_CV_0.XA3.CEIN VGND 1.53184f
C2039 SUNSAR_SAR8B_CV_0.XA1.XA12.A VGND 1.07013f
C2040 SUNSAR_SAR8B_CV_0.XA2.CEIN VGND 1.7182f
C2041 SUNSAR_SAR8B_CV_0.XA0.XA12.A VGND 1.12334f
C2042 SUNSAR_SAR8B_CV_0.XA1.CEIN VGND 1.53659f
C2043 a_21402_37180# VGND 0.475717f $ **FLOATING
C2044 a_17730_37180# VGND 0.475516f $ **FLOATING
C2045 a_16362_37180# VGND 0.477063f $ **FLOATING
C2046 a_12690_37180# VGND 0.475497f $ **FLOATING
C2047 a_11322_37180# VGND 0.477061f $ **FLOATING
C2048 a_7650_37180# VGND 0.475501f $ **FLOATING
C2049 a_6282_37180# VGND 0.477063f $ **FLOATING
C2050 a_2610_37180# VGND 0.475473f $ **FLOATING
C2051 a_21402_37532# VGND 0.547813f $ **FLOATING
C2052 a_17730_37532# VGND 0.55015f $ **FLOATING
C2053 a_16362_37532# VGND 0.548796f $ **FLOATING
C2054 a_12690_37532# VGND 0.549979f $ **FLOATING
C2055 a_11322_37532# VGND 0.548796f $ **FLOATING
C2056 a_7650_37532# VGND 0.550021f $ **FLOATING
C2057 a_6282_37532# VGND 0.548798f $ **FLOATING
C2058 a_2610_37532# VGND 0.548506f $ **FLOATING
C2059 a_27575_39955# VGND 0.440387f $ **FLOATING
C2060 a_27575_40307# VGND 0.408627f $ **FLOATING
C2061 tt_um_TT06_SAR_done_0.x3.MP1.G VGND 1.07773f
C2062 a_27575_40659# VGND 0.389133f $ **FLOATING
C2063 tt_um_TT06_SAR_done_0.x4.MP0.G VGND 0.822801f
C2064 a_27575_41011# VGND 0.472703f $ **FLOATING
C2065 a_27575_41363# VGND 0.532318f $ **FLOATING
C2066 a_22790_40296# VGND 0.546732f $ **FLOATING
C2067 a_21422_40296# VGND 0.54563f $ **FLOATING
C2068 a_17750_40296# VGND 0.546813f $ **FLOATING
C2069 a_16382_40296# VGND 0.547966f $ **FLOATING
C2070 a_12710_40296# VGND 0.546813f $ **FLOATING
C2071 a_11342_40296# VGND 0.547969f $ **FLOATING
C2072 a_7670_40296# VGND 0.54681f $ **FLOATING
C2073 a_6302_40296# VGND 0.547966f $ **FLOATING
C2074 a_2630_40296# VGND 0.54539f $ **FLOATING
C2075 a_22790_40648# VGND 0.492438f $ **FLOATING
C2076 a_21422_40648# VGND 0.49034f $ **FLOATING
C2077 a_17750_40648# VGND 0.492453f $ **FLOATING
C2078 a_16382_40648# VGND 0.490883f $ **FLOATING
C2079 a_12710_40648# VGND 0.492453f $ **FLOATING
C2080 a_11342_40648# VGND 0.490883f $ **FLOATING
C2081 a_7670_40648# VGND 0.492453f $ **FLOATING
C2082 a_6302_40648# VGND 0.490883f $ **FLOATING
C2083 a_2630_40648# VGND 0.492826f $ **FLOATING
C2084 tt_um_TT06_SAR_done_0.DONE VGND 22.5616f
C2085 a_22790_41000# VGND 0.388777f $ **FLOATING
C2086 a_21422_41000# VGND 0.388174f $ **FLOATING
C2087 a_17750_41000# VGND 0.388174f $ **FLOATING
C2088 a_16382_41000# VGND 0.388174f $ **FLOATING
C2089 a_12710_41000# VGND 0.388174f $ **FLOATING
C2090 a_11342_41000# VGND 0.388174f $ **FLOATING
C2091 a_7670_41000# VGND 0.388174f $ **FLOATING
C2092 a_6302_41000# VGND 0.388174f $ **FLOATING
C2093 a_2630_41000# VGND 0.388638f $ **FLOATING
C2094 a_22790_41352# VGND 0.374594f $ **FLOATING
C2095 a_21422_41352# VGND 0.393558f $ **FLOATING
C2096 a_17750_41352# VGND 0.393558f $ **FLOATING
C2097 a_16382_41352# VGND 0.393558f $ **FLOATING
C2098 a_12710_41352# VGND 0.393558f $ **FLOATING
C2099 a_11342_41352# VGND 0.393558f $ **FLOATING
C2100 a_7670_41352# VGND 0.393558f $ **FLOATING
C2101 a_6302_41352# VGND 0.393558f $ **FLOATING
C2102 a_2630_41352# VGND 0.394022f $ **FLOATING
C2103 SUNSAR_CAPT8B_CV_0.XA4.MP1.G VGND 0.803097f
C2104 SUNSAR_CAPT8B_CV_0.XI14.XA3.MN1.S VGND 0.107737f
C2105 SUNSAR_SAR8B_CV_0.D<0> VGND 5.89609f
C2106 SUNSAR_SAR8B_CV_0.D<1> VGND 13.8115f
C2107 SUNSAR_CAPT8B_CV_0.XH13.XA3.MN1.S VGND 0.107643f
C2108 SUNSAR_CAPT8B_CV_0.XG12.XA3.MN1.S VGND 0.107643f
C2109 SUNSAR_SAR8B_CV_0.D<2> VGND 12.6061f
C2110 SUNSAR_SAR8B_CV_0.D<3> VGND 11.4617f
C2111 SUNSAR_CAPT8B_CV_0.XF11.XA3.MN1.S VGND 0.107643f
C2112 SUNSAR_CAPT8B_CV_0.XE10.XA3.MN1.S VGND 0.107643f
C2113 SUNSAR_SAR8B_CV_0.D<4> VGND 11.8531f
C2114 SUNSAR_SAR8B_CV_0.D<5> VGND 12.723499f
C2115 SUNSAR_CAPT8B_CV_0.XD09.XA3.MN1.S VGND 0.107643f
C2116 SUNSAR_CAPT8B_CV_0.XC08.XA3.MN1.S VGND 0.107643f
C2117 SUNSAR_SAR8B_CV_0.D<6> VGND 12.0371f
C2118 SUNSAR_SAR8B_CV_0.D<7> VGND 17.848501f
C2119 SUNSAR_CAPT8B_CV_0.XB07.XA3.MN1.S VGND 0.107643f
C2120 a_22790_41880# VGND 0.394408f $ **FLOATING
C2121 a_21422_41880# VGND 0.395138f $ **FLOATING
C2122 a_17750_41880# VGND 0.395707f $ **FLOATING
C2123 a_16382_41880# VGND 0.395707f $ **FLOATING
C2124 a_12710_41880# VGND 0.395707f $ **FLOATING
C2125 a_11342_41880# VGND 0.395707f $ **FLOATING
C2126 a_7670_41880# VGND 0.395707f $ **FLOATING
C2127 a_6302_41880# VGND 0.395707f $ **FLOATING
C2128 a_2630_41880# VGND 0.396052f $ **FLOATING
C2129 SUNSAR_CAPT8B_CV_0.XA5.B VGND 1.95346f
C2130 a_22790_42408# VGND 0.410698f $ **FLOATING
C2131 a_21422_42408# VGND 0.389697f $ **FLOATING
C2132 a_17750_42408# VGND 0.390266f $ **FLOATING
C2133 a_16382_42408# VGND 0.390266f $ **FLOATING
C2134 a_12710_42408# VGND 0.390266f $ **FLOATING
C2135 a_11342_42408# VGND 0.390266f $ **FLOATING
C2136 a_7670_42408# VGND 0.390266f $ **FLOATING
C2137 a_6302_42408# VGND 0.390266f $ **FLOATING
C2138 a_2630_42408# VGND 0.390612f $ **FLOATING
C2139 SUNSAR_CAPT8B_CV_0.XA5.XA2.A VGND 1.03543f
C2140 SUNSAR_CAPT8B_CV_0.XI14.XA5.A VGND 1.28758f
C2141 SUNSAR_CAPT8B_CV_0.XH13.XA5.A VGND 1.27933f
C2142 SUNSAR_CAPT8B_CV_0.XG12.XA5.A VGND 1.27933f
C2143 SUNSAR_CAPT8B_CV_0.XF11.XA5.A VGND 1.27933f
C2144 SUNSAR_CAPT8B_CV_0.XE10.XA5.A VGND 1.27933f
C2145 SUNSAR_CAPT8B_CV_0.XD09.XA5.A VGND 1.27933f
C2146 SUNSAR_CAPT8B_CV_0.XC08.XA5.A VGND 1.27933f
C2147 SUNSAR_CAPT8B_CV_0.XB07.XA5.A VGND 1.29578f
C2148 a_22790_42760# VGND 0.378208f $ **FLOATING
C2149 a_21422_42760# VGND 0.393027f $ **FLOATING
C2150 a_17750_42760# VGND 0.393596f $ **FLOATING
C2151 a_16382_42760# VGND 0.393596f $ **FLOATING
C2152 a_12710_42760# VGND 0.393596f $ **FLOATING
C2153 a_11342_42760# VGND 0.393596f $ **FLOATING
C2154 a_7670_42760# VGND 0.393596f $ **FLOATING
C2155 a_6302_42760# VGND 0.393596f $ **FLOATING
C2156 a_2630_42760# VGND 0.393942f $ **FLOATING
C2157 SUNSAR_SAR8B_CV_0.CK_SAMPLE VGND 23.7311f
C2158 SUNSAR_SAR8B_CV_0.EN VGND 10.740701f
C2159 a_22790_43112# VGND 0.388427f $ **FLOATING
C2160 SUNSAR_CAPT8B_CV_0.XI14.XA6.A VGND 1.29446f
C2161 SUNSAR_CAPT8B_CV_0.XH13.XA6.A VGND 1.29655f
C2162 SUNSAR_CAPT8B_CV_0.XG12.XA6.A VGND 1.29655f
C2163 SUNSAR_CAPT8B_CV_0.XF11.XA6.A VGND 1.29655f
C2164 SUNSAR_CAPT8B_CV_0.XE10.XA6.A VGND 1.29655f
C2165 SUNSAR_CAPT8B_CV_0.XD09.XA6.A VGND 1.29655f
C2166 SUNSAR_CAPT8B_CV_0.XC08.XA6.A VGND 1.29655f
C2167 SUNSAR_CAPT8B_CV_0.XB07.XA6.A VGND 1.29893f
C2168 SUNSAR_CAPT8B_CV_0.XA6.A VGND 2.38038f
C2169 a_21422_43288# VGND 0.394124f $ **FLOATING
C2170 a_17750_43288# VGND 0.394693f $ **FLOATING
C2171 a_16382_43288# VGND 0.394693f $ **FLOATING
C2172 a_12710_43288# VGND 0.394693f $ **FLOATING
C2173 a_11342_43288# VGND 0.394693f $ **FLOATING
C2174 a_7670_43288# VGND 0.394693f $ **FLOATING
C2175 a_6302_43288# VGND 0.394693f $ **FLOATING
C2176 a_2630_43288# VGND 0.395039f $ **FLOATING
C2177 SUNSAR_CAPT8B_CV_0.XA6.XA1.MN1.S VGND 0.103608f
C2178 SUNSAR_CAPT8B_CV_0.XA6.B VGND 1.64884f
C2179 a_22790_43640# VGND 0.387806f $ **FLOATING
C2180 SUNSAR_CAPT8B_CV_0.XI14.XA7.MN1.S VGND 0.112889f
C2181 SUNSAR_CAPT8B_CV_0.XI14.XA7.C VGND 2.58298f
C2182 SUNSAR_CAPT8B_CV_0.XI14.XA7.CN VGND 1.69058f
C2183 SUNSAR_CAPT8B_CV_0.XH13.XA7.MN1.S VGND 0.112889f
C2184 SUNSAR_CAPT8B_CV_0.XH13.XA7.CN VGND 1.69315f
C2185 SUNSAR_CAPT8B_CV_0.XH13.XA7.C VGND 2.56583f
C2186 SUNSAR_CAPT8B_CV_0.XG12.XA7.MN1.S VGND 0.112889f
C2187 SUNSAR_CAPT8B_CV_0.XG12.XA7.C VGND 2.61645f
C2188 SUNSAR_CAPT8B_CV_0.XG12.XA7.CN VGND 1.69315f
C2189 SUNSAR_CAPT8B_CV_0.XF11.XA7.MN1.S VGND 0.112889f
C2190 SUNSAR_CAPT8B_CV_0.XF11.XA7.CN VGND 1.69315f
C2191 SUNSAR_CAPT8B_CV_0.XF11.XA7.C VGND 2.61645f
C2192 SUNSAR_CAPT8B_CV_0.XE10.XA7.MN1.S VGND 0.112889f
C2193 SUNSAR_CAPT8B_CV_0.XE10.XA7.C VGND 2.5725f
C2194 SUNSAR_CAPT8B_CV_0.XE10.XA7.CN VGND 1.69797f
C2195 SUNSAR_CAPT8B_CV_0.XD09.XA7.MN1.S VGND 0.112889f
C2196 SUNSAR_CAPT8B_CV_0.XD09.XA7.CN VGND 1.69797f
C2197 SUNSAR_CAPT8B_CV_0.XD09.XA7.C VGND 2.5725f
C2198 SUNSAR_CAPT8B_CV_0.XC08.XA7.MN1.S VGND 0.112889f
C2199 SUNSAR_CAPT8B_CV_0.XC08.XA7.C VGND 2.61716f
C2200 SUNSAR_CAPT8B_CV_0.XC08.XA7.CN VGND 1.69797f
C2201 SUNSAR_CAPT8B_CV_0.XB07.XA7.MN1.S VGND 0.112889f
C2202 SUNSAR_CAPT8B_CV_0.XB07.XA7.CN VGND 1.69726f
C2203 SUNSAR_CAPT8B_CV_0.XB07.XA7.C VGND 2.68306f
C2204 SUNSAR_CAPT8B_CV_0.XA6.XA2.A VGND 0.88269f
C2205 a_21422_43816# VGND 0.390629f $ **FLOATING
C2206 a_17750_43816# VGND 0.391198f $ **FLOATING
C2207 a_16382_43816# VGND 0.391198f $ **FLOATING
C2208 a_12710_43816# VGND 0.391198f $ **FLOATING
C2209 a_11342_43816# VGND 0.391198f $ **FLOATING
C2210 a_7670_43816# VGND 0.391198f $ **FLOATING
C2211 a_6302_43816# VGND 0.391198f $ **FLOATING
C2212 a_2630_43816# VGND 0.391544f $ **FLOATING
C2213 SUNSAR_SAR8B_CV_0.CK_SAMPLE_BSSW VGND 24.501099f
C2214 a_22790_43992# VGND 0.384235f $ **FLOATING
C2215 SUNSAR_CAPT8B_CV_0.XI14.QN VGND 1.23582f
C2216 SUNSAR_CAPT8B_CV_0.XH13.QN VGND 1.23517f
C2217 SUNSAR_CAPT8B_CV_0.XG12.QN VGND 1.23517f
C2218 SUNSAR_CAPT8B_CV_0.XF11.QN VGND 1.23517f
C2219 SUNSAR_CAPT8B_CV_0.XE10.QN VGND 1.26123f
C2220 SUNSAR_CAPT8B_CV_0.XD09.QN VGND 1.26291f
C2221 SUNSAR_CAPT8B_CV_0.XC08.QN VGND 1.26291f
C2222 SUNSAR_CAPT8B_CV_0.XB07.QN VGND 1.26299f
C2223 SUNSAR_CAPT8B_CV_0.XA2.MP0.G VGND 0.5774f
C2224 a_21422_44168# VGND 0.425534f $ **FLOATING
C2225 a_17750_44168# VGND 0.425449f $ **FLOATING
C2226 a_16382_44168# VGND 0.425864f $ **FLOATING
C2227 a_12710_44168# VGND 0.425449f $ **FLOATING
C2228 a_11342_44168# VGND 0.425864f $ **FLOATING
C2229 a_7670_44168# VGND 0.425449f $ **FLOATING
C2230 a_6302_44168# VGND 0.425864f $ **FLOATING
C2231 a_2630_44168# VGND 0.426034f $ **FLOATING
C2232 TIE_L VGND 6.36945f
C2233 a_22790_44344# VGND 0.423601f $ **FLOATING
.ends

