magic
tech sky130A
magscale 1 2
timestamp 1712844206
<< locali >>
rect 12024 44858 27288 44864
rect 12024 44810 12030 44858
rect 12078 44810 27288 44858
rect 12024 44804 27288 44810
rect 22528 44658 27042 44664
rect 22528 44610 22534 44658
rect 22582 44610 27042 44658
rect 22528 44604 27042 44610
rect 29374 44316 31318 44404
rect 24918 40102 26422 40170
rect 26658 39684 26726 43886
rect 27042 41671 29310 41677
rect 27042 41623 27048 41671
rect 27096 41623 29310 41671
rect 27042 41617 29310 41623
rect 26658 39628 26664 39684
rect 26720 39628 26726 39684
rect 26658 39586 26726 39628
<< viali >>
rect 12030 44810 12078 44858
rect 27288 44804 27348 44864
rect 22534 44610 22582 44658
rect 27042 44604 27102 44664
rect 31318 44316 31406 44404
rect 26658 43886 26726 43954
rect 22372 40112 22428 40168
rect 26422 40102 26490 40170
rect 27048 41623 27096 41671
rect 29310 41617 29370 41677
rect 26664 39628 26720 39684
<< metal1 >>
rect 12242 44892 12302 44898
rect 11933 44804 11939 44864
rect 11999 44858 12090 44864
rect 11999 44810 12030 44858
rect 12078 44810 12090 44858
rect 11999 44804 12090 44810
rect 7358 44714 7418 44720
rect 12242 44714 12302 44832
rect 27282 44864 27354 44876
rect 27282 44804 27288 44864
rect 27348 44804 27354 44864
rect 27282 44792 27354 44804
rect 7418 44654 12302 44714
rect 22396 44664 22456 44670
rect 27036 44664 27108 44676
rect 7358 44648 7418 44654
rect 22456 44658 22594 44664
rect 22456 44610 22534 44658
rect 22582 44610 22594 44658
rect 22456 44604 22594 44610
rect 27036 44604 27042 44664
rect 27102 44604 27108 44664
rect 22396 44598 22456 44604
rect 27036 44592 27108 44604
rect 17370 44482 17376 44542
rect 17436 44482 23300 44542
rect 23360 44482 23366 44542
rect 26652 43954 26732 43966
rect 26500 43886 26506 43954
rect 26574 43886 26658 43954
rect 26726 43886 26732 43954
rect 26652 43874 26732 43886
rect 27042 41671 27102 44592
rect 27042 41623 27048 41671
rect 27096 41623 27102 41671
rect 27042 41597 27102 41623
rect 27288 40558 27348 44792
rect 31312 44404 31412 44416
rect 31312 44316 31318 44404
rect 31406 44316 31412 44404
rect 31312 44304 31412 44316
rect 31318 44216 31406 44304
rect 31318 44122 31406 44128
rect 29304 41677 29376 41689
rect 29304 41617 29310 41677
rect 29370 41617 29376 41677
rect 29304 41605 29376 41617
rect 29310 40910 29370 41605
rect 22366 40168 22434 40180
rect 22366 40112 22372 40168
rect 22428 40112 22434 40168
rect 22366 40034 22434 40112
rect 26416 40170 26496 40182
rect 26416 40102 26422 40170
rect 26490 40102 27336 40170
rect 26416 40090 26496 40102
rect 22360 39966 22366 40034
rect 22434 39966 22440 40034
rect 26658 39684 26726 39696
rect 26658 39628 26664 39684
rect 26720 39628 26726 39684
rect 26658 39468 26726 39628
rect 14848 7490 14946 7716
<< via1 >>
rect 11939 44804 11999 44864
rect 12242 44832 12302 44892
rect 7358 44654 7418 44714
rect 22396 44604 22456 44664
rect 17376 44482 17436 44542
rect 23300 44482 23360 44542
rect 26506 43886 26574 43954
rect 31318 44128 31406 44216
rect 22366 39966 22434 40034
<< metal2 >>
rect 11494 44921 11581 44937
rect 11939 44933 11999 44935
rect 11494 44865 11503 44921
rect 11559 44865 11581 44921
rect 11932 44877 11941 44933
rect 11997 44877 12006 44933
rect 11494 44855 11581 44865
rect 11939 44864 11999 44877
rect 3150 44588 3210 44780
rect 7193 44696 7202 44756
rect 7262 44714 7271 44756
rect 8172 44750 8228 44757
rect 8170 44748 8230 44750
rect 7262 44696 7358 44714
rect 7202 44654 7358 44696
rect 7418 44654 7424 44714
rect 8170 44692 8172 44748
rect 8228 44692 8230 44748
rect 3150 44532 3152 44588
rect 3208 44532 3210 44588
rect 3150 44336 3210 44532
rect 6472 44450 6528 44457
rect 6470 44448 6530 44450
rect 6470 44392 6472 44448
rect 6528 44392 6530 44448
rect 6470 44328 6530 44392
rect 8170 44318 8230 44692
rect 11501 44730 11561 44855
rect 12236 44832 12242 44892
rect 12302 44832 12326 44892
rect 12386 44832 12395 44892
rect 17378 44888 17434 44895
rect 17376 44886 17436 44888
rect 11939 44798 11999 44804
rect 17376 44830 17378 44886
rect 17434 44830 17436 44886
rect 11501 44670 11880 44730
rect 11820 44609 11880 44670
rect 11512 44590 11568 44597
rect 11510 44588 11570 44590
rect 11510 44532 11512 44588
rect 11568 44532 11570 44588
rect 11820 44549 15945 44609
rect 16532 44590 16588 44597
rect 11510 44338 11570 44532
rect 13212 44450 13268 44457
rect 13210 44448 13270 44450
rect 13210 44392 13212 44448
rect 13268 44392 13270 44448
rect 13210 44334 13270 44392
rect 15885 44408 15945 44549
rect 15885 44339 15945 44348
rect 16530 44588 16590 44590
rect 16530 44532 16532 44588
rect 16588 44532 16590 44588
rect 16530 44338 16590 44532
rect 17376 44542 17436 44830
rect 21612 44848 21668 44888
rect 21610 44792 21612 44828
rect 21668 44792 21670 44828
rect 18250 44708 18310 44710
rect 18243 44652 18252 44708
rect 18308 44652 18317 44708
rect 17376 44476 17436 44482
rect 18250 44342 18310 44652
rect 21610 44334 21670 44792
rect 22266 44662 22396 44664
rect 22259 44606 22268 44662
rect 22324 44606 22396 44662
rect 22266 44604 22396 44606
rect 22456 44604 22462 44664
rect 23298 44548 23358 44828
rect 23298 44542 23360 44548
rect 23298 44482 23300 44542
rect 23298 44476 23360 44482
rect 23298 44328 23358 44476
rect 31312 44128 31318 44216
rect 31406 44128 31412 44216
rect 31318 44052 31406 44128
rect 26506 43954 26574 43960
rect 31318 43955 31406 43964
rect 24746 43886 26506 43954
rect 26506 43880 26574 43886
rect 24846 43069 26214 43074
rect 24846 43011 26151 43069
rect 26209 43011 26218 43069
rect 24846 43006 26214 43011
rect 24846 42646 25272 42714
rect 25340 42646 25349 42714
rect 22366 40034 22434 40040
rect 22366 39889 22434 39966
rect 22362 39831 22371 39889
rect 22429 39831 22438 39889
rect 22366 39826 22434 39831
rect 2646 39595 2706 39599
rect 2641 39590 2795 39595
rect 2641 39530 2646 39590
rect 2706 39530 2795 39590
rect 6862 39531 6871 39589
rect 6929 39531 6938 39589
rect 7766 39569 7834 39674
rect 2641 39525 2795 39530
rect 2646 39521 2706 39525
rect 7762 39511 7771 39569
rect 7829 39511 7838 39569
rect 11922 39551 11931 39609
rect 11989 39551 11998 39609
rect 12782 39551 12791 39609
rect 12849 39551 12858 39609
rect 16942 39551 16951 39609
rect 17009 39551 17018 39609
rect 17822 39551 17831 39609
rect 17889 39551 17898 39609
rect 21982 39531 21991 39589
rect 22049 39531 22058 39589
rect 7766 39506 7834 39511
rect 22851 39414 22909 39418
rect 22846 39409 29506 39414
rect 22846 39351 22851 39409
rect 22909 39351 29506 39409
rect 22846 39346 29506 39351
rect 29574 39346 29583 39414
rect 22851 39342 22909 39346
rect 20515 39214 20573 39218
rect 20510 39209 26146 39214
rect 20510 39151 20515 39209
rect 20573 39151 26146 39209
rect 20510 39146 26146 39151
rect 26214 39146 26223 39214
rect 20515 39142 20573 39146
rect 8377 39114 8435 39118
rect 6166 39109 6866 39114
rect 6166 39051 6216 39109
rect 6274 39051 6866 39109
rect 6166 39046 6866 39051
rect 6934 39046 6943 39114
rect 7757 39046 7766 39114
rect 7834 39109 8440 39114
rect 7834 39051 8377 39109
rect 8435 39051 8440 39109
rect 11256 39094 11314 39098
rect 11926 39094 11994 39103
rect 7834 39046 8440 39051
rect 11251 39089 11926 39094
rect 8377 39042 8435 39046
rect 11251 39031 11256 39089
rect 11314 39031 11926 39089
rect 11251 39026 11926 39031
rect 12777 39026 12786 39094
rect 12854 39089 13480 39094
rect 12854 39031 13417 39089
rect 13475 39031 13484 39089
rect 16277 39046 16286 39114
rect 16354 39109 17014 39114
rect 16354 39051 16951 39109
rect 17009 39051 17018 39109
rect 17826 39094 17894 39103
rect 16354 39046 17014 39051
rect 12854 39026 13480 39031
rect 17894 39089 18520 39094
rect 17894 39031 18457 39089
rect 18515 39031 18524 39089
rect 17894 39026 18520 39031
rect 11256 39022 11314 39026
rect 11926 39017 11994 39026
rect 17826 39017 17894 39026
rect 22572 35824 22640 35833
rect 22572 35747 22640 35756
rect 25014 34112 25340 34116
rect 22044 34111 25342 34112
rect 22044 34053 25277 34111
rect 25335 34053 25344 34111
rect 22044 34044 25342 34053
rect 20114 30124 20510 30192
rect 20578 30124 20587 30192
rect 12694 413 12814 2926
rect 14498 695 14618 2932
rect 14498 585 14503 695
rect 14613 585 14618 695
rect 14498 580 14618 585
rect 14503 576 14613 580
rect 12690 303 12699 413
rect 12809 303 12818 413
rect 12694 298 12814 303
<< via2 >>
rect 11503 44865 11559 44921
rect 11941 44877 11997 44933
rect 7202 44696 7262 44756
rect 8172 44692 8228 44748
rect 3152 44532 3208 44588
rect 6472 44392 6528 44448
rect 12326 44832 12386 44892
rect 17378 44830 17434 44886
rect 11512 44532 11568 44588
rect 13212 44392 13268 44448
rect 15885 44348 15945 44408
rect 16532 44532 16588 44588
rect 21612 44792 21668 44848
rect 18252 44652 18308 44708
rect 22268 44606 22324 44662
rect 31318 43964 31406 44052
rect 26151 43011 26209 43069
rect 25272 42646 25340 42714
rect 22371 39831 22429 39889
rect 2646 39530 2706 39590
rect 6871 39531 6929 39589
rect 7771 39511 7829 39569
rect 11931 39551 11989 39609
rect 12791 39551 12849 39609
rect 16951 39551 17009 39609
rect 17831 39551 17889 39609
rect 21991 39531 22049 39589
rect 22851 39351 22909 39409
rect 29506 39346 29574 39414
rect 20515 39151 20573 39209
rect 26146 39146 26214 39214
rect 6216 39051 6274 39109
rect 6866 39046 6934 39114
rect 7766 39046 7834 39114
rect 8377 39051 8435 39109
rect 11256 39031 11314 39089
rect 11926 39026 11994 39094
rect 12786 39026 12854 39094
rect 13417 39031 13475 39089
rect 16286 39046 16354 39114
rect 16951 39051 17009 39109
rect 17826 39026 17894 39094
rect 18457 39031 18515 39089
rect 22572 35756 22640 35824
rect 25277 34053 25335 34111
rect 20510 30124 20578 30192
rect 14503 585 14613 695
rect 12699 303 12809 413
<< metal3 >>
rect 11830 44937 12002 44938
rect 5942 44861 5948 44925
rect 6012 44923 6018 44925
rect 11494 44923 11581 44937
rect 6012 44921 11581 44923
rect 6012 44865 11503 44921
rect 11559 44865 11581 44921
rect 11830 44873 11836 44937
rect 11900 44933 12002 44937
rect 11900 44877 11941 44933
rect 11997 44877 12002 44933
rect 12321 44892 12391 44897
rect 12321 44888 12326 44892
rect 11900 44873 12002 44877
rect 11830 44872 12002 44873
rect 6012 44863 11581 44865
rect 6012 44861 6018 44863
rect 11494 44855 11581 44863
rect 12218 44832 12326 44888
rect 12386 44888 12391 44892
rect 17373 44888 17439 44891
rect 12386 44886 17439 44888
rect 12386 44832 17378 44886
rect 12218 44830 17378 44832
rect 17434 44830 17439 44886
rect 12218 44828 17439 44830
rect 12321 44827 12391 44828
rect 17373 44825 17439 44828
rect 17718 44788 17724 44852
rect 17788 44850 17794 44852
rect 21607 44850 21673 44853
rect 17788 44848 21673 44850
rect 17788 44792 21612 44848
rect 21668 44792 21673 44848
rect 17788 44790 21673 44792
rect 17788 44788 17794 44790
rect 21607 44787 21673 44790
rect 6978 44694 6984 44758
rect 7048 44756 7054 44758
rect 7197 44756 7267 44761
rect 7048 44696 7202 44756
rect 7262 44696 7267 44756
rect 7048 44694 7054 44696
rect 7197 44691 7267 44696
rect 8167 44750 8233 44753
rect 14038 44750 14044 44752
rect 8167 44748 14044 44750
rect 8167 44692 8172 44748
rect 8228 44692 14044 44748
rect 8167 44690 14044 44692
rect 8167 44687 8233 44690
rect 14038 44688 14044 44690
rect 14108 44688 14114 44752
rect 16982 44648 16988 44712
rect 17052 44710 17058 44712
rect 18247 44710 18313 44713
rect 17052 44708 18313 44710
rect 17052 44652 18252 44708
rect 18308 44652 18313 44708
rect 17052 44650 18313 44652
rect 17052 44648 17058 44650
rect 18247 44647 18313 44650
rect 22263 44662 22329 44667
rect 22263 44606 22268 44662
rect 22324 44606 22329 44662
rect 22263 44601 22329 44606
rect 22894 44664 22962 44694
rect 3147 44590 3213 44593
rect 11162 44590 11168 44592
rect 3147 44588 11168 44590
rect 3147 44532 3152 44588
rect 3208 44532 11168 44588
rect 3147 44530 11168 44532
rect 3147 44527 3213 44530
rect 11162 44528 11168 44530
rect 11232 44528 11238 44592
rect 11507 44590 11573 44593
rect 16252 44592 16316 44598
rect 14774 44590 14780 44592
rect 11507 44588 14780 44590
rect 11507 44532 11512 44588
rect 11568 44532 14780 44588
rect 11507 44530 14780 44532
rect 11507 44527 11573 44530
rect 14774 44528 14780 44530
rect 14844 44528 14850 44592
rect 16527 44590 16593 44593
rect 16316 44588 16593 44590
rect 16316 44532 16532 44588
rect 16588 44532 16593 44588
rect 16316 44530 16593 44532
rect 16252 44522 16316 44528
rect 16527 44527 16593 44530
rect 6467 44450 6533 44453
rect 12862 44450 12868 44452
rect 6467 44448 12868 44450
rect 6467 44392 6472 44448
rect 6528 44392 12868 44448
rect 6467 44390 12868 44392
rect 6467 44387 6533 44390
rect 12862 44388 12868 44390
rect 12932 44388 12938 44452
rect 13207 44450 13273 44453
rect 15510 44450 15516 44452
rect 13207 44448 15516 44450
rect 13207 44392 13212 44448
rect 13268 44392 15516 44448
rect 13207 44390 15516 44392
rect 13207 44387 13273 44390
rect 15510 44388 15516 44390
rect 15580 44388 15586 44452
rect 15880 44408 15950 44413
rect 22266 44408 22326 44601
rect 15880 44348 15885 44408
rect 15945 44348 22326 44408
rect 22894 44596 27006 44664
rect 15880 44343 15950 44348
rect 22894 44294 22962 44596
rect 26938 44186 27006 44596
rect 26488 44118 30966 44186
rect 31034 44118 31040 44186
rect 31313 44052 31411 44057
rect 31313 43964 31318 44052
rect 31406 43964 31411 44052
rect 31313 43959 31411 43964
rect 31318 43852 31406 43959
rect 31318 43758 31406 43764
rect 26146 43069 26214 43074
rect 26146 43011 26151 43069
rect 26209 43011 26214 43069
rect 25267 42714 25345 42719
rect 25267 42646 25272 42714
rect 25340 42646 25345 42714
rect 25267 42641 25345 42646
rect 2641 39590 2711 39595
rect 2641 39530 2646 39590
rect 2706 39530 2711 39590
rect 2641 29275 2711 39530
rect 4500 39424 5100 39480
rect 4410 39423 5210 39424
rect 4410 39125 4651 39423
rect 4949 39125 5210 39423
rect 6211 39134 6279 39246
rect 4410 39124 5210 39125
rect 4500 39100 5100 39124
rect 6146 39109 6279 39134
rect 6146 39051 6216 39109
rect 6274 39051 6279 39109
rect 6146 39026 6279 39051
rect 3888 38448 5778 38632
rect 3042 38312 3226 38318
rect 3042 37708 3226 38128
rect 6211 30970 6279 39026
rect 6406 38318 6590 40792
rect 6866 39589 6934 39594
rect 6866 39531 6871 39589
rect 6929 39531 6934 39589
rect 6866 39119 6934 39531
rect 7766 39569 7834 39574
rect 7766 39511 7771 39569
rect 7829 39511 7834 39569
rect 7766 39119 7834 39511
rect 6861 39114 6939 39119
rect 6861 39046 6866 39114
rect 6934 39046 6939 39114
rect 6861 39041 6939 39046
rect 7761 39114 7839 39119
rect 7761 39046 7766 39114
rect 7834 39046 7839 39114
rect 7761 39041 7839 39046
rect 6386 38312 6590 38318
rect 6570 38128 6590 38312
rect 8102 38278 8286 40572
rect 9450 39423 10270 39424
rect 6386 38088 6590 38128
rect 8082 38272 8286 38278
rect 8266 38088 8286 38272
rect 6386 37768 6570 38088
rect 8082 37988 8286 38088
rect 8372 39109 8440 39286
rect 9450 39125 9691 39423
rect 9989 39125 10270 39423
rect 9450 39124 10270 39125
rect 8372 39051 8377 39109
rect 8435 39051 8440 39109
rect 8082 37848 8266 37988
rect 8372 27636 8440 39051
rect 11251 39089 11319 39126
rect 11251 39031 11256 39089
rect 11314 39031 11319 39089
rect 8908 38428 10818 38612
rect 11251 28232 11319 39031
rect 11446 38338 11630 40612
rect 11926 39609 11994 39614
rect 11926 39551 11931 39609
rect 11989 39551 11994 39609
rect 11926 39099 11994 39551
rect 12786 39609 12854 39614
rect 12786 39551 12791 39609
rect 12849 39551 12854 39609
rect 12786 39099 12854 39551
rect 11921 39094 11999 39099
rect 11921 39026 11926 39094
rect 11994 39026 11999 39094
rect 11921 39021 11999 39026
rect 12781 39094 12859 39099
rect 12781 39026 12786 39094
rect 12854 39026 12859 39094
rect 12781 39021 12859 39026
rect 11426 38332 11630 38338
rect 11610 38148 11630 38332
rect 11426 38108 11630 38148
rect 11426 37808 11610 38108
rect 13142 38048 13326 40632
rect 14640 39424 15180 39460
rect 13412 39089 13480 39186
rect 14640 39124 14730 39424
rect 15030 39124 15180 39424
rect 14640 39100 15180 39124
rect 16291 39119 16359 39266
rect 16281 39114 16359 39119
rect 13412 39031 13417 39089
rect 13475 39031 13480 39089
rect 16281 39046 16286 39114
rect 16354 39046 16359 39114
rect 16281 39041 16359 39046
rect 13122 38012 13306 38018
rect 13122 37822 13306 37828
rect 13412 26386 13480 39031
rect 13914 38468 15832 38652
rect 16291 29204 16359 39041
rect 16486 38298 16670 40172
rect 16946 39609 17014 39614
rect 16946 39551 16951 39609
rect 17009 39551 17014 39609
rect 16946 39109 17014 39551
rect 16946 39051 16951 39109
rect 17009 39051 17014 39109
rect 17826 39609 17894 39614
rect 17826 39551 17831 39609
rect 17889 39551 17894 39609
rect 17826 39099 17894 39551
rect 16946 39046 17014 39051
rect 17821 39094 17899 39099
rect 17821 39026 17826 39094
rect 17894 39026 17899 39094
rect 17821 39021 17899 39026
rect 18182 38338 18366 40172
rect 22366 39889 22434 39894
rect 22366 39831 22371 39889
rect 22429 39831 22434 39889
rect 21986 39589 22054 39594
rect 21986 39531 21991 39589
rect 22049 39531 22054 39589
rect 19530 39423 20310 39424
rect 16466 38292 16670 38298
rect 16650 38108 16670 38292
rect 16466 38088 16670 38108
rect 18162 38332 18366 38338
rect 18346 38148 18366 38332
rect 16466 37848 16650 38088
rect 18162 37888 18366 38148
rect 18182 37848 18366 37888
rect 18452 39089 18520 39206
rect 19530 39125 19751 39423
rect 20049 39125 20310 39423
rect 21986 39354 22054 39531
rect 21331 39286 22054 39354
rect 19530 39124 20310 39125
rect 20510 39209 20578 39214
rect 20510 39151 20515 39209
rect 20573 39151 20578 39209
rect 18452 39031 18457 39089
rect 18515 39031 18520 39089
rect 18452 26436 18520 39031
rect 18954 38488 20292 38672
rect 20510 30197 20578 39151
rect 21331 31422 21399 39286
rect 22366 38434 22434 39831
rect 22846 39409 22914 39594
rect 22846 39351 22851 39409
rect 22909 39351 22914 39409
rect 22846 39346 22914 39351
rect 22366 38366 22640 38434
rect 21506 38312 21690 38318
rect 21506 37928 21690 38128
rect 22572 35829 22640 38366
rect 23202 38352 23386 40172
rect 23202 37588 23386 38168
rect 22567 35824 22645 35829
rect 22567 35756 22572 35824
rect 22640 35756 22645 35824
rect 22567 35751 22645 35756
rect 25272 34111 25340 42641
rect 26146 39219 26214 43011
rect 26141 39214 26219 39219
rect 26141 39146 26146 39214
rect 26214 39146 26219 39214
rect 26141 39141 26219 39146
rect 28007 38336 28207 40248
rect 28799 39118 28999 40176
rect 29506 39654 29574 39660
rect 29506 39419 29574 39586
rect 29501 39414 29579 39419
rect 29501 39346 29506 39414
rect 29574 39346 29579 39414
rect 29501 39341 29579 39346
rect 28799 39081 29260 39118
rect 28799 38783 28939 39081
rect 29237 38783 29260 39081
rect 28799 38759 29260 38783
rect 28906 38758 29260 38759
rect 28007 38130 28207 38136
rect 28938 37006 29238 38758
rect 28938 36700 29238 36706
rect 25272 34053 25277 34111
rect 25335 34053 25340 34111
rect 25272 34048 25340 34053
rect 20505 30192 20583 30197
rect 20505 30124 20510 30192
rect 20578 30124 20583 30192
rect 20505 30119 20583 30124
rect 22748 22486 22862 22726
rect 23032 22486 23146 22726
rect 22760 22152 22970 22248
rect 12304 7488 12406 7714
rect 14848 7490 14946 7716
rect 12306 3738 12416 3966
rect 14846 3736 14956 3964
rect 31313 700 31431 705
rect 14498 699 31432 700
rect 14498 695 31313 699
rect 14498 585 14503 695
rect 14613 585 31313 695
rect 14498 581 31313 585
rect 31431 581 31432 699
rect 14498 580 31432 581
rect 31313 575 31431 580
rect 12694 417 27016 418
rect 12694 413 26897 417
rect 12694 303 12699 413
rect 12809 303 26897 413
rect 12694 299 26897 303
rect 27015 299 27021 417
rect 12694 298 27016 299
<< via3 >>
rect 5948 44861 6012 44925
rect 11836 44873 11900 44937
rect 17724 44788 17788 44852
rect 6984 44694 7048 44758
rect 14044 44688 14108 44752
rect 16988 44648 17052 44712
rect 11168 44528 11232 44592
rect 14780 44528 14844 44592
rect 16252 44528 16316 44592
rect 12868 44388 12932 44452
rect 15516 44388 15580 44452
rect 30966 44118 31034 44186
rect 31318 43764 31406 43852
rect 4651 39125 4949 39423
rect 3042 38128 3226 38312
rect 6386 38128 6570 38312
rect 8082 38088 8266 38272
rect 9691 39125 9989 39423
rect 11426 38148 11610 38332
rect 14730 39124 15030 39424
rect 13122 37828 13306 38012
rect 16466 38108 16650 38292
rect 18162 38148 18346 38332
rect 19751 39125 20049 39423
rect 21506 38128 21690 38312
rect 23202 38168 23386 38352
rect 29506 39586 29574 39654
rect 28939 38783 29237 39081
rect 28007 38136 28207 38336
rect 28938 36706 29238 37006
rect 31313 581 31431 699
rect 26897 299 27015 417
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44982 1594 45152
rect 1534 44892 1594 44922
rect 2270 44982 2330 45152
rect 2270 44892 2330 44922
rect 3006 44984 3066 45152
rect 3006 44892 3066 44924
rect 3742 44988 3802 45152
rect 3742 44892 3802 44928
rect 4478 44984 4538 45152
rect 4478 44892 4538 44924
rect 5214 44986 5274 45152
rect 5950 44926 6010 45152
rect 6686 44986 6746 45152
rect 5214 44892 5274 44926
rect 5947 44925 6013 44926
rect 798 44832 5799 44892
rect 5947 44861 5948 44925
rect 6012 44861 6013 44925
rect 6686 44892 6746 44926
rect 7422 44982 7482 45152
rect 7422 44892 7482 44922
rect 8158 44984 8218 45152
rect 8158 44892 8218 44924
rect 8894 44982 8954 45152
rect 8894 44892 8954 44922
rect 9630 44982 9690 45152
rect 9630 44892 9690 44922
rect 10366 44982 10426 45152
rect 10366 44892 10426 44922
rect 11102 44988 11162 45152
rect 11838 44938 11898 45152
rect 11102 44892 11162 44928
rect 11835 44937 11901 44938
rect 5947 44860 6013 44861
rect 6610 44832 11445 44892
rect 11835 44873 11836 44937
rect 11900 44873 11901 44937
rect 11835 44872 11901 44873
rect 5739 44756 6820 44772
rect 6983 44758 7049 44759
rect 6983 44756 6984 44758
rect 5739 44712 6984 44756
rect 6606 44696 6984 44712
rect 6983 44694 6984 44696
rect 7048 44694 7049 44758
rect 12574 44730 12634 45152
rect 13310 44873 13370 45152
rect 12867 44807 13373 44873
rect 6983 44693 7049 44694
rect 11170 44670 12634 44730
rect 11170 44593 11230 44670
rect 11167 44592 11233 44593
rect 11167 44528 11168 44592
rect 11232 44528 11233 44592
rect 11167 44527 11233 44528
rect 12870 44453 12930 44807
rect 14046 44753 14106 45152
rect 14043 44752 14109 44753
rect 14043 44688 14044 44752
rect 14108 44688 14109 44752
rect 14043 44687 14109 44688
rect 14782 44593 14842 45152
rect 14779 44592 14845 44593
rect 14779 44528 14780 44592
rect 14844 44528 14845 44592
rect 14779 44527 14845 44528
rect 15518 44453 15578 45152
rect 16254 44593 16314 45152
rect 16990 44713 17050 45152
rect 17726 44853 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 45014 29562 45152
rect 29502 44900 29574 45014
rect 30238 44952 30298 45152
rect 30974 45054 31034 45152
rect 17723 44852 17789 44853
rect 17723 44788 17724 44852
rect 17788 44788 17789 44852
rect 17723 44787 17789 44788
rect 16987 44712 17053 44713
rect 16987 44648 16988 44712
rect 17052 44648 17053 44712
rect 16987 44647 17053 44648
rect 16251 44592 16317 44593
rect 16251 44528 16252 44592
rect 16316 44528 16317 44592
rect 16251 44527 16317 44528
rect 12867 44452 12933 44453
rect 12867 44388 12868 44452
rect 12932 44388 12933 44452
rect 12867 44387 12933 44388
rect 15515 44452 15581 44453
rect 15515 44388 15516 44452
rect 15580 44388 15581 44452
rect 15515 44387 15581 44388
rect 200 39424 500 44152
rect 29506 39655 29574 44900
rect 30966 44187 31034 45054
rect 31710 44952 31770 45152
rect 30965 44186 31035 44187
rect 30965 44118 30966 44186
rect 31034 44118 31035 44186
rect 30965 44117 31035 44118
rect 31200 43852 31500 44152
rect 31200 43764 31318 43852
rect 31406 43764 31500 43852
rect 29505 39654 29575 39655
rect 29505 39586 29506 39654
rect 29574 39586 29575 39654
rect 29505 39585 29575 39586
rect 14729 39424 15031 39425
rect 200 39423 14730 39424
rect 200 39125 4651 39423
rect 4949 39125 9691 39423
rect 9989 39125 14730 39423
rect 200 39124 14730 39125
rect 15030 39423 24250 39424
rect 15030 39125 19751 39423
rect 20049 39125 24250 39423
rect 15030 39124 24250 39125
rect 200 1000 500 39124
rect 14729 39123 15031 39124
rect 23950 39082 24250 39124
rect 23950 39081 30928 39082
rect 23950 38783 28939 39081
rect 29237 38783 30928 39081
rect 23950 38782 30928 38783
rect 31200 38382 31500 43764
rect 1490 38352 31500 38382
rect 1490 38332 23202 38352
rect 1490 38312 11426 38332
rect 1490 38128 3042 38312
rect 3226 38128 6386 38312
rect 6570 38272 11426 38312
rect 6570 38128 8082 38272
rect 1490 38088 8082 38128
rect 8266 38148 11426 38272
rect 11610 38292 18162 38332
rect 11610 38148 16466 38292
rect 8266 38108 16466 38148
rect 16650 38148 18162 38292
rect 18346 38312 23202 38332
rect 18346 38148 21506 38312
rect 16650 38128 21506 38148
rect 21690 38168 23202 38312
rect 23386 38336 31500 38352
rect 23386 38168 28007 38336
rect 21690 38136 28007 38168
rect 28207 38136 31500 38336
rect 21690 38128 31500 38136
rect 16650 38108 31500 38128
rect 8266 38088 31500 38108
rect 1490 38082 31500 38088
rect 13122 38013 13306 38082
rect 13121 38012 13307 38013
rect 13121 37828 13122 38012
rect 13306 37828 13307 38012
rect 13121 37827 13307 37828
rect 26976 36316 27080 38082
rect 28937 37006 29239 37007
rect 28937 36706 28938 37006
rect 29238 36706 29239 37006
rect 28937 36705 29239 36706
rect 28938 36398 29238 36705
rect 22748 22486 22862 22726
rect 23032 22486 23146 22726
rect 22752 22152 22974 22256
rect 12304 7488 12406 7714
rect 12306 3738 12416 3966
rect 14846 3736 14956 3964
rect 31200 1000 31500 38082
rect 31312 699 31432 700
rect 31312 581 31313 699
rect 31431 581 31432 699
rect 26896 417 27016 418
rect 26896 299 26897 417
rect 27015 299 27016 417
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 299
rect 31312 0 31432 581
<< rmetal4 >>
rect 798 44892 858 44952
rect 1534 44922 1594 44982
rect 2270 44922 2330 44982
rect 3006 44924 3066 44984
rect 3742 44928 3802 44988
rect 4478 44924 4538 44984
rect 5214 44926 5274 44986
rect 6686 44926 6746 44986
rect 7422 44922 7482 44982
rect 8158 44924 8218 44984
rect 8894 44922 8954 44982
rect 9630 44922 9690 44982
rect 10366 44922 10426 44982
rect 11102 44928 11162 44988
rect 5739 44772 5799 44832
rect 6696 44772 6756 44832
use sky130_fd_pr__cap_mim_m3_1_XS736D  sky130_fd_pr__cap_mim_m3_1_XS736D_0
timestamp 1710669355
transform -1 0 28962 0 1 18780
box -1986 -17640 1986 17640
use SUNSAR_CAPT8B_CV  SUNSAR_CAPT8B_CV_0 ../SUN_SAR9B_SKY130NM
timestamp 1712843141
transform 1 0 2306 0 1 40314
box -225 -788 22902 4180
use SUNSAR_SAR8B_CV  SUNSAR_SAR8B_CV_0 ../SUN_SAR9B_SKY130NM
timestamp 1712843141
transform 1 0 2448 0 1 2648
box -1922 -1864 24278 37062
use tt_um_TT06_SAR_done  tt_um_TT06_SAR_done_0
timestamp 1712843141
transform 1 0 27251 0 1 39973
box -180 -132 2700 1540
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 31200 1000 31500 44152 0 FreeSans 2000 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 6250 44712 6310 44772 0 FreeSans 320 0 0 0 TIE_L
flabel metal4 5398 44832 5458 44892 0 FreeSans 320 0 0 0 TIE_L2
flabel metal4 6864 44832 6924 44892 0 FreeSans 320 0 0 0 TIE_L1
flabel metal4 s 200 1000 500 44152 0 FreeSans 2000 90 0 0 VPWR
port 51 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
